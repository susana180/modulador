// This is the unpowered netlist.
module OQPSK_PS_RCOSINE2 (BitIn,
    CLK,
    EN,
    RST,
    I,
    Q,
    addI,
    addQ);
 input BitIn;
 input CLK;
 input EN;
 input RST;
 output [12:0] I;
 output [12:0] Q;
 output [5:0] addI;
 output [5:0] addQ;

 wire \Reg_Delay_Q.In ;
 wire \Reg_Delay_Q.Out ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire \bit2symb.regi ;
 wire \p_shaping_I.bit_in ;
 wire \p_shaping_I.bit_in_1 ;
 wire \p_shaping_I.bit_in_2 ;
 wire \p_shaping_I.counter[0] ;
 wire \p_shaping_I.counter[1] ;
 wire \p_shaping_I.ctl_1 ;
 wire \p_shaping_Q.bit_in_1 ;
 wire \p_shaping_Q.bit_in_2 ;
 wire \p_shaping_Q.counter[0] ;
 wire \p_shaping_Q.counter[1] ;
 wire \p_shaping_Q.ctl_1 ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire clknet_0_CLK;
 wire clknet_1_0__leaf_CLK;
 wire clknet_1_1__leaf_CLK;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1444_ (.I(net30),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1445_ (.I(_1258_),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1446_ (.I(_1269_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1447_ (.I(net47),
    .Z(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1448_ (.I(net34),
    .Z(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1449_ (.I(_1302_),
    .Z(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1450_ (.I(net31),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1451_ (.I(_1324_),
    .Z(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1452_ (.I(net33),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1453_ (.I(_1346_),
    .Z(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1454_ (.I(net32),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1455_ (.I(_1368_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1456_ (.A1(_1335_),
    .A2(_1357_),
    .A3(_1379_),
    .ZN(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1457_ (.A1(_1280_),
    .A2(_1291_),
    .A3(_1313_),
    .A4(_1389_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1458_ (.I(_1400_),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1459_ (.I(_1411_),
    .Z(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1460_ (.I(net46),
    .Z(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1461_ (.I(_1432_),
    .Z(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1462_ (.I(_1443_),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1463_ (.I(_0036_),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1464_ (.I(net37),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1465_ (.I(_0058_),
    .Z(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1466_ (.I(_0069_),
    .Z(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1467_ (.I(net39),
    .Z(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1468_ (.I(_0091_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1469_ (.I(_0102_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1470_ (.I(net38),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1471_ (.I(_0124_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1472_ (.I(_0135_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1473_ (.A1(_0080_),
    .A2(_0113_),
    .A3(_0145_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1474_ (.A1(_0047_),
    .A2(_0156_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1475_ (.I(net45),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1476_ (.I(net44),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1477_ (.I(_0189_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1478_ (.A1(_0178_),
    .A2(_0200_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1479_ (.I(_0210_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1480_ (.I(_0058_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1481_ (.I(_0232_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1482_ (.I(_0091_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1483_ (.I(_0254_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1484_ (.A1(_0243_),
    .A2(_0265_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1485_ (.A1(_0091_),
    .A2(_0135_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1486_ (.I(_0287_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1487_ (.I(net46),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1488_ (.I(_0308_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1489_ (.A1(_0319_),
    .A2(_0145_),
    .B(_0113_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1490_ (.A1(_0276_),
    .A2(_0297_),
    .A3(_0330_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1491_ (.I(_0069_),
    .Z(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1492_ (.I(_0351_),
    .Z(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1493_ (.I(_0102_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1494_ (.I(_0373_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1495_ (.I(net38),
    .Z(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1496_ (.I(_0395_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1497_ (.I(_0406_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1498_ (.I(net45),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1499_ (.I(_0427_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1500_ (.A1(_0362_),
    .A2(_0384_),
    .A3(_0416_),
    .B(_0438_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1501_ (.A1(_0200_),
    .A2(_0449_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1502_ (.I(_0069_),
    .Z(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1503_ (.I(_0470_),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1504_ (.I(_0135_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1505_ (.I(_0491_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1506_ (.A1(_0481_),
    .A2(_0502_),
    .B(_0438_),
    .C(_0384_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1507_ (.A1(_0200_),
    .A2(_0513_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1508_ (.A1(_0221_),
    .A2(_0341_),
    .B(_0459_),
    .C(_0522_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1509_ (.I(_0533_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1510_ (.A1(_0167_),
    .A2(_0544_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1511_ (.I(_0554_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1512_ (.I(\p_shaping_I.bit_in_1 ),
    .Z(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1513_ (.I(_0570_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1514_ (.I(_0578_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1515_ (.I(_1400_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1516_ (.I(_0592_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1517_ (.I(\p_shaping_I.bit_in ),
    .Z(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1518_ (.I(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1519_ (.I(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1520_ (.I(net48),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1521_ (.A1(\p_shaping_I.ctl_1 ),
    .A2(net57),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1522_ (.A1(_0603_),
    .A2(_0604_),
    .B(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1523_ (.A1(_0599_),
    .A2(_0606_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1524_ (.A1(_0586_),
    .A2(_0599_),
    .B(_0607_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1525_ (.I(\p_shaping_Q.bit_in_1 ),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1526_ (.I(_0608_),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1527_ (.I(\Reg_Delay_Q.Out ),
    .ZN(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1528_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1529_ (.I(_0611_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1530_ (.A1(net48),
    .A2(\p_shaping_Q.ctl_1 ),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1531_ (.A1(_0604_),
    .A2(_0612_),
    .B(_0613_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1532_ (.A1(_0554_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1533_ (.A1(_0609_),
    .A2(_0554_),
    .B(_0615_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1534_ (.A1(_0604_),
    .A2(_0599_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1535_ (.I(_0616_),
    .Z(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1536_ (.A1(_0604_),
    .A2(_0554_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1537_ (.I(_0617_),
    .Z(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1538_ (.I(_0200_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1539_ (.I(_0618_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1540_ (.I(_0091_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1541_ (.I(_0620_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1542_ (.I(_0621_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1543_ (.I(net46),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1544_ (.I(_0623_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1545_ (.I(_0624_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1546_ (.I(_0124_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1547_ (.I(_0626_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1548_ (.I(_0627_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1549_ (.A1(_0625_),
    .A2(_0628_),
    .ZN(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1550_ (.I(_0623_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1551_ (.A1(_0351_),
    .A2(_0630_),
    .B(_0406_),
    .ZN(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1552_ (.I(_0058_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1553_ (.A1(_0632_),
    .A2(_0308_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1554_ (.A1(_1432_),
    .A2(_0135_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1555_ (.A1(_0351_),
    .A2(_0627_),
    .B(_0634_),
    .C(_0254_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1556_ (.A1(_0622_),
    .A2(_0629_),
    .A3(_0631_),
    .B1(_0633_),
    .B2(_0635_),
    .ZN(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1557_ (.A1(_1443_),
    .A2(_0491_),
    .B(_0254_),
    .ZN(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1558_ (.I(_0637_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1559_ (.A1(net45),
    .A2(net44),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1560_ (.I(_0639_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1561_ (.A1(_0638_),
    .A2(_0640_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1562_ (.A1(_0618_),
    .A2(_0449_),
    .B(_0641_),
    .ZN(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1563_ (.I(net39),
    .ZN(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1564_ (.I(_0643_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1565_ (.I(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1566_ (.A1(_0243_),
    .A2(_0628_),
    .B(_0645_),
    .ZN(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1567_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1568_ (.I(_0124_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1569_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1570_ (.I(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1571_ (.A1(_0058_),
    .A2(net46),
    .ZN(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1572_ (.I(_0651_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1573_ (.I(_0652_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1574_ (.A1(_0362_),
    .A2(_0625_),
    .A3(_0416_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1575_ (.I(_0621_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1576_ (.A1(_0650_),
    .A2(_0653_),
    .B(_0654_),
    .C(_0655_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1577_ (.I(net45),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1578_ (.I(_0657_),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1579_ (.I(net44),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1580_ (.A1(_0658_),
    .A2(_0659_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1581_ (.I(_0660_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1582_ (.A1(_0647_),
    .A2(_0656_),
    .B(_0661_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1583_ (.A1(_0619_),
    .A2(_0636_),
    .B(_0642_),
    .C(_0662_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1584_ (.I(_0663_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1585_ (.I(\p_shaping_Q.counter[1] ),
    .Z(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1586_ (.I(_0665_),
    .Z(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1587_ (.I(_0178_),
    .Z(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1588_ (.I(_0667_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1589_ (.I(net44),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1590_ (.I(_0669_),
    .Z(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1591_ (.A1(_0069_),
    .A2(_0308_),
    .A3(_0102_),
    .A4(_0648_),
    .Z(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1592_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1593_ (.A1(_0670_),
    .A2(_0672_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1594_ (.I(_0624_),
    .Z(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1595_ (.I(_0674_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1596_ (.A1(_0632_),
    .A2(_0308_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1597_ (.A1(_0470_),
    .A2(_0145_),
    .B(_0373_),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _1598_ (.A1(_0675_),
    .A2(_0297_),
    .B1(_0676_),
    .B2(_0677_),
    .C(_0670_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1599_ (.A1(_0673_),
    .A2(_0678_),
    .Z(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1600_ (.I(_0628_),
    .Z(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1601_ (.A1(_0675_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1602_ (.A1(_0351_),
    .A2(_0406_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1603_ (.I(_0682_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1604_ (.A1(_0080_),
    .A2(_0674_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1605_ (.A1(_0650_),
    .A2(_0684_),
    .B(_0655_),
    .ZN(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1606_ (.A1(_0681_),
    .A2(_0683_),
    .A3(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1607_ (.I(_0640_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1608_ (.I(_0395_),
    .Z(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1609_ (.A1(_0232_),
    .A2(_0688_),
    .ZN(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1610_ (.A1(_0265_),
    .A2(_0689_),
    .A3(_0653_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1611_ (.A1(_0687_),
    .A2(_0690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1612_ (.I(_0643_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1613_ (.I(_0692_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1614_ (.I(_0693_),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1615_ (.I(_0626_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1616_ (.I(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1617_ (.A1(_0362_),
    .A2(_0696_),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _1618_ (.I0(_0694_),
    .I1(_0647_),
    .S(_0697_),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _1619_ (.A1(_0668_),
    .A2(_0679_),
    .B1(_0686_),
    .B2(_0691_),
    .C1(_0698_),
    .C2(_0673_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1620_ (.A1(_0620_),
    .A2(_0427_),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1621_ (.A1(_0669_),
    .A2(_0700_),
    .ZN(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1622_ (.I(net37),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1623_ (.A1(_0702_),
    .A2(_0623_),
    .B(_0124_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1624_ (.A1(_0620_),
    .A2(_0658_),
    .A3(_0669_),
    .A4(_0703_),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1625_ (.A1(_0232_),
    .A2(_0624_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1626_ (.A1(_0701_),
    .A2(_0704_),
    .B(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1627_ (.A1(_0658_),
    .A2(_0189_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1628_ (.A1(_0702_),
    .A2(_1432_),
    .Z(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1629_ (.A1(_0632_),
    .A2(_0648_),
    .B(_0102_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1630_ (.A1(_0491_),
    .A2(_0708_),
    .B(_0709_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1631_ (.A1(_0695_),
    .A2(_0676_),
    .B(_0373_),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1632_ (.A1(_0427_),
    .A2(_0189_),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1633_ (.A1(_0632_),
    .A2(_0648_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1634_ (.A1(_0630_),
    .A2(_0713_),
    .B(_0254_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1635_ (.A1(_0707_),
    .A2(_0710_),
    .A3(_0711_),
    .B1(_0712_),
    .B2(_0714_),
    .ZN(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1636_ (.A1(_0706_),
    .A2(_0715_),
    .Z(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1637_ (.I(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1638_ (.A1(_0666_),
    .A2(_0699_),
    .A3(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1639_ (.I(_0665_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1640_ (.A1(_0706_),
    .A2(_0715_),
    .ZN(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1641_ (.I(\p_shaping_Q.counter[1] ),
    .Z(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1642_ (.A1(_0721_),
    .A2(\p_shaping_Q.counter[0] ),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1643_ (.I(_0722_),
    .Z(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1644_ (.I(_0659_),
    .Z(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1645_ (.I(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1646_ (.A1(_0725_),
    .A2(_0672_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1647_ (.I(_0702_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1648_ (.I(_0727_),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1649_ (.I(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1650_ (.I(_0655_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1651_ (.I(_0650_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1652_ (.A1(_0729_),
    .A2(_0730_),
    .A3(_0731_),
    .ZN(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1653_ (.A1(_0647_),
    .A2(_0697_),
    .B(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1654_ (.A1(_0646_),
    .A2(_0629_),
    .A3(_0631_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1655_ (.A1(_0687_),
    .A2(_0690_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1656_ (.A1(_0673_),
    .A2(_0678_),
    .B(_0668_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1657_ (.A1(_0726_),
    .A2(_0733_),
    .B1(_0734_),
    .B2(_0735_),
    .C(_0736_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1658_ (.A1(_0719_),
    .A2(_0720_),
    .B1(_0723_),
    .B2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1659_ (.A1(_0718_),
    .A2(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1660_ (.A1(_0664_),
    .A2(_0739_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1661_ (.I(_0740_),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1662_ (.A1(_0664_),
    .A2(_0739_),
    .ZN(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1663_ (.A1(_0718_),
    .A2(_0741_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1664_ (.I(_0723_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1665_ (.I(_0721_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1666_ (.I(\p_shaping_Q.bit_in_2 ),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1667_ (.I(_0730_),
    .Z(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1668_ (.I(_0630_),
    .Z(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1669_ (.A1(_0470_),
    .A2(_0747_),
    .B(_0695_),
    .ZN(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1670_ (.I(_0297_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1671_ (.I(_0705_),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1672_ (.A1(_0749_),
    .A2(_0750_),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1673_ (.A1(_0746_),
    .A2(_0748_),
    .B(_0751_),
    .ZN(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1674_ (.I(_0667_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1675_ (.A1(_0753_),
    .A2(_0672_),
    .B(_0619_),
    .ZN(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1676_ (.I(_0727_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1677_ (.I(_0755_),
    .Z(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1678_ (.I(_0731_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1679_ (.A1(_0756_),
    .A2(_0757_),
    .B(_0638_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1680_ (.A1(_0502_),
    .A2(_0708_),
    .B(_0384_),
    .ZN(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1681_ (.I(_0657_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1682_ (.I(_0760_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1683_ (.I(_0761_),
    .Z(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1684_ (.A1(_0758_),
    .A2(_0759_),
    .B(_0762_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1685_ (.I(_0724_),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1686_ (.I(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1687_ (.I(_0644_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1688_ (.A1(_0766_),
    .A2(_0658_),
    .A3(_0652_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1689_ (.A1(_0765_),
    .A2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1690_ (.A1(_0752_),
    .A2(_0754_),
    .B1(_0763_),
    .B2(_0768_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1691_ (.A1(_0745_),
    .A2(_0720_),
    .B(_0769_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1692_ (.I(\p_shaping_Q.bit_in_2 ),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1693_ (.I(_0771_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1694_ (.A1(_0695_),
    .A2(_0652_),
    .B(_0692_),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1695_ (.A1(_0635_),
    .A2(_0773_),
    .B(_0178_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1696_ (.A1(_0727_),
    .A2(_1443_),
    .B(_0620_),
    .C(_0688_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1697_ (.A1(_0297_),
    .A2(_0705_),
    .B(_0775_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1698_ (.A1(_0427_),
    .A2(_0671_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1699_ (.A1(_0659_),
    .A2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1700_ (.A1(_0670_),
    .A2(_0774_),
    .A3(_0767_),
    .B1(_0776_),
    .B2(_0778_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1701_ (.A1(_0772_),
    .A2(_0717_),
    .A3(_0779_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1702_ (.A1(_0744_),
    .A2(_0770_),
    .A3(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1703_ (.I(_0764_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1704_ (.I(_0782_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1705_ (.I(_0761_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1706_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1707_ (.A1(_0755_),
    .A2(_0649_),
    .B(_0319_),
    .ZN(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _1708_ (.A1(_0629_),
    .A2(_0631_),
    .B1(_0786_),
    .B2(_0746_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1709_ (.A1(_0749_),
    .A2(_0633_),
    .Z(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1710_ (.A1(_0668_),
    .A2(_0788_),
    .Z(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _1711_ (.A1(_0785_),
    .A2(_0787_),
    .B(_0789_),
    .C(_0732_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1712_ (.I(_0694_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1713_ (.A1(_0362_),
    .A2(_0036_),
    .B(_0416_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1714_ (.I(_0792_),
    .Z(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1715_ (.A1(_0680_),
    .A2(_0653_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1716_ (.I(_0794_),
    .Z(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _1717_ (.A1(_0319_),
    .A2(_0649_),
    .Z(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1718_ (.I(_0438_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1719_ (.A1(_0756_),
    .A2(_0796_),
    .B(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1720_ (.A1(_0791_),
    .A2(_0793_),
    .B(_0795_),
    .C(_0798_),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1721_ (.A1(_0764_),
    .A2(_0449_),
    .Z(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1722_ (.A1(_0799_),
    .A2(_0800_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1723_ (.A1(_0783_),
    .A2(_0790_),
    .B(_0801_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1724_ (.I(\p_shaping_Q.bit_in_1 ),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1725_ (.A1(_0803_),
    .A2(_0737_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1726_ (.A1(_0802_),
    .A2(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1727_ (.A1(_0781_),
    .A2(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1728_ (.A1(_0612_),
    .A2(_0664_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1729_ (.A1(_0481_),
    .A2(_0502_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1730_ (.I(_0080_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1731_ (.A1(_0623_),
    .A2(_0395_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1732_ (.A1(_0809_),
    .A2(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1733_ (.I(_0747_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1734_ (.A1(_0809_),
    .A2(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1735_ (.I(_0766_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _1736_ (.I0(_0808_),
    .I1(_0654_),
    .I2(_0811_),
    .I3(_0813_),
    .S0(_0760_),
    .S1(_0814_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1737_ (.I(_0703_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1738_ (.I(_0816_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1739_ (.I(_0773_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1740_ (.A1(_0817_),
    .A2(_0818_),
    .B(_0221_),
    .C(_0635_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1741_ (.A1(_0764_),
    .A2(_0815_),
    .B(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1742_ (.A1(_0807_),
    .A2(_0820_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1743_ (.A1(_0743_),
    .A2(_0806_),
    .A3(_0821_),
    .Z(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1744_ (.I(_0722_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1745_ (.I(_0823_),
    .Z(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1746_ (.A1(_0824_),
    .A2(_0806_),
    .B(_0821_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1747_ (.A1(_0742_),
    .A2(_0822_),
    .A3(_0825_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1748_ (.I(_0721_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1749_ (.I(_0827_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1750_ (.A1(_0828_),
    .A2(_0770_),
    .A3(_0780_),
    .A4(_0805_),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1751_ (.A1(_0743_),
    .A2(_0806_),
    .A3(_0821_),
    .B(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1752_ (.A1(_0720_),
    .A2(_0769_),
    .B(_0745_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1753_ (.A1(_0625_),
    .A2(_0287_),
    .B1(_0631_),
    .B2(_0645_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1754_ (.A1(_0627_),
    .A2(_0633_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1755_ (.A1(_0702_),
    .A2(_1432_),
    .A3(_0395_),
    .Z(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _1756_ (.A1(_0834_),
    .A2(_0816_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1757_ (.A1(_0657_),
    .A2(_0669_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1758_ (.A1(_0621_),
    .A2(_0833_),
    .B1(_0835_),
    .B2(_0775_),
    .C(_0836_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1759_ (.A1(_0624_),
    .A2(_0688_),
    .ZN(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1760_ (.A1(_0766_),
    .A2(_0838_),
    .ZN(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1761_ (.A1(_0728_),
    .A2(_0319_),
    .A3(_0287_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1762_ (.A1(_0839_),
    .A2(_0639_),
    .A3(_0748_),
    .A4(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1763_ (.A1(_0660_),
    .A2(_0832_),
    .B(_0837_),
    .C(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1764_ (.A1(_0831_),
    .A2(_0842_),
    .Z(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1765_ (.A1(_0243_),
    .A2(_0838_),
    .B(_0645_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1766_ (.I(_0243_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1767_ (.A1(_0845_),
    .A2(_0810_),
    .B(_0730_),
    .ZN(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1768_ (.A1(_0786_),
    .A2(_0844_),
    .B(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1769_ (.I(_0689_),
    .Z(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1770_ (.A1(_0812_),
    .A2(_0384_),
    .A3(_0848_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1771_ (.I(_0836_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1772_ (.I(_0850_),
    .Z(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1773_ (.I(_0747_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1774_ (.I(_0766_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1775_ (.I(_0145_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1776_ (.A1(_0809_),
    .A2(_0852_),
    .A3(_0853_),
    .A4(_0854_),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1777_ (.A1(_0851_),
    .A2(_0855_),
    .Z(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1778_ (.I(_0036_),
    .Z(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1779_ (.A1(_0857_),
    .A2(_0724_),
    .A3(_0156_),
    .ZN(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1780_ (.A1(_0818_),
    .A2(_0846_),
    .B1(_0858_),
    .B2(_0661_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1781_ (.A1(_0687_),
    .A2(_0847_),
    .B1(_0849_),
    .B2(_0856_),
    .C(_0859_),
    .ZN(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1782_ (.A1(_0610_),
    .A2(_0613_),
    .Z(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1783_ (.A1(_0167_),
    .A2(_0544_),
    .A3(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1784_ (.I(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1785_ (.A1(_0728_),
    .A2(_0649_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1786_ (.I(_0864_),
    .Z(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1787_ (.I(_0853_),
    .Z(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1788_ (.A1(_0852_),
    .A2(_0865_),
    .B(_0796_),
    .C(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1789_ (.A1(_0809_),
    .A2(_0696_),
    .B(_0852_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1790_ (.A1(_0865_),
    .A2(_0868_),
    .B(_0784_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1791_ (.A1(_0797_),
    .A2(_0788_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1792_ (.A1(_0470_),
    .A2(_0692_),
    .A3(_0627_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1793_ (.A1(_0867_),
    .A2(_0869_),
    .B(_0870_),
    .C(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _1794_ (.A1(_0619_),
    .A2(_0872_),
    .B1(_0799_),
    .B2(_0800_),
    .C(_0699_),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1795_ (.I(_0803_),
    .Z(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1796_ (.A1(_0860_),
    .A2(_0863_),
    .B1(_0873_),
    .B2(_0874_),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1797_ (.A1(_0755_),
    .A2(_0796_),
    .B(_0265_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1798_ (.I(_0634_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1799_ (.A1(_0729_),
    .A2(_0877_),
    .B(_0853_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1800_ (.A1(_0868_),
    .A2(_0876_),
    .B(_0878_),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1801_ (.A1(_0625_),
    .A2(_0659_),
    .A3(_0156_),
    .Z(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1802_ (.A1(_0759_),
    .A2(_0878_),
    .B1(_0880_),
    .B2(_0210_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1803_ (.A1(_0850_),
    .A2(_0849_),
    .A3(_0855_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1804_ (.A1(_0707_),
    .A2(_0879_),
    .B(_0881_),
    .C(_0882_),
    .ZN(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1805_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1806_ (.A1(_0167_),
    .A2(_0533_),
    .A3(_0861_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1807_ (.I(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _1808_ (.A1(_0765_),
    .A2(_0790_),
    .B(_0801_),
    .C(_0737_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _1809_ (.A1(_0609_),
    .A2(_0884_),
    .A3(_0886_),
    .A4(_0887_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1810_ (.A1(_0666_),
    .A2(_0843_),
    .B1(_0875_),
    .B2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1811_ (.A1(_0666_),
    .A2(_0843_),
    .A3(_0875_),
    .A4(_0888_),
    .Z(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1812_ (.A1(_0664_),
    .A2(_0820_),
    .B(_0611_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1813_ (.A1(_0833_),
    .A2(_0876_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1814_ (.A1(_0265_),
    .A2(_0684_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1815_ (.A1(_0622_),
    .A2(_0680_),
    .B(_0667_),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1816_ (.A1(_0618_),
    .A2(_0893_),
    .A3(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1817_ (.A1(_0047_),
    .A2(_0694_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1818_ (.A1(_0865_),
    .A2(_0896_),
    .B(_0714_),
    .C(_0210_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1819_ (.A1(_0845_),
    .A2(_0680_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1820_ (.I(_0626_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1821_ (.A1(_0674_),
    .A2(_0899_),
    .B(_0113_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1822_ (.A1(_0898_),
    .A2(_0900_),
    .B(_0794_),
    .C(_0850_),
    .ZN(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1823_ (.A1(_0892_),
    .A2(_0895_),
    .B(_0897_),
    .C(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1824_ (.A1(_0891_),
    .A2(_0902_),
    .Z(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1825_ (.A1(_0743_),
    .A2(_0889_),
    .A3(_0890_),
    .A4(_0903_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1826_ (.A1(_0824_),
    .A2(_0889_),
    .A3(_0890_),
    .B(_0903_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1827_ (.A1(_0830_),
    .A2(_0904_),
    .A3(_0905_),
    .Z(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1828_ (.A1(_0904_),
    .A2(_0905_),
    .B(_0830_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1829_ (.A1(_0906_),
    .A2(_0907_),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1830_ (.A1(_0826_),
    .A2(_0908_),
    .Z(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1831_ (.I(_0909_),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1832_ (.A1(_0828_),
    .A2(_0843_),
    .A3(_0875_),
    .A4(_0888_),
    .ZN(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1833_ (.A1(_0824_),
    .A2(_0889_),
    .A3(_0903_),
    .B(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1834_ (.A1(_0232_),
    .A2(_0810_),
    .B(_0644_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1835_ (.A1(_0688_),
    .A2(_0651_),
    .B(_0810_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1836_ (.A1(_0912_),
    .A2(_0913_),
    .Z(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1837_ (.A1(_0728_),
    .A2(_1443_),
    .B(_0644_),
    .C(_0406_),
    .ZN(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1838_ (.A1(_0871_),
    .A2(_0915_),
    .B(_0705_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1839_ (.A1(_0080_),
    .A2(_0899_),
    .B(_0838_),
    .C(_0373_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1840_ (.A1(_0864_),
    .A2(_0917_),
    .B(_0836_),
    .ZN(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1841_ (.A1(_0630_),
    .A2(_0491_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1842_ (.A1(_0692_),
    .A2(_0689_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1843_ (.A1(_0919_),
    .A2(_0920_),
    .B1(_0835_),
    .B2(_0637_),
    .C(_0639_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _1844_ (.A1(_0660_),
    .A2(_0914_),
    .B1(_0916_),
    .B2(_0918_),
    .C(_0921_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1845_ (.A1(_0717_),
    .A2(_0779_),
    .A3(_0842_),
    .B(_0771_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1846_ (.A1(_0922_),
    .A2(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1847_ (.A1(_0628_),
    .A2(_0652_),
    .B(_0682_),
    .C(_0621_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1848_ (.A1(_0760_),
    .A2(_0871_),
    .A3(_0925_),
    .A4(_0915_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1849_ (.A1(_0760_),
    .A2(_0330_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1850_ (.A1(_0714_),
    .A2(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1851_ (.A1(_0729_),
    .A2(_0502_),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1852_ (.A1(_0696_),
    .A2(_0708_),
    .B(_0693_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1853_ (.A1(_0729_),
    .A2(_0812_),
    .A3(_0854_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1854_ (.A1(_0814_),
    .A2(_0929_),
    .B1(_0930_),
    .B2(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _1855_ (.A1(_0724_),
    .A2(_0926_),
    .A3(_0928_),
    .B1(_0778_),
    .B2(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1856_ (.A1(_0862_),
    .A2(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1857_ (.A1(_0609_),
    .A2(_0884_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1858_ (.A1(_0874_),
    .A2(_0873_),
    .B(_0934_),
    .C(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1859_ (.A1(_0884_),
    .A2(_0887_),
    .B1(_0933_),
    .B2(_0863_),
    .C(_0609_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1860_ (.A1(_0827_),
    .A2(_0924_),
    .B1(_0936_),
    .B2(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1861_ (.A1(_0827_),
    .A2(_0924_),
    .A3(_0936_),
    .A4(_0937_),
    .Z(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1862_ (.A1(_0823_),
    .A2(_0938_),
    .A3(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1863_ (.A1(_0663_),
    .A2(_0820_),
    .A3(_0902_),
    .Z(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1864_ (.A1(_0611_),
    .A2(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1865_ (.I(_0899_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1866_ (.A1(_0845_),
    .A2(_0047_),
    .A3(_0943_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _1867_ (.A1(_0747_),
    .A2(_0416_),
    .B(_0693_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1868_ (.A1(_0866_),
    .A2(_0676_),
    .B1(_0944_),
    .B2(_0945_),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1869_ (.A1(_0675_),
    .A2(_0848_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1870_ (.I(_0655_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1871_ (.I(_0707_),
    .Z(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _1872_ (.A1(_0330_),
    .A2(_0929_),
    .B1(_0947_),
    .B2(_0948_),
    .C(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1873_ (.A1(_0851_),
    .A2(_0946_),
    .B(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1874_ (.I(_0653_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1875_ (.I(_0622_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1876_ (.A1(_0952_),
    .A2(_0638_),
    .B1(_0795_),
    .B2(_0953_),
    .C(_0221_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1877_ (.A1(_0858_),
    .A2(_0951_),
    .A3(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1878_ (.A1(_0942_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1879_ (.A1(_0940_),
    .A2(_0956_),
    .Z(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1880_ (.A1(_0826_),
    .A2(_0908_),
    .B(_0906_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1881_ (.A1(_0911_),
    .A2(_0957_),
    .A3(_0958_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1882_ (.I(_0959_),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1883_ (.A1(_0823_),
    .A2(_0938_),
    .A3(_0939_),
    .A4(_0956_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1884_ (.A1(_0939_),
    .A2(_0960_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1885_ (.I(_0722_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1886_ (.A1(_0716_),
    .A2(_0779_),
    .A3(_0842_),
    .A4(_0922_),
    .Z(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1887_ (.A1(_0690_),
    .A2(_0818_),
    .B(_0660_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1888_ (.A1(_0178_),
    .A2(_0677_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1889_ (.A1(_0893_),
    .A2(_0965_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1890_ (.A1(_0674_),
    .A2(_0899_),
    .B(_0755_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1891_ (.A1(_0786_),
    .A2(_0844_),
    .B1(_0900_),
    .B2(_0967_),
    .C(_0438_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1892_ (.A1(_0966_),
    .A2(_0968_),
    .B(_0670_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1893_ (.A1(_0964_),
    .A2(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1894_ (.A1(_0772_),
    .A2(_0963_),
    .B(_0970_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _1895_ (.A1(_0717_),
    .A2(_0779_),
    .A3(_0842_),
    .A4(_0922_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1896_ (.A1(_0964_),
    .A2(_0969_),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1897_ (.A1(_0745_),
    .A2(_0972_),
    .A3(_0973_),
    .B(_0721_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1898_ (.A1(_0884_),
    .A2(_0933_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1899_ (.A1(_0852_),
    .A2(_0732_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1900_ (.A1(_0756_),
    .A2(_0857_),
    .B(_0712_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1901_ (.A1(_0746_),
    .A2(_0683_),
    .A3(_0848_),
    .ZN(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1902_ (.A1(_0276_),
    .A2(_0949_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1903_ (.A1(_0976_),
    .A2(_0977_),
    .B1(_0978_),
    .B2(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1904_ (.I(_0845_),
    .Z(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1905_ (.A1(_0981_),
    .A2(_0838_),
    .B(_0948_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1906_ (.A1(_0683_),
    .A2(_0793_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1907_ (.A1(_0786_),
    .A2(_0982_),
    .B(_0983_),
    .C(_0784_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1908_ (.A1(_0754_),
    .A2(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1909_ (.A1(_0885_),
    .A2(_0980_),
    .A3(_0985_),
    .Z(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1910_ (.A1(_0873_),
    .A2(_0975_),
    .B(_0986_),
    .C(_0803_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1911_ (.I(_0608_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1912_ (.A1(_0731_),
    .A2(_0952_),
    .B(_0948_),
    .ZN(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1913_ (.A1(_0989_),
    .A2(_0944_),
    .B(_0647_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1914_ (.A1(_0785_),
    .A2(_0871_),
    .A3(_0925_),
    .A4(_0915_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1915_ (.A1(_0714_),
    .A2(_0927_),
    .B(_0725_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1916_ (.A1(_0754_),
    .A2(_0990_),
    .B1(_0991_),
    .B2(_0992_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _1917_ (.A1(_0860_),
    .A2(_0993_),
    .B(\p_shaping_Q.bit_in_1 ),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1918_ (.A1(_0886_),
    .A2(_0980_),
    .A3(_0985_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _1919_ (.A1(_0988_),
    .A2(_0887_),
    .B(_0994_),
    .C(_0995_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _1920_ (.A1(_0971_),
    .A2(_0974_),
    .B1(_0987_),
    .B2(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1921_ (.A1(_0971_),
    .A2(_0974_),
    .A3(_0987_),
    .A4(_0996_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1922_ (.A1(_0962_),
    .A2(_0997_),
    .A3(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1923_ (.A1(_0981_),
    .A2(_0791_),
    .A3(_0919_),
    .B(_0839_),
    .ZN(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1924_ (.A1(_0981_),
    .A2(_0965_),
    .B1(_1000_),
    .B2(_0753_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1925_ (.I(_0221_),
    .Z(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1926_ (.A1(_0683_),
    .A2(_0877_),
    .A3(_0793_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1927_ (.A1(_0953_),
    .A2(_1003_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1928_ (.A1(_0791_),
    .A2(_0684_),
    .A3(_0877_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1929_ (.A1(_1002_),
    .A2(_1004_),
    .A3(_1005_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1930_ (.A1(_0782_),
    .A2(_1001_),
    .B(_1006_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1931_ (.A1(_0941_),
    .A2(_0955_),
    .B(_0611_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1932_ (.A1(_1007_),
    .A2(_1008_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1933_ (.A1(_0999_),
    .A2(_1009_),
    .Z(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1934_ (.A1(_0961_),
    .A2(_1010_),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1935_ (.I(_0911_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1936_ (.A1(_1012_),
    .A2(_0957_),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1937_ (.A1(_0742_),
    .A2(_0822_),
    .A3(_0825_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1938_ (.A1(_0830_),
    .A2(_0904_),
    .A3(_0905_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _1939_ (.A1(_1014_),
    .A2(_0907_),
    .B1(_1012_),
    .B2(_0957_),
    .C(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1940_ (.A1(_1013_),
    .A2(_1016_),
    .Z(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _1941_ (.A1(_1011_),
    .A2(_1017_),
    .Z(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1942_ (.I(_1018_),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1943_ (.A1(_0962_),
    .A2(_0997_),
    .Z(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1944_ (.A1(_0971_),
    .A2(_0974_),
    .A3(_0987_),
    .A4(_0996_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1945_ (.A1(_1019_),
    .A2(_1009_),
    .B(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1946_ (.A1(_0808_),
    .A2(_0750_),
    .A3(_0920_),
    .B(_0690_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1947_ (.A1(_0851_),
    .A2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1948_ (.A1(_0113_),
    .A2(_0834_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1949_ (.A1(_0645_),
    .A2(_0816_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1950_ (.A1(_1024_),
    .A2(_1025_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1951_ (.A1(_0661_),
    .A2(_1026_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1952_ (.A1(_0734_),
    .A2(_0945_),
    .B(_0640_),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1953_ (.A1(_1023_),
    .A2(_1027_),
    .A3(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1954_ (.A1(_0963_),
    .A2(_0970_),
    .B(_1029_),
    .C(_0772_),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1955_ (.A1(_1023_),
    .A2(_1027_),
    .A3(_1028_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1956_ (.A1(_0964_),
    .A2(_0969_),
    .B(_0772_),
    .ZN(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _1957_ (.A1(_0745_),
    .A2(_0972_),
    .B(_1031_),
    .C(_1032_),
    .ZN(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1958_ (.A1(_0665_),
    .A2(_1030_),
    .A3(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1959_ (.A1(_0813_),
    .A2(_0876_),
    .B(_0945_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _1960_ (.A1(_0675_),
    .A2(_0814_),
    .A3(_0713_),
    .ZN(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1961_ (.A1(_0814_),
    .A2(_0817_),
    .Z(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1962_ (.A1(_1036_),
    .A2(_1037_),
    .B(_0850_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1963_ (.A1(_0853_),
    .A2(_0816_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1964_ (.A1(_0640_),
    .A2(_0849_),
    .A3(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1965_ (.A1(_0854_),
    .A2(_0750_),
    .B(_0693_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1966_ (.A1(_0481_),
    .A2(_0812_),
    .B(_0696_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _1967_ (.A1(_0694_),
    .A2(_0877_),
    .B1(_1041_),
    .B2(_1042_),
    .C(_0210_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _1968_ (.A1(_1035_),
    .A2(_1038_),
    .B(_1040_),
    .C(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1969_ (.A1(_0988_),
    .A2(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1970_ (.A1(_0994_),
    .A2(_1044_),
    .ZN(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _1971_ (.A1(_0883_),
    .A2(_0933_),
    .A3(_1044_),
    .B(_0608_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1972_ (.I(_1047_),
    .Z(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1973_ (.A1(_0862_),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1974_ (.A1(_0863_),
    .A2(_1045_),
    .A3(_1046_),
    .B(_1049_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1975_ (.A1(_1034_),
    .A2(_1050_),
    .Z(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1976_ (.A1(_1034_),
    .A2(_1050_),
    .B(_0723_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1977_ (.A1(_1051_),
    .A2(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1978_ (.I(_0866_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _1979_ (.I(_0797_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1980_ (.A1(_0753_),
    .A2(_0920_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _1981_ (.A1(_1054_),
    .A2(_0757_),
    .A3(_1055_),
    .B1(_0867_),
    .B2(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1982_ (.I(_0708_),
    .Z(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1983_ (.A1(_0650_),
    .A2(_1058_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1984_ (.A1(_0668_),
    .A2(_0749_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1985_ (.A1(_0839_),
    .A2(_1059_),
    .B(_1060_),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1986_ (.A1(_0673_),
    .A2(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _1987_ (.A1(_0765_),
    .A2(_1057_),
    .B(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1988_ (.I(\Reg_Delay_Q.Out ),
    .Z(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _1989_ (.A1(_0941_),
    .A2(_0955_),
    .A3(_1007_),
    .ZN(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1990_ (.A1(_1064_),
    .A2(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1991_ (.A1(_1063_),
    .A2(_1066_),
    .ZN(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _1992_ (.A1(_1021_),
    .A2(_1053_),
    .A3(_1067_),
    .Z(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1993_ (.A1(_0961_),
    .A2(_1010_),
    .ZN(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1994_ (.A1(_1011_),
    .A2(_1017_),
    .B(_1069_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _1995_ (.A1(_1068_),
    .A2(_1070_),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1996_ (.I(_1071_),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _1997_ (.A1(_1034_),
    .A2(_1050_),
    .Z(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1998_ (.A1(_1051_),
    .A2(_1052_),
    .A3(_1067_),
    .Z(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _1999_ (.A1(_1072_),
    .A2(_1073_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2000_ (.A1(_0330_),
    .A2(_0833_),
    .ZN(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2001_ (.A1(_0481_),
    .A2(_0036_),
    .A3(_0854_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _2002_ (.A1(_0761_),
    .A2(_0796_),
    .A3(_0713_),
    .A4(_1076_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2003_ (.A1(_0622_),
    .A2(_0761_),
    .A3(_0898_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2004_ (.A1(_1075_),
    .A2(_1078_),
    .B(_1077_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2005_ (.A1(_1075_),
    .A2(_1077_),
    .B(_1079_),
    .C(_0725_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2006_ (.A1(_1002_),
    .A2(_1024_),
    .B(_1080_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2007_ (.A1(_0963_),
    .A2(_0970_),
    .A3(_1029_),
    .B(_0771_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2008_ (.A1(_1081_),
    .A2(_1082_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2009_ (.A1(_0885_),
    .A2(_1047_),
    .Z(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2010_ (.A1(_0656_),
    .A2(_0947_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2011_ (.A1(_0785_),
    .A2(_1085_),
    .B(_0619_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2012_ (.A1(_0047_),
    .A2(_0730_),
    .A3(_0943_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2013_ (.A1(_0667_),
    .A2(_0792_),
    .A3(_0748_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2014_ (.A1(_0797_),
    .A2(_1059_),
    .A3(_0900_),
    .B1(_1088_),
    .B2(_1087_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2015_ (.A1(_1087_),
    .A2(_1088_),
    .B(_1089_),
    .C(_0725_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2016_ (.A1(_1086_),
    .A2(_1090_),
    .Z(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2017_ (.I0(_1047_),
    .I1(_1084_),
    .S(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2018_ (.A1(_0744_),
    .A2(_1083_),
    .B(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2019_ (.A1(_0665_),
    .A2(_1083_),
    .A3(_1092_),
    .Z(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2020_ (.A1(_0722_),
    .A2(_1093_),
    .A3(_1094_),
    .Z(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2021_ (.A1(_1063_),
    .A2(_1065_),
    .B(\Reg_Delay_Q.Out ),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2022_ (.A1(_0757_),
    .A2(_0952_),
    .B(_0709_),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2023_ (.A1(_1056_),
    .A2(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2024_ (.A1(_0783_),
    .A2(_1060_),
    .A3(_1098_),
    .B1(_0661_),
    .B2(_1035_),
    .ZN(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2025_ (.A1(_1096_),
    .A2(_1099_),
    .ZN(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2026_ (.A1(_1095_),
    .A2(_1100_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2027_ (.A1(_1074_),
    .A2(_1101_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2028_ (.A1(_1013_),
    .A2(_1011_),
    .A3(_1016_),
    .A4(_1068_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2029_ (.A1(_1051_),
    .A2(_1052_),
    .B(_1067_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2030_ (.A1(_1021_),
    .A2(_1073_),
    .A3(_1104_),
    .ZN(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2031_ (.A1(_1073_),
    .A2(_1104_),
    .B(_1021_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2032_ (.A1(_1069_),
    .A2(_1105_),
    .B(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2033_ (.A1(_1103_),
    .A2(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2034_ (.A1(_1102_),
    .A2(_1108_),
    .Z(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2035_ (.I(_1109_),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2036_ (.A1(_0828_),
    .A2(_1083_),
    .A3(_1092_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2037_ (.A1(_1095_),
    .A2(_1100_),
    .B(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2038_ (.A1(_0731_),
    .A2(_1058_),
    .B(_1076_),
    .C(_0791_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2039_ (.A1(_0681_),
    .A2(_0677_),
    .B(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2040_ (.A1(_0818_),
    .A2(_1059_),
    .B(_0917_),
    .C(_1055_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2041_ (.A1(_1055_),
    .A2(_1113_),
    .B(_1114_),
    .ZN(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2042_ (.A1(_0276_),
    .A2(_0710_),
    .B1(_0880_),
    .B2(_1002_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2043_ (.A1(_0765_),
    .A2(_1115_),
    .B(_1116_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2044_ (.A1(_0994_),
    .A2(_1045_),
    .A3(_1117_),
    .Z(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2045_ (.A1(_0988_),
    .A2(_1117_),
    .B(_0862_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2046_ (.A1(_0868_),
    .A2(_0876_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2047_ (.A1(_0866_),
    .A2(_1076_),
    .Z(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2048_ (.A1(_0929_),
    .A2(_0833_),
    .A3(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2049_ (.A1(_0894_),
    .A2(_1120_),
    .B1(_1122_),
    .B2(_1055_),
    .C(_0782_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2050_ (.A1(_1082_),
    .A2(_1123_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2051_ (.A1(_0873_),
    .A2(_0975_),
    .B(_0803_),
    .C(_0885_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2052_ (.I(_1125_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2053_ (.A1(_1118_),
    .A2(_1119_),
    .B1(_1124_),
    .B2(_0744_),
    .C(_1126_),
    .ZN(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2054_ (.A1(_1118_),
    .A2(_1119_),
    .B(_1125_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2055_ (.I(_1082_),
    .Z(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2056_ (.A1(_1129_),
    .A2(_1123_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2057_ (.A1(_0719_),
    .A2(_1128_),
    .A3(_1130_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2058_ (.A1(_0723_),
    .A2(_1127_),
    .A3(_1131_),
    .ZN(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2059_ (.A1(_0709_),
    .A2(_0712_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2060_ (.A1(_1002_),
    .A2(_0880_),
    .B(_1078_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2061_ (.A1(_0700_),
    .A2(_0835_),
    .B(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2062_ (.A1(_0793_),
    .A2(_1133_),
    .B(_1135_),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2063_ (.A1(_1096_),
    .A2(_1136_),
    .Z(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2064_ (.A1(_1132_),
    .A2(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2065_ (.A1(_1111_),
    .A2(_1138_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2066_ (.A1(_1074_),
    .A2(_1101_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2067_ (.A1(_1102_),
    .A2(_1108_),
    .B(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2068_ (.A1(_1139_),
    .A2(_1141_),
    .ZN(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2069_ (.I(_1142_),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2070_ (.I(_1131_),
    .ZN(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2071_ (.A1(_0824_),
    .A2(_1127_),
    .A3(_1137_),
    .B(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2072_ (.I(_0753_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2073_ (.A1(_0759_),
    .A2(_0795_),
    .B(_0778_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2074_ (.A1(_0757_),
    .A2(_1058_),
    .B(_0865_),
    .C(_0953_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2075_ (.A1(_0948_),
    .A2(_0750_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2076_ (.A1(_0953_),
    .A2(_0848_),
    .B1(_1148_),
    .B2(_0681_),
    .C(_0784_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2077_ (.A1(_0785_),
    .A2(_1147_),
    .B(_1149_),
    .C(_0782_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2078_ (.A1(_1145_),
    .A2(_0638_),
    .A3(_1042_),
    .B1(_1146_),
    .B2(_1150_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2079_ (.I0(_0988_),
    .I1(_1048_),
    .S(_1151_),
    .Z(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2080_ (.A1(_0886_),
    .A2(_1152_),
    .B(_1126_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2081_ (.A1(_0962_),
    .A2(_1153_),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2082_ (.I(\p_shaping_Q.bit_in_2 ),
    .Z(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2083_ (.A1(_0685_),
    .A2(_0795_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2084_ (.A1(_0894_),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2085_ (.I(_0618_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2086_ (.A1(_1158_),
    .A2(_1121_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2087_ (.A1(_0949_),
    .A2(_1159_),
    .ZN(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2088_ (.A1(_0762_),
    .A2(_1039_),
    .B(_1157_),
    .C(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2089_ (.A1(_0777_),
    .A2(_0984_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2090_ (.A1(_1155_),
    .A2(_1162_),
    .B(_1129_),
    .C(_1161_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2091_ (.A1(_1155_),
    .A2(_1161_),
    .B(_1163_),
    .C(_0744_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2092_ (.A1(_1154_),
    .A2(_1164_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2093_ (.A1(_1064_),
    .A2(_0544_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2094_ (.A1(_1063_),
    .A2(_1065_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2095_ (.A1(_0981_),
    .A2(_0945_),
    .B1(_1003_),
    .B2(_1054_),
    .C(_1145_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2096_ (.A1(_1064_),
    .A2(_0544_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2097_ (.A1(_1167_),
    .A2(_1168_),
    .B(_1169_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2098_ (.A1(_1166_),
    .A2(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2099_ (.A1(_1165_),
    .A2(_1171_),
    .Z(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2100_ (.A1(_1144_),
    .A2(_1172_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2101_ (.A1(_1103_),
    .A2(_1107_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2102_ (.A1(_1102_),
    .A2(_1139_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2103_ (.A1(_1111_),
    .A2(_1138_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2104_ (.A1(_1111_),
    .A2(_1138_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2105_ (.A1(_1140_),
    .A2(_1176_),
    .B(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2106_ (.A1(_1174_),
    .A2(_1175_),
    .B(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2107_ (.A1(_1173_),
    .A2(_1179_),
    .Z(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2108_ (.I(_1180_),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2109_ (.A1(_1154_),
    .A2(_1164_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2110_ (.A1(_1165_),
    .A2(_1171_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2111_ (.A1(_1181_),
    .A2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2112_ (.I(_0962_),
    .Z(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2113_ (.A1(_0943_),
    .A2(_1058_),
    .B(_0713_),
    .C(_1054_),
    .ZN(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2114_ (.A1(_0949_),
    .A2(_0685_),
    .A3(_1184_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2115_ (.A1(_0851_),
    .A2(_1039_),
    .B1(_1168_),
    .B2(_0783_),
    .C(_1185_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2116_ (.A1(_1048_),
    .A2(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2117_ (.A1(_0874_),
    .A2(_1186_),
    .B(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2118_ (.A1(_0886_),
    .A2(_1188_),
    .B(_1126_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2119_ (.A1(_0022_),
    .A2(_1189_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2120_ (.A1(_0749_),
    .A2(_1024_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2121_ (.A1(_1191_),
    .A2(_1076_),
    .B(_0762_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2122_ (.A1(_1160_),
    .A2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2123_ (.A1(_1129_),
    .A2(_1193_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2124_ (.A1(_1155_),
    .A2(_1193_),
    .B(_1194_),
    .C(_0827_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2125_ (.A1(_0459_),
    .A2(_0522_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2126_ (.A1(_1158_),
    .A2(_0341_),
    .B(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2127_ (.A1(_1096_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2128_ (.A1(_0612_),
    .A2(_1197_),
    .B(_1198_),
    .ZN(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2129_ (.A1(_1190_),
    .A2(_1195_),
    .A3(_1199_),
    .Z(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2130_ (.A1(_1183_),
    .A2(_1200_),
    .ZN(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2131_ (.A1(_1144_),
    .A2(_1172_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2132_ (.A1(_1173_),
    .A2(_1179_),
    .B(_1202_),
    .ZN(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2133_ (.A1(_1201_),
    .A2(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2134_ (.I(_1204_),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2135_ (.A1(_0746_),
    .A2(_0817_),
    .B(_1060_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2136_ (.A1(_0687_),
    .A2(_1026_),
    .B1(_1205_),
    .B2(_0783_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2137_ (.A1(_1084_),
    .A2(_1206_),
    .B(_0823_),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2138_ (.A1(_1084_),
    .A2(_1206_),
    .B(_1207_),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2139_ (.A1(_1145_),
    .A2(_0672_),
    .B(_1160_),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2140_ (.A1(_1129_),
    .A2(_1209_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2141_ (.A1(_1155_),
    .A2(_1209_),
    .B(_1210_),
    .C(_0666_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2142_ (.A1(_1208_),
    .A2(_1211_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2143_ (.A1(_1064_),
    .A2(_0522_),
    .B1(_1196_),
    .B2(_1096_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2144_ (.A1(_1212_),
    .A2(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2145_ (.A1(_1190_),
    .A2(_1195_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2146_ (.A1(_1190_),
    .A2(_1195_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2147_ (.A1(_1215_),
    .A2(_1199_),
    .B(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2148_ (.A1(_1214_),
    .A2(_1217_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2149_ (.I(_1201_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2150_ (.A1(_1181_),
    .A2(_1182_),
    .B(_1200_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2151_ (.A1(_1202_),
    .A2(_1220_),
    .Z(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2152_ (.A1(_1181_),
    .A2(_1182_),
    .A3(_1200_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2153_ (.A1(_1173_),
    .A2(_1179_),
    .A3(_1219_),
    .B1(_1221_),
    .B2(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2154_ (.A1(_1218_),
    .A2(_1223_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2155_ (.I(_1224_),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2156_ (.A1(_1208_),
    .A2(_1211_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2157_ (.A1(_1212_),
    .A2(_1213_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2158_ (.A1(_1225_),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2159_ (.A1(_0743_),
    .A2(_1126_),
    .Z(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2160_ (.A1(_1145_),
    .A2(_1025_),
    .B(_1158_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2161_ (.A1(_0701_),
    .A2(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2162_ (.A1(_1048_),
    .A2(_1230_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2163_ (.A1(_0874_),
    .A2(_1230_),
    .B(_1231_),
    .C(_0863_),
    .ZN(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2164_ (.A1(_1228_),
    .A2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2165_ (.A1(_1213_),
    .A2(_1233_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2166_ (.A1(_1213_),
    .A2(_1233_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2167_ (.A1(_1234_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2168_ (.A1(_1211_),
    .A2(_1236_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2169_ (.A1(_1227_),
    .A2(_1237_),
    .ZN(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2170_ (.A1(_1214_),
    .A2(_1217_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2171_ (.A1(_1218_),
    .A2(_1223_),
    .B(_1239_),
    .ZN(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2172_ (.A1(_1238_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2173_ (.I(_1241_),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2174_ (.A1(_1218_),
    .A2(_1223_),
    .A3(_1238_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2175_ (.A1(_1225_),
    .A2(_1226_),
    .B(_1237_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2176_ (.A1(_1225_),
    .A2(_1226_),
    .A3(_1237_),
    .B(_1239_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2177_ (.A1(_1243_),
    .A2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2178_ (.A1(_1211_),
    .A2(_1234_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2179_ (.A1(_1235_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2180_ (.A1(_0022_),
    .A2(_1084_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2181_ (.A1(_1242_),
    .A2(_1245_),
    .A3(_1247_),
    .B(_1248_),
    .ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2182_ (.A1(_0822_),
    .A2(_0825_),
    .B(_0742_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2183_ (.A1(_0826_),
    .A2(_1249_),
    .ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2184_ (.I(_1335_),
    .Z(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2185_ (.A1(_1250_),
    .A2(_1280_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2186_ (.I(_1324_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2187_ (.I(_1252_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2188_ (.I(_1379_),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2189_ (.I(_1368_),
    .Z(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2190_ (.A1(_1269_),
    .A2(_1255_),
    .B(_1357_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2191_ (.A1(_1253_),
    .A2(_1254_),
    .B(_1256_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2192_ (.A1(_1251_),
    .A2(_1257_),
    .ZN(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2193_ (.I(net34),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2194_ (.I(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2195_ (.I(_1261_),
    .Z(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2196_ (.I(net30),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2197_ (.I(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2198_ (.I(net32),
    .Z(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2199_ (.I(_1265_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2200_ (.A1(_1264_),
    .A2(_1266_),
    .Z(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2201_ (.I(_1252_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2202_ (.I(_1264_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2203_ (.A1(_1268_),
    .A2(_1270_),
    .A3(_1254_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2204_ (.A1(_1357_),
    .A2(_1302_),
    .ZN(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2205_ (.I(_1272_),
    .Z(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2206_ (.I(_1256_),
    .Z(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2207_ (.A1(_1273_),
    .A2(_1274_),
    .Z(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2208_ (.A1(_1262_),
    .A2(_1267_),
    .A3(_1271_),
    .B(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2209_ (.I(net47),
    .Z(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2210_ (.I(_1277_),
    .Z(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2211_ (.A1(_1259_),
    .A2(_1276_),
    .B(_1278_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _2212_ (.I(net47),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2213_ (.I(_1281_),
    .Z(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2214_ (.A1(_1262_),
    .A2(_1389_),
    .Z(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2215_ (.I(_1346_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2216_ (.I(_1284_),
    .Z(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2217_ (.I(_1285_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2218_ (.I(_1379_),
    .Z(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2219_ (.A1(_1268_),
    .A2(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2220_ (.I(net32),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2221_ (.I(_1289_),
    .Z(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2222_ (.I(_1290_),
    .Z(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2223_ (.I(net31),
    .Z(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2224_ (.A1(_1293_),
    .A2(_1263_),
    .Z(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2225_ (.A1(_1292_),
    .A2(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2226_ (.I(_1346_),
    .Z(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2227_ (.I(_1296_),
    .Z(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2228_ (.I(_1293_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2229_ (.I(_1298_),
    .Z(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2230_ (.I(_1258_),
    .Z(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2231_ (.I(_1300_),
    .Z(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2232_ (.I(_1265_),
    .Z(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2233_ (.A1(_1299_),
    .A2(_1301_),
    .A3(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2234_ (.A1(_1297_),
    .A2(_1304_),
    .Z(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2235_ (.A1(_1286_),
    .A2(_1288_),
    .B1(_1295_),
    .B2(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2236_ (.A1(_1291_),
    .A2(_1261_),
    .ZN(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2237_ (.I(_1307_),
    .Z(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2238_ (.A1(_1282_),
    .A2(_1283_),
    .B1(_1306_),
    .B2(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2239_ (.A1(_1279_),
    .A2(_1309_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2240_ (.I(\p_shaping_I.counter[1] ),
    .Z(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2241_ (.A1(_1311_),
    .A2(\p_shaping_I.counter[0] ),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2242_ (.I(_1312_),
    .Z(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2243_ (.I(_1314_),
    .Z(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2244_ (.A1(_1253_),
    .A2(_1270_),
    .B(_1292_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2245_ (.I(_1266_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2246_ (.I(_1346_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2247_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2248_ (.A1(_1317_),
    .A2(_1251_),
    .B(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2249_ (.I(_1284_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2250_ (.I(_1321_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2251_ (.I(_1368_),
    .Z(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2252_ (.A1(_1298_),
    .A2(_1323_),
    .Z(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2253_ (.A1(_1322_),
    .A2(_1325_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2254_ (.A1(_1293_),
    .A2(_1258_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2255_ (.I(_1327_),
    .Z(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2256_ (.I(_1313_),
    .Z(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2257_ (.A1(_1316_),
    .A2(_1320_),
    .B1(_1326_),
    .B2(_1328_),
    .C(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2258_ (.I(_1357_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2259_ (.I(_1331_),
    .Z(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2260_ (.I(_1267_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2261_ (.I(_1335_),
    .Z(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2262_ (.A1(_1334_),
    .A2(_1270_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2263_ (.A1(_1250_),
    .A2(_1287_),
    .B(_1331_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2264_ (.A1(_1332_),
    .A2(_1333_),
    .B1(_1336_),
    .B2(_1337_),
    .C(_1262_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2265_ (.I(net34),
    .Z(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2266_ (.I(_1293_),
    .Z(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2267_ (.I(net33),
    .Z(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _2268_ (.A1(_1340_),
    .A2(_1300_),
    .A3(_1341_),
    .A4(_1323_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2269_ (.A1(_1339_),
    .A2(_1342_),
    .ZN(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2270_ (.A1(_1277_),
    .A2(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2271_ (.I(_1334_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2272_ (.I(_1285_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2273_ (.I(_1287_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2274_ (.A1(_1347_),
    .A2(_1348_),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2275_ (.I(_1288_),
    .Z(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2276_ (.I(_1289_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2277_ (.I(_1351_),
    .Z(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2278_ (.I(_1341_),
    .Z(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2279_ (.I(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2280_ (.A1(_1334_),
    .A2(_1352_),
    .B(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2281_ (.A1(_1345_),
    .A2(_1349_),
    .B1(_1350_),
    .B2(_1355_),
    .ZN(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2282_ (.A1(_1278_),
    .A2(_1330_),
    .A3(_1338_),
    .B1(_1344_),
    .B2(_1356_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2283_ (.I(_1311_),
    .Z(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2284_ (.I(_1296_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2285_ (.I(_1258_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2286_ (.A1(_1340_),
    .A2(_1361_),
    .ZN(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2287_ (.A1(_1266_),
    .A2(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2288_ (.A1(_1290_),
    .A2(_1327_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2289_ (.A1(_1340_),
    .A2(_1265_),
    .Z(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2290_ (.A1(_1318_),
    .A2(_1365_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2291_ (.A1(_1360_),
    .A2(_1363_),
    .B1(_1364_),
    .B2(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2292_ (.A1(net47),
    .A2(_1339_),
    .ZN(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2293_ (.A1(_1340_),
    .A2(_1300_),
    .B(_1368_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2294_ (.A1(_1296_),
    .A2(_1362_),
    .A3(_1370_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2295_ (.A1(_1298_),
    .A2(_1323_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2296_ (.A1(_1264_),
    .A2(_1372_),
    .B(_1321_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _2297_ (.A1(_1281_),
    .A2(_1339_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2298_ (.A1(_1341_),
    .A2(_1302_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2299_ (.A1(_1362_),
    .A2(_1375_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2300_ (.I(_1281_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2301_ (.A1(_1371_),
    .A2(_1373_),
    .A3(_1374_),
    .B1(_1376_),
    .B2(_1377_),
    .ZN(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2302_ (.A1(_1367_),
    .A2(_1369_),
    .B(_1378_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2303_ (.I(_1380_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2304_ (.A1(_1359_),
    .A2(_1381_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2305_ (.A1(_1358_),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2306_ (.A1(_1315_),
    .A2(_1383_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2307_ (.A1(_1310_),
    .A2(_1384_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2308_ (.I(_1385_),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2309_ (.I(_1312_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2310_ (.I(_1386_),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2311_ (.A1(_1313_),
    .A2(_1342_),
    .B(_1281_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2312_ (.I(_1324_),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2313_ (.I(_1289_),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2314_ (.A1(_1390_),
    .A2(_1391_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2315_ (.A1(_1253_),
    .A2(_1348_),
    .B(_1347_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2316_ (.I(_1297_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2317_ (.I(_1351_),
    .Z(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2318_ (.A1(_1345_),
    .A2(_1394_),
    .A3(_1395_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2319_ (.A1(_1392_),
    .A2(_1393_),
    .B(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2320_ (.I(_1263_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2321_ (.I(_1398_),
    .Z(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2322_ (.I(_1399_),
    .Z(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2323_ (.A1(_1334_),
    .A2(_1401_),
    .B(_1348_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2324_ (.A1(_1324_),
    .A2(_1263_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2325_ (.I(_1403_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2326_ (.A1(_1352_),
    .A2(_1404_),
    .B(_1286_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2327_ (.I(_1372_),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2328_ (.A1(_1354_),
    .A2(_1406_),
    .A3(_1328_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2329_ (.I(_1261_),
    .Z(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2330_ (.A1(_1402_),
    .A2(_1405_),
    .B(_1407_),
    .C(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2331_ (.I(_1291_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2332_ (.I(_1410_),
    .Z(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2333_ (.A1(_1412_),
    .A2(_1338_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _2334_ (.A1(_1388_),
    .A2(_1397_),
    .B1(_1409_),
    .B2(_1413_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _2335_ (.A1(_1310_),
    .A2(_1387_),
    .A3(_1383_),
    .B1(_1414_),
    .B2(_1382_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2336_ (.I(_1311_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2337_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2338_ (.I(\p_shaping_I.counter[0] ),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2339_ (.I(_1311_),
    .Z(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2340_ (.I(_1369_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2341_ (.I(_1420_),
    .Z(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2342_ (.I(_1421_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2343_ (.I(\p_shaping_I.bit_in_2 ),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2344_ (.A1(_1367_),
    .A2(_1422_),
    .B(_1378_),
    .C(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2345_ (.A1(_1296_),
    .A2(_1379_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2346_ (.A1(_1299_),
    .A2(_1425_),
    .ZN(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2347_ (.A1(_1252_),
    .A2(_1264_),
    .B(_1318_),
    .C(_1266_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2348_ (.A1(_1399_),
    .A2(_1426_),
    .B(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2349_ (.A1(_1361_),
    .A2(_1255_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2350_ (.A1(_1299_),
    .A2(_1391_),
    .B(_1429_),
    .C(_1353_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2351_ (.A1(_1391_),
    .A2(_1327_),
    .B(_1321_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2352_ (.I(_1302_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2353_ (.A1(_1430_),
    .A2(_1431_),
    .B(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2354_ (.A1(_1272_),
    .A2(_1328_),
    .B(_1377_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2355_ (.A1(_1344_),
    .A2(_1428_),
    .B1(_1434_),
    .B2(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2356_ (.I(_1436_),
    .Z(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2357_ (.A1(_1424_),
    .A2(_1437_),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2358_ (.A1(_1419_),
    .A2(_1438_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2359_ (.I(_1398_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2360_ (.A1(_1390_),
    .A2(_1440_),
    .B(_1290_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2361_ (.I(_1441_),
    .Z(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2362_ (.I(_1322_),
    .Z(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2363_ (.A1(_1363_),
    .A2(_1442_),
    .B(_0026_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2364_ (.I(_1433_),
    .Z(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2365_ (.A1(_0028_),
    .A2(_1333_),
    .A3(_1271_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2366_ (.I(_1304_),
    .Z(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2367_ (.A1(_1332_),
    .A2(_0030_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2368_ (.A1(_0031_),
    .A2(_1393_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2369_ (.I(_1329_),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2370_ (.I(_1410_),
    .Z(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2371_ (.A1(_0027_),
    .A2(_0029_),
    .B1(_0032_),
    .B2(_0033_),
    .C(_0034_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2372_ (.I(_1284_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2373_ (.I(_0037_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2374_ (.A1(_1298_),
    .A2(_1361_),
    .B(_1323_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2375_ (.I(_0039_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2376_ (.A1(_1351_),
    .A2(_1327_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2377_ (.I(_0041_),
    .Z(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2378_ (.I(_1339_),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2379_ (.A1(_1253_),
    .A2(_1267_),
    .B(_0043_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2380_ (.A1(_0038_),
    .A2(_0040_),
    .B(_0042_),
    .C(_0044_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2381_ (.A1(_1412_),
    .A2(_1283_),
    .A3(_0045_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2382_ (.A1(_0035_),
    .A2(_0046_),
    .B(_0586_),
    .C(_1358_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2383_ (.I(_0570_),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2384_ (.A1(_1333_),
    .A2(_1271_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2385_ (.A1(_1335_),
    .A2(_1290_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _2386_ (.I(_0051_),
    .Z(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2387_ (.I(_1252_),
    .Z(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2388_ (.I(_1269_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2389_ (.A1(_0053_),
    .A2(_1287_),
    .B(_0054_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2390_ (.A1(_0052_),
    .A2(_0055_),
    .B(_1354_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2391_ (.A1(_0034_),
    .A2(_1305_),
    .A3(_1355_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2392_ (.A1(_0033_),
    .A2(_0050_),
    .A3(_0056_),
    .B1(_0057_),
    .B2(_1421_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2393_ (.A1(_1412_),
    .A2(_1283_),
    .A3(_0045_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2394_ (.A1(_0049_),
    .A2(_1414_),
    .B(_0059_),
    .C(_0060_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2395_ (.A1(_0048_),
    .A2(_0061_),
    .Z(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2396_ (.A1(_1359_),
    .A2(_1438_),
    .B1(_0048_),
    .B2(_0061_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2397_ (.A1(_1417_),
    .A2(_1418_),
    .B1(_1439_),
    .B2(_0062_),
    .C(_0063_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2398_ (.I(_1294_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2399_ (.I(_1370_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2400_ (.A1(_1317_),
    .A2(_0065_),
    .B(_0066_),
    .C(_1319_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2401_ (.A1(_0043_),
    .A2(_1257_),
    .A3(_0067_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2402_ (.A1(_1250_),
    .A2(_1440_),
    .B(_1331_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2403_ (.A1(_1305_),
    .A2(_0070_),
    .B(_1369_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2404_ (.A1(_1291_),
    .A2(_1260_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2405_ (.I(_0072_),
    .Z(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2406_ (.A1(_1300_),
    .A2(_1265_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2407_ (.A1(_1390_),
    .A2(_0074_),
    .B(_1321_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2408_ (.A1(_1366_),
    .A2(_0073_),
    .A3(_0075_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2409_ (.A1(_1282_),
    .A2(_0068_),
    .B(_0071_),
    .C(_0076_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2410_ (.I(_0601_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2411_ (.A1(_0078_),
    .A2(_1310_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2412_ (.A1(_0077_),
    .A2(_0079_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2413_ (.A1(_0064_),
    .A2(_0081_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2414_ (.A1(_1415_),
    .A2(_0082_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2415_ (.A1(_1439_),
    .A2(_0062_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2416_ (.A1(_1387_),
    .A2(_0063_),
    .A3(_0081_),
    .B(_0084_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2417_ (.I(\p_shaping_I.bit_in_2 ),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2418_ (.I(_0086_),
    .Z(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2419_ (.A1(_1381_),
    .A2(_1437_),
    .B(_0087_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2420_ (.A1(_1354_),
    .A2(_1267_),
    .B1(_0070_),
    .B2(_1292_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2421_ (.A1(_1301_),
    .A2(_1325_),
    .B(_0066_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2422_ (.A1(_1391_),
    .A2(_1404_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _2423_ (.A1(_1427_),
    .A2(_0090_),
    .B1(_0092_),
    .B2(_1319_),
    .C(_0072_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2424_ (.I(_1429_),
    .Z(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2425_ (.A1(_1269_),
    .A2(_1255_),
    .B(_1341_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2426_ (.A1(_1277_),
    .A2(_1313_),
    .A3(_0095_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2427_ (.A1(_1268_),
    .A2(_0054_),
    .A3(_1360_),
    .A4(_1254_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2428_ (.A1(_0094_),
    .A2(_0052_),
    .A3(_0096_),
    .A4(_0097_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2429_ (.A1(_1307_),
    .A2(_0089_),
    .B(_0093_),
    .C(_0098_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2430_ (.I(_0099_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2431_ (.A1(_0088_),
    .A2(_0100_),
    .Z(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2432_ (.A1(_0088_),
    .A2(_0100_),
    .B(_1416_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _2433_ (.A1(_1377_),
    .A2(_0043_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2434_ (.I(_1431_),
    .Z(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2435_ (.A1(_1250_),
    .A2(_0074_),
    .B(_1360_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2436_ (.A1(_0105_),
    .A2(_0106_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2437_ (.I(_1353_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2438_ (.A1(_1361_),
    .A2(_1255_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2439_ (.A1(_1390_),
    .A2(_0109_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2440_ (.I(_0110_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2441_ (.A1(_0108_),
    .A2(_0055_),
    .A3(_0111_),
    .B(_0106_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2442_ (.A1(_1268_),
    .A2(_0054_),
    .A3(_1331_),
    .A4(_1292_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2443_ (.A1(_1280_),
    .A2(_1285_),
    .A3(_1325_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2444_ (.A1(_1374_),
    .A2(_0114_),
    .A3(_0115_),
    .B(_1400_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2445_ (.A1(_0104_),
    .A2(_0107_),
    .B1(_0112_),
    .B2(_1420_),
    .C(_0116_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2446_ (.I(_0117_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2447_ (.A1(\p_shaping_I.bit_in ),
    .A2(_0605_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2448_ (.A1(_0592_),
    .A2(_0119_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2449_ (.A1(_0118_),
    .A2(_0120_),
    .ZN(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2450_ (.A1(_1358_),
    .A2(_0035_),
    .A3(_0046_),
    .B(_0578_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2451_ (.A1(_0121_),
    .A2(_0122_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2452_ (.A1(_0101_),
    .A2(_0103_),
    .A3(_0123_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2453_ (.A1(_0101_),
    .A2(_0103_),
    .B(_0123_),
    .ZN(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2454_ (.A1(_1279_),
    .A2(_1309_),
    .B(_0077_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2455_ (.A1(_0603_),
    .A2(_0127_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2456_ (.A1(_1440_),
    .A2(_1325_),
    .B(_1318_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2457_ (.A1(_1401_),
    .A2(_1393_),
    .B(_0129_),
    .C(_0104_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2458_ (.A1(_1301_),
    .A2(_1351_),
    .B(_1353_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2459_ (.A1(_1392_),
    .A2(_0131_),
    .B(_0042_),
    .C(_0073_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2460_ (.A1(_1286_),
    .A2(_0092_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2461_ (.A1(_0111_),
    .A2(_0133_),
    .B(_0031_),
    .C(_1420_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _2462_ (.A1(_0130_),
    .A2(_0132_),
    .A3(_0134_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2463_ (.A1(_0128_),
    .A2(_0136_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2464_ (.A1(_1314_),
    .A2(_0125_),
    .A3(_0126_),
    .A4(_0137_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2465_ (.A1(_1387_),
    .A2(_0125_),
    .A3(_0126_),
    .B(_0137_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2466_ (.A1(_0085_),
    .A2(_0138_),
    .A3(_0139_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2467_ (.A1(_0138_),
    .A2(_0139_),
    .B(_0085_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2468_ (.A1(_0140_),
    .A2(_0141_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2469_ (.A1(_0083_),
    .A2(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2470_ (.I(_0143_),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2471_ (.I(_1314_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2472_ (.A1(_0101_),
    .A2(_0103_),
    .A3(_0123_),
    .ZN(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2473_ (.A1(_0144_),
    .A2(_0126_),
    .A3(_0137_),
    .B(_0146_),
    .ZN(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2474_ (.I(\p_shaping_I.counter[1] ),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2475_ (.A1(_1440_),
    .A2(_1303_),
    .B1(_1403_),
    .B2(_0039_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2476_ (.A1(_0075_),
    .A2(_0149_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2477_ (.A1(_1308_),
    .A2(_0150_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2478_ (.A1(_1274_),
    .A2(_0090_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2479_ (.A1(_1399_),
    .A2(_1254_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2480_ (.A1(_0037_),
    .A2(_1406_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2481_ (.A1(_0153_),
    .A2(_0154_),
    .B(_1369_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2482_ (.A1(_0152_),
    .A2(_0155_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2483_ (.A1(_1322_),
    .A2(_1442_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2484_ (.A1(_0053_),
    .A2(_1301_),
    .B(_1303_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2485_ (.I(_1362_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2486_ (.A1(_0052_),
    .A2(_0159_),
    .B(_0160_),
    .C(_0108_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2487_ (.A1(_0052_),
    .A2(_0158_),
    .B(_0161_),
    .C(_1374_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _2488_ (.A1(_0151_),
    .A2(_0157_),
    .A3(_0162_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2489_ (.A1(_1381_),
    .A2(_1437_),
    .A3(_0099_),
    .B(_0086_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2490_ (.A1(_0163_),
    .A2(_0164_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2491_ (.I(_0118_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2492_ (.A1(_1414_),
    .A2(_0059_),
    .A3(_0060_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2493_ (.A1(_1400_),
    .A2(_0119_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2494_ (.A1(_1297_),
    .A2(_1392_),
    .ZN(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2495_ (.A1(_0039_),
    .A2(_0041_),
    .B(_0037_),
    .ZN(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2496_ (.A1(_0170_),
    .A2(_0171_),
    .B(_1388_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2497_ (.I(_0172_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2498_ (.A1(_1364_),
    .A2(_1366_),
    .ZN(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2499_ (.A1(_0051_),
    .A2(_0159_),
    .B(_1360_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2500_ (.A1(_1260_),
    .A2(_0095_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2501_ (.A1(_0129_),
    .A2(_0176_),
    .B(_1277_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2502_ (.A1(_1433_),
    .A2(_0174_),
    .A3(_0175_),
    .B(_0177_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2503_ (.I(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2504_ (.A1(_0169_),
    .A2(_0173_),
    .A3(_0180_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2505_ (.I(_0578_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2506_ (.A1(_0166_),
    .A2(_0168_),
    .B(_0181_),
    .C(_0182_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2507_ (.I(_0570_),
    .Z(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2508_ (.A1(_0169_),
    .A2(_0173_),
    .A3(_0180_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2509_ (.A1(_0184_),
    .A2(_0118_),
    .B(_0122_),
    .C(_0185_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2510_ (.A1(_0148_),
    .A2(_0165_),
    .B1(_0183_),
    .B2(_0186_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2511_ (.A1(_0148_),
    .A2(_0165_),
    .A3(_0183_),
    .A4(_0186_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2512_ (.A1(_1332_),
    .A2(_1352_),
    .B(_0160_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2513_ (.A1(_1336_),
    .A2(_0131_),
    .B(_1262_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2514_ (.A1(_0043_),
    .A2(_0129_),
    .B1(_1441_),
    .B2(_1375_),
    .C(_1377_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2515_ (.A1(_0190_),
    .A2(_0191_),
    .B(_0192_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2516_ (.A1(_1322_),
    .A2(_0074_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2517_ (.A1(_1317_),
    .A2(_0065_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2518_ (.A1(_0194_),
    .A2(_0065_),
    .B1(_0195_),
    .B2(_0038_),
    .C(_1307_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _2519_ (.A1(_1411_),
    .A2(_0193_),
    .A3(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2520_ (.A1(_0127_),
    .A2(_0136_),
    .B(_0602_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2521_ (.A1(_0197_),
    .A2(_0198_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2522_ (.A1(_1312_),
    .A2(_0187_),
    .A3(_0188_),
    .A4(_0199_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2523_ (.A1(_0144_),
    .A2(_0187_),
    .A3(_0188_),
    .B(_0199_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2524_ (.A1(_0201_),
    .A2(_0202_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2525_ (.A1(_0083_),
    .A2(_0142_),
    .B(_0140_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2526_ (.A1(_0147_),
    .A2(_0203_),
    .A3(_0204_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2527_ (.I(_0205_),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2528_ (.I(_0148_),
    .Z(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2529_ (.A1(_0206_),
    .A2(_0165_),
    .A3(_0183_),
    .A4(_0186_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2530_ (.A1(_0207_),
    .A2(_0201_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2531_ (.A1(_1381_),
    .A2(_1437_),
    .A3(_0099_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2532_ (.A1(_0163_),
    .A2(_0209_),
    .B(_1423_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2533_ (.A1(_1347_),
    .A2(_1404_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2534_ (.I(_1337_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2535_ (.A1(_0212_),
    .A2(_0213_),
    .B(_1420_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2536_ (.A1(_1410_),
    .A2(_1407_),
    .A3(_0105_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2537_ (.A1(_0108_),
    .A2(_0055_),
    .A3(_0111_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2538_ (.A1(_1299_),
    .A2(_1303_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2539_ (.A1(_1270_),
    .A2(_1406_),
    .B(_0217_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2540_ (.A1(_1347_),
    .A2(_0218_),
    .B(_1282_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2541_ (.A1(_0216_),
    .A2(_0219_),
    .B(_0028_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2542_ (.A1(_0214_),
    .A2(_0215_),
    .A3(_0220_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2543_ (.A1(_0211_),
    .A2(_0222_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2544_ (.I(_0169_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2545_ (.A1(_0053_),
    .A2(_1280_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2546_ (.A1(_1319_),
    .A2(_0225_),
    .A3(_0110_),
    .B(_0131_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2547_ (.A1(_1399_),
    .A2(_1297_),
    .A3(_1406_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2548_ (.A1(_0037_),
    .A2(_0066_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2549_ (.A1(_0227_),
    .A2(_0228_),
    .B(_1261_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2550_ (.A1(_1285_),
    .A2(_0066_),
    .Z(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2551_ (.A1(_1433_),
    .A2(_0115_),
    .A3(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2552_ (.A1(_0226_),
    .A2(_0229_),
    .B(_0231_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2553_ (.A1(_0194_),
    .A2(_0056_),
    .B(_1408_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2554_ (.I0(_0233_),
    .I1(_0234_),
    .S(_1278_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2555_ (.A1(_0117_),
    .A2(_0172_),
    .A3(_0179_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2556_ (.A1(_0235_),
    .A2(_0236_),
    .B(_0570_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2557_ (.I(_0237_),
    .Z(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2558_ (.A1(_0224_),
    .A2(_0238_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2559_ (.I(_1278_),
    .Z(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2560_ (.I(_1365_),
    .Z(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2561_ (.A1(_0241_),
    .A2(_0040_),
    .B(_1329_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2562_ (.A1(_1274_),
    .A2(_0225_),
    .A3(_0111_),
    .B(_0242_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2563_ (.A1(_1343_),
    .A2(_0244_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2564_ (.A1(_0026_),
    .A2(_1271_),
    .Z(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2565_ (.A1(_1345_),
    .A2(_1401_),
    .B(_0073_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2566_ (.I(_0053_),
    .Z(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2567_ (.A1(_0248_),
    .A2(_0026_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2568_ (.A1(_0249_),
    .A2(_1350_),
    .A3(_1396_),
    .A4(_1421_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2569_ (.A1(_0246_),
    .A2(_0247_),
    .B(_0250_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2570_ (.A1(_0240_),
    .A2(_0245_),
    .B(_0251_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2571_ (.A1(_0049_),
    .A2(_0236_),
    .B(_0252_),
    .C(_0122_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2572_ (.A1(_0117_),
    .A2(_0173_),
    .A3(_0180_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2573_ (.A1(_1388_),
    .A2(_0244_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2574_ (.A1(_0256_),
    .A2(_0251_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2575_ (.A1(_0168_),
    .A2(_0255_),
    .B(_0257_),
    .C(_0182_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2576_ (.A1(_0224_),
    .A2(_0253_),
    .A3(_0258_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2577_ (.A1(_1359_),
    .A2(_0223_),
    .B(_0239_),
    .C(_0259_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2578_ (.A1(_0184_),
    .A2(_0118_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2579_ (.A1(_0226_),
    .A2(_0229_),
    .B(_0231_),
    .C(_1410_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2580_ (.A1(_0034_),
    .A2(_0234_),
    .B(_0262_),
    .C(\p_shaping_I.bit_in_1 ),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2581_ (.A1(_0173_),
    .A2(_0180_),
    .B(_0184_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2582_ (.A1(_0169_),
    .A2(_0261_),
    .A3(_0263_),
    .A4(_0264_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2583_ (.I(_0224_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2584_ (.A1(_0267_),
    .A2(_0253_),
    .A3(_0258_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2585_ (.A1(_0211_),
    .A2(_0222_),
    .B(_1419_),
    .ZN(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2586_ (.A1(_0211_),
    .A2(_0222_),
    .B1(_0266_),
    .B2(_0268_),
    .C(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2587_ (.A1(_1314_),
    .A2(_0260_),
    .A3(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2588_ (.I(_0108_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2589_ (.A1(_1365_),
    .A2(_0094_),
    .A3(_0039_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2590_ (.A1(_0272_),
    .A2(_0273_),
    .B(_1308_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2591_ (.A1(_0272_),
    .A2(_1404_),
    .A3(_0074_),
    .B(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2592_ (.A1(_0248_),
    .A2(_0213_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2593_ (.I(_1372_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2594_ (.A1(_1332_),
    .A2(_0278_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2595_ (.A1(_1363_),
    .A2(_0279_),
    .B(_0176_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2596_ (.I(_1282_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2597_ (.A1(_0033_),
    .A2(_0277_),
    .B(_0280_),
    .C(_0281_),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2598_ (.A1(_0275_),
    .A2(_0282_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2599_ (.A1(_0127_),
    .A2(_0136_),
    .A3(_0197_),
    .B(_0602_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2600_ (.A1(_0283_),
    .A2(_0284_),
    .Z(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _2601_ (.A1(_0208_),
    .A2(_0271_),
    .A3(_0285_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2602_ (.A1(_0146_),
    .A2(_0138_),
    .A3(_0203_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2603_ (.A1(_1415_),
    .A2(_0082_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2604_ (.A1(_0147_),
    .A2(_0201_),
    .A3(_0202_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2605_ (.A1(_0085_),
    .A2(_0138_),
    .A3(_0139_),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _2606_ (.A1(_0289_),
    .A2(_0141_),
    .B(_0290_),
    .C(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2607_ (.A1(_0288_),
    .A2(_0292_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2608_ (.A1(_0286_),
    .A2(_0293_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2609_ (.I(_0294_),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2610_ (.A1(_0239_),
    .A2(_0259_),
    .B(_0206_),
    .C(_0223_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2611_ (.A1(_1386_),
    .A2(_0260_),
    .A3(_0285_),
    .B(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2612_ (.I(_1317_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2613_ (.I(_1286_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _2614_ (.A1(_1401_),
    .A2(_0298_),
    .B(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2615_ (.A1(_1402_),
    .A2(_1405_),
    .B(_1421_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2616_ (.I(_0028_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2617_ (.A1(_0038_),
    .A2(_0030_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2618_ (.A1(_1394_),
    .A2(_1365_),
    .A3(_0094_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2619_ (.A1(_0303_),
    .A2(_0304_),
    .ZN(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2620_ (.A1(_0302_),
    .A2(_0305_),
    .B(_1412_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2621_ (.A1(_0241_),
    .A2(_1336_),
    .A3(_0213_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _2622_ (.A1(_0302_),
    .A2(_1407_),
    .A3(_0307_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _2623_ (.A1(_0300_),
    .A2(_0301_),
    .B(_0306_),
    .C(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2624_ (.A1(_0151_),
    .A2(_0157_),
    .A3(_0162_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2625_ (.A1(_1380_),
    .A2(_1436_),
    .A3(_0099_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2626_ (.A1(_0311_),
    .A2(_0312_),
    .A3(_0222_),
    .B(_0087_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2627_ (.A1(_0310_),
    .A2(_0313_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2628_ (.A1(_0049_),
    .A2(_0236_),
    .B(_0235_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2629_ (.A1(_0120_),
    .A2(_0263_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2630_ (.A1(_1359_),
    .A2(_0314_),
    .B1(_0315_),
    .B2(_0316_),
    .C(_0239_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2631_ (.A1(_0310_),
    .A2(_0313_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2632_ (.I(_0120_),
    .Z(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2633_ (.A1(_0578_),
    .A2(_0255_),
    .B(_0263_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2634_ (.A1(_0320_),
    .A2(_0321_),
    .B1(_0315_),
    .B2(_0316_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2635_ (.I(_1312_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2636_ (.A1(_1416_),
    .A2(_0318_),
    .A3(_0322_),
    .B(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2637_ (.A1(_0317_),
    .A2(_0324_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2638_ (.A1(_0272_),
    .A2(_0298_),
    .B1(_0095_),
    .B2(_0042_),
    .C(_0302_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2639_ (.A1(_0240_),
    .A2(_1342_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2640_ (.A1(_0038_),
    .A2(_0298_),
    .B(_1408_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2641_ (.A1(_1273_),
    .A2(_0050_),
    .B(_0154_),
    .C(_0328_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2642_ (.A1(_0281_),
    .A2(_0329_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2643_ (.A1(_0326_),
    .A2(_0327_),
    .B(_0331_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _2644_ (.A1(_0127_),
    .A2(_0136_),
    .A3(_0197_),
    .A4(_0283_),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2645_ (.A1(_0601_),
    .A2(_0333_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2646_ (.A1(_0332_),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2647_ (.A1(_0296_),
    .A2(_0325_),
    .A3(_0335_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _2648_ (.A1(_1387_),
    .A2(_0260_),
    .A3(_0270_),
    .A4(_0285_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2649_ (.A1(_0144_),
    .A2(_0260_),
    .A3(_0270_),
    .B(_0285_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2650_ (.A1(_0208_),
    .A2(_0337_),
    .A3(_0338_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2651_ (.A1(_0286_),
    .A2(_0293_),
    .B(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2652_ (.A1(_0336_),
    .A2(_0340_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2653_ (.I(_0342_),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2654_ (.A1(_1417_),
    .A2(_0318_),
    .A3(_0322_),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2655_ (.A1(_0325_),
    .A2(_0335_),
    .B(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2656_ (.I(_1423_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2657_ (.A1(_0214_),
    .A2(_0215_),
    .A3(_0220_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2658_ (.A1(_0163_),
    .A2(_0209_),
    .A3(_0346_),
    .A4(_0310_),
    .Z(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2659_ (.I(_0104_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2660_ (.A1(_0299_),
    .A2(_0348_),
    .A3(_0030_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2661_ (.A1(_1395_),
    .A2(_0160_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2662_ (.A1(_0033_),
    .A2(_0350_),
    .A3(_0040_),
    .Z(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2663_ (.I(_1408_),
    .Z(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2664_ (.A1(_0353_),
    .A2(_1426_),
    .B1(_0092_),
    .B2(_0095_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2665_ (.A1(_1333_),
    .A2(_0133_),
    .B(_0352_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2666_ (.I(_0281_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2667_ (.A1(_0352_),
    .A2(_0354_),
    .B(_0355_),
    .C(_0356_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2668_ (.A1(_0349_),
    .A2(_0357_),
    .Z(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2669_ (.A1(_0345_),
    .A2(_0347_),
    .B(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2670_ (.I(_0087_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2671_ (.A1(_0349_),
    .A2(_0357_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2672_ (.A1(_0163_),
    .A2(_0209_),
    .A3(_0346_),
    .A4(_0310_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2673_ (.A1(_0360_),
    .A2(_0361_),
    .A3(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2674_ (.I(_0054_),
    .Z(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2675_ (.A1(_0365_),
    .A2(_1394_),
    .A3(_1352_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2676_ (.A1(_0248_),
    .A2(_1329_),
    .A3(_0109_),
    .A4(_0094_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2677_ (.A1(_0366_),
    .A2(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2678_ (.A1(_0028_),
    .A2(_0195_),
    .A3(_0131_),
    .B1(_0367_),
    .B2(_0366_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2679_ (.A1(_0368_),
    .A2(_0369_),
    .B(_0281_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2680_ (.A1(_0365_),
    .A2(_0278_),
    .B1(_1295_),
    .B2(_1305_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2681_ (.A1(_0365_),
    .A2(_1394_),
    .A3(_0278_),
    .A4(_1295_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2682_ (.A1(_1308_),
    .A2(_0371_),
    .A3(_0372_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2683_ (.A1(_0370_),
    .A2(_0374_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2684_ (.A1(_0182_),
    .A2(_0255_),
    .B(_0375_),
    .C(_0263_),
    .ZN(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2685_ (.A1(_0370_),
    .A2(_0374_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2686_ (.A1(_0235_),
    .A2(_0236_),
    .B(_0377_),
    .C(_0184_),
    .ZN(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2687_ (.A1(_0320_),
    .A2(_0376_),
    .A3(_0378_),
    .B(_0266_),
    .ZN(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2688_ (.A1(_1419_),
    .A2(_0359_),
    .A3(_0364_),
    .A4(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2689_ (.A1(_0360_),
    .A2(_0363_),
    .B(_0361_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2690_ (.A1(_1423_),
    .A2(_0358_),
    .A3(_0347_),
    .B(_0148_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2691_ (.A1(_0320_),
    .A2(_0376_),
    .A3(_0378_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2692_ (.A1(_0381_),
    .A2(_0382_),
    .B(_0383_),
    .C(_0266_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2693_ (.A1(_0323_),
    .A2(_0380_),
    .A3(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2694_ (.A1(_0332_),
    .A2(_0333_),
    .B(_0601_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2695_ (.I(_0353_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2696_ (.I(_0272_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2697_ (.A1(_0298_),
    .A2(_1328_),
    .B(_0217_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2698_ (.A1(_0389_),
    .A2(_0390_),
    .B(_0213_),
    .C(_0353_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2699_ (.A1(_0388_),
    .A2(_1425_),
    .B(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2700_ (.I(_0356_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2701_ (.A1(_0348_),
    .A2(_0226_),
    .B1(_0392_),
    .B2(_0393_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2702_ (.A1(_0387_),
    .A2(_0394_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2703_ (.A1(_0386_),
    .A2(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2704_ (.A1(_0344_),
    .A2(_0397_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _2705_ (.A1(_0288_),
    .A2(_0286_),
    .A3(_0292_),
    .A4(_0336_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2706_ (.A1(_0317_),
    .A2(_0324_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2707_ (.I(_0335_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2708_ (.A1(_0400_),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2709_ (.A1(_0400_),
    .A2(_0401_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2710_ (.A1(_0317_),
    .A2(_0324_),
    .A3(_0401_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2711_ (.A1(_0317_),
    .A2(_0324_),
    .B(_0401_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2712_ (.A1(_0295_),
    .A2(_0337_),
    .B1(_0404_),
    .B2(_0405_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2713_ (.A1(_0296_),
    .A2(_0402_),
    .A3(_0403_),
    .B1(_0407_),
    .B2(_0339_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2714_ (.A1(_0399_),
    .A2(_0408_),
    .Z(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2715_ (.A1(_0398_),
    .A2(_0409_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2716_ (.I(_0410_),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2717_ (.A1(_0386_),
    .A2(_0396_),
    .B(_0380_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2718_ (.I(_0073_),
    .Z(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _2719_ (.A1(_0299_),
    .A2(_1442_),
    .B1(_0195_),
    .B2(_0105_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _2720_ (.A1(_1364_),
    .A2(_1366_),
    .B(_0249_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2721_ (.A1(_1348_),
    .A2(_1336_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2722_ (.A1(_0026_),
    .A2(_0415_),
    .A3(_1364_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2723_ (.I(_0365_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2724_ (.A1(_0418_),
    .A2(_0034_),
    .A3(_1389_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2725_ (.A1(_0155_),
    .A2(_0417_),
    .B(_0419_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2726_ (.A1(_0412_),
    .A2(_0413_),
    .B1(_0414_),
    .B2(_0104_),
    .C(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2727_ (.A1(_0182_),
    .A2(_0421_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2728_ (.A1(_0237_),
    .A2(_0421_),
    .B(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2729_ (.A1(_0267_),
    .A2(_0423_),
    .Z(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2730_ (.A1(_0087_),
    .A2(_0363_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2731_ (.I(_0302_),
    .Z(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2732_ (.A1(_1350_),
    .A2(_0092_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2733_ (.A1(_1273_),
    .A2(_0415_),
    .B(_0356_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2734_ (.A1(_0426_),
    .A2(_0428_),
    .B(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2735_ (.A1(_0216_),
    .A2(_0328_),
    .B(_0430_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2736_ (.A1(_0345_),
    .A2(_0347_),
    .A3(_0431_),
    .B(_1419_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2737_ (.A1(_0425_),
    .A2(_0431_),
    .B(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2738_ (.A1(_0424_),
    .A2(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _2739_ (.I(_0299_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2740_ (.A1(_0435_),
    .A2(_0090_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2741_ (.A1(_0435_),
    .A2(_1350_),
    .B(_0436_),
    .C(_0348_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2742_ (.I(_0389_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _2743_ (.A1(_0439_),
    .A2(_0241_),
    .A3(_0040_),
    .A4(_0412_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2744_ (.A1(_0592_),
    .A2(_0437_),
    .A3(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2745_ (.A1(_0387_),
    .A2(_0441_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2746_ (.A1(_0144_),
    .A2(_0434_),
    .A3(_0442_),
    .Z(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2747_ (.A1(_1315_),
    .A2(_0434_),
    .B(_0442_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2748_ (.A1(_0411_),
    .A2(_0443_),
    .A3(_0444_),
    .Z(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2749_ (.A1(_0443_),
    .A2(_0444_),
    .B(_0411_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2750_ (.A1(_0445_),
    .A2(_0446_),
    .ZN(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _2751_ (.A1(_0344_),
    .A2(_0397_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2752_ (.A1(_0398_),
    .A2(_0409_),
    .B(_0448_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2753_ (.A1(_0447_),
    .A2(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2754_ (.I(_0451_),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2755_ (.A1(_0424_),
    .A2(_0433_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2756_ (.A1(_0452_),
    .A2(_0443_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2757_ (.A1(_0105_),
    .A2(_0195_),
    .B(_1388_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2758_ (.A1(_0389_),
    .A2(_0153_),
    .A3(_0160_),
    .B(_0279_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _2759_ (.A1(_1375_),
    .A2(_0390_),
    .B1(_0455_),
    .B2(_0388_),
    .C(_0356_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2760_ (.A1(_1274_),
    .A2(_1442_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2761_ (.A1(_0454_),
    .A2(_0456_),
    .B1(_0457_),
    .B2(_0388_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2762_ (.A1(_0586_),
    .A2(_0458_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2763_ (.A1(_0238_),
    .A2(_0458_),
    .B(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2764_ (.A1(_0238_),
    .A2(_0421_),
    .B(_0422_),
    .C(_0224_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2765_ (.A1(_0267_),
    .A2(_0461_),
    .B(_0462_),
    .C(_1386_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2766_ (.A1(_1320_),
    .A2(_0042_),
    .B(_0328_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2767_ (.A1(_0426_),
    .A2(_0230_),
    .B(_0429_),
    .C(_0464_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2768_ (.A1(_0360_),
    .A2(_0245_),
    .B(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2769_ (.A1(_0425_),
    .A2(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2770_ (.A1(_0360_),
    .A2(_0465_),
    .B(_1417_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2771_ (.A1(_0467_),
    .A2(_0468_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2772_ (.A1(_0463_),
    .A2(_0469_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2773_ (.A1(_1425_),
    .A2(_0303_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2774_ (.A1(_0393_),
    .A2(_1283_),
    .ZN(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2775_ (.A1(_0435_),
    .A2(_0388_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2776_ (.I(_0240_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2777_ (.A1(_0241_),
    .A2(_0474_),
    .B(_0475_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _2778_ (.A1(_0348_),
    .A2(_0472_),
    .B(_0473_),
    .C(_0476_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2779_ (.A1(_0078_),
    .A2(_0477_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2780_ (.A1(_0332_),
    .A2(_0333_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _2781_ (.A1(_1345_),
    .A2(_0300_),
    .B1(_0273_),
    .B2(_0435_),
    .C(_0426_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2782_ (.A1(_0078_),
    .A2(_0477_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2783_ (.A1(_0479_),
    .A2(_0480_),
    .B(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2784_ (.A1(_0478_),
    .A2(_0483_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2785_ (.A1(_0471_),
    .A2(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2786_ (.A1(_0453_),
    .A2(_0485_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2787_ (.A1(_0399_),
    .A2(_0408_),
    .B(_0398_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2788_ (.A1(_0448_),
    .A2(_0446_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _2789_ (.A1(_0487_),
    .A2(_0447_),
    .B(_0488_),
    .C(_0445_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2790_ (.A1(_0486_),
    .A2(_0489_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2791_ (.I(_0490_),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2792_ (.A1(_0463_),
    .A2(_0467_),
    .A3(_0468_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _2793_ (.A1(_0471_),
    .A2(_0484_),
    .B(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2794_ (.A1(_1295_),
    .A2(_1326_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _2795_ (.A1(_1405_),
    .A2(_1422_),
    .A3(_0494_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _2796_ (.A1(_0412_),
    .A2(_0228_),
    .B1(_0480_),
    .B2(_0475_),
    .C(_0495_),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2797_ (.A1(_0238_),
    .A2(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2798_ (.A1(_0586_),
    .A2(_0496_),
    .B(_0267_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2799_ (.A1(_1386_),
    .A2(_0462_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2800_ (.A1(_0497_),
    .A2(_0498_),
    .B(_0499_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2801_ (.I(_0429_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2802_ (.I(_0426_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2803_ (.A1(_0472_),
    .A2(_0350_),
    .B(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2804_ (.A1(_0501_),
    .A2(_0504_),
    .B(_0425_),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _2805_ (.A1(_0345_),
    .A2(_0501_),
    .A3(_0504_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2806_ (.A1(_0206_),
    .A2(_0505_),
    .A3(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2807_ (.A1(_0500_),
    .A2(_0507_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2808_ (.A1(_0473_),
    .A2(_0476_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2809_ (.A1(_0393_),
    .A2(_0472_),
    .B(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2810_ (.A1(_0387_),
    .A2(_0510_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2811_ (.A1(_0603_),
    .A2(_0510_),
    .B(_0511_),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2812_ (.A1(_0508_),
    .A2(_0512_),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2813_ (.A1(_0493_),
    .A2(_0514_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2814_ (.A1(_0452_),
    .A2(_0443_),
    .B(_0485_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2815_ (.A1(_0486_),
    .A2(_0489_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2816_ (.A1(_0516_),
    .A2(_0517_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2817_ (.A1(_0515_),
    .A2(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2818_ (.I(_0519_),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2819_ (.I(_0323_),
    .Z(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2820_ (.A1(_0120_),
    .A2(_0321_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _2821_ (.A1(_0389_),
    .A2(_1251_),
    .B(_0353_),
    .C(_1395_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2822_ (.A1(_1422_),
    .A2(_0305_),
    .B1(_0521_),
    .B2(_0240_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2823_ (.A1(_0520_),
    .A2(_0523_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2824_ (.A1(_0025_),
    .A2(_0524_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2825_ (.A1(_0503_),
    .A2(_1342_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2826_ (.A1(_0501_),
    .A2(_0526_),
    .B(_0425_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _2827_ (.A1(_0345_),
    .A2(_0501_),
    .A3(_0526_),
    .B(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _2828_ (.A1(_1417_),
    .A2(_0528_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2829_ (.A1(_0525_),
    .A2(_0529_),
    .Z(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2830_ (.A1(_0078_),
    .A2(_0476_),
    .B1(_0509_),
    .B2(_0387_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _2831_ (.I(_0531_),
    .Z(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2832_ (.A1(_0530_),
    .A2(_0532_),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2833_ (.A1(_0508_),
    .A2(_0512_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2834_ (.A1(_0500_),
    .A2(_0507_),
    .B(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _2835_ (.A1(_0534_),
    .A2(_0536_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2836_ (.I(_0537_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2837_ (.A1(_0493_),
    .A2(_0514_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2838_ (.A1(_0493_),
    .A2(_0514_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2839_ (.A1(_0516_),
    .A2(_0539_),
    .B(_0540_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _2840_ (.A1(_0486_),
    .A2(_0489_),
    .A3(_0515_),
    .B(_0541_),
    .ZN(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2841_ (.A1(_0538_),
    .A2(_0542_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2842_ (.I(_0543_),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2843_ (.A1(_0025_),
    .A2(_0524_),
    .A3(_0529_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2844_ (.A1(_0530_),
    .A2(_0532_),
    .B(_0545_),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _2845_ (.A1(_0475_),
    .A2(_1375_),
    .B1(_0304_),
    .B2(_1422_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2846_ (.A1(_0049_),
    .A2(_0547_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2847_ (.A1(_0321_),
    .A2(_0547_),
    .B(_0548_),
    .ZN(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2848_ (.A1(_0320_),
    .A2(_0549_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _2849_ (.A1(_1315_),
    .A2(_0462_),
    .A3(_0550_),
    .ZN(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _2850_ (.A1(_0529_),
    .A2(_0531_),
    .A3(_0551_),
    .Z(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2851_ (.A1(_0546_),
    .A2(_0552_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2852_ (.A1(_0534_),
    .A2(_0536_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2853_ (.A1(_0538_),
    .A2(_0542_),
    .B(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2854_ (.A1(_0553_),
    .A2(_0556_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2855_ (.I(_0557_),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2856_ (.A1(_0537_),
    .A2(_0553_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2857_ (.A1(_0542_),
    .A2(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2858_ (.I(_0552_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2859_ (.A1(_0546_),
    .A2(_0560_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2860_ (.A1(_0546_),
    .A2(_0560_),
    .B(_0555_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2861_ (.A1(_0561_),
    .A2(_0562_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2862_ (.A1(_0532_),
    .A2(_0551_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2863_ (.A1(_0532_),
    .A2(_0551_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2864_ (.A1(_0529_),
    .A2(_0564_),
    .B(_0565_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2865_ (.A1(_0559_),
    .A2(_0563_),
    .A3(_0566_),
    .B1(_0520_),
    .B2(_1315_),
    .ZN(net7));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2866_ (.A1(_1415_),
    .A2(_0082_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2867_ (.I(_0567_),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2868_ (.A1(\bit2symb.regi ),
    .A2(_1411_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2869_ (.A1(_0603_),
    .A2(net42),
    .B(_0568_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2870_ (.I0(net1),
    .I1(\Reg_Delay_Q.In ),
    .S(_0599_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2871_ (.I(_0569_),
    .Z(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _2872_ (.A1(_0439_),
    .A2(_0415_),
    .A3(_0412_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2873_ (.I(_0571_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2874_ (.A1(\Reg_Delay_Q.In ),
    .A2(_0572_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2875_ (.A1(_0612_),
    .A2(_0572_),
    .B(_0573_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2876_ (.I(net2),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2877_ (.A1(_0418_),
    .A2(_0574_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2878_ (.I(_0575_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2879_ (.I(_0574_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2880_ (.A1(_0574_),
    .A2(_0065_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2881_ (.A1(_0248_),
    .A2(_0576_),
    .B1(net42),
    .B2(_0577_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2882_ (.A1(_0418_),
    .A2(net2),
    .ZN(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _2883_ (.A1(_0278_),
    .A2(_0579_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2884_ (.I(_0580_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _2885_ (.A1(_1395_),
    .A2(_0579_),
    .B(_0581_),
    .C(_0217_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _2886_ (.A1(_0439_),
    .A2(_0581_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2887_ (.I(_0582_),
    .Z(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2888_ (.A1(_0439_),
    .A2(_0580_),
    .B(_0503_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _2889_ (.A1(_0574_),
    .A2(net42),
    .B1(_0581_),
    .B2(_0474_),
    .C(_0583_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2890_ (.I(net2),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _2891_ (.A1(_0418_),
    .A2(_0503_),
    .A3(_0584_),
    .A4(_1389_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _2892_ (.I(_0584_),
    .ZN(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _2893_ (.A1(_0393_),
    .A2(_0587_),
    .A3(_0030_),
    .A4(_1273_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2894_ (.A1(_0474_),
    .A2(_0581_),
    .B(_0475_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _2895_ (.A1(_0585_),
    .A2(_0588_),
    .A3(_0589_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2896_ (.A1(_0584_),
    .A2(_0571_),
    .ZN(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2897_ (.A1(_0857_),
    .A2(_0587_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _2898_ (.A1(_0857_),
    .A2(_0590_),
    .B(_0591_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2899_ (.A1(_0756_),
    .A2(_0576_),
    .B1(_0952_),
    .B2(_0590_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2900_ (.A1(_0834_),
    .A2(_0817_),
    .A3(_0590_),
    .B1(_0576_),
    .B2(_0943_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _2901_ (.A1(_1024_),
    .A2(_0788_),
    .A3(_0590_),
    .B1(_0576_),
    .B2(_1054_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _2902_ (.A1(_0584_),
    .A2(_0571_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2903_ (.A1(_0788_),
    .A2(_0593_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2904_ (.A1(_0870_),
    .A2(_0572_),
    .B(_0587_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _2905_ (.A1(_0762_),
    .A2(_0594_),
    .B(_0595_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _2906_ (.A1(_1158_),
    .A2(_0595_),
    .B1(_0594_),
    .B2(_0712_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2907_ (.A1(_0828_),
    .A2(\p_shaping_Q.counter[0] ),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2908_ (.A1(_0022_),
    .A2(_0596_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2909_ (.A1(_0592_),
    .A2(_0572_),
    .ZN(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _2910_ (.I0(\bit2symb.regi ),
    .I1(net1),
    .S(_0597_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _2911_ (.I(_0598_),
    .Z(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2912_ (.A1(_0206_),
    .A2(\p_shaping_I.counter[0] ),
    .ZN(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _2913_ (.A1(_0025_),
    .A2(_0600_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2914_ (.D(_0006_),
    .RN(net53),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(\p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2915_ (.D(_0007_),
    .RN(net52),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(\Reg_Delay_Q.In ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2916_ (.D(_0008_),
    .RN(net52),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(\Reg_Delay_Q.Out ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2917_ (.D(_0009_),
    .RN(net54),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2918_ (.D(_0010_),
    .RN(net53),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2919_ (.D(_0011_),
    .RN(net54),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2920_ (.D(_0012_),
    .RN(net54),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2921_ (.D(_0013_),
    .RN(net55),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2922_ (.D(_0014_),
    .RN(net54),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2923_ (.D(_0015_),
    .RN(net51),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2924_ (.D(_0016_),
    .RN(net51),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2925_ (.D(_0017_),
    .RN(net51),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2926_ (.D(_0018_),
    .RN(net51),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2927_ (.D(_0019_),
    .RN(net52),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2928_ (.D(_0020_),
    .RN(net55),
    .CLK(clknet_1_1__leaf_CLK),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2929_ (.D(_0021_),
    .RN(net48),
    .CLK(_0005_),
    .Q(\p_shaping_Q.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2930_ (.D(_0022_),
    .RN(net48),
    .CLK(_0005_),
    .Q(\p_shaping_Q.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2931_ (.D(\p_shaping_I.bit_in ),
    .RN(net57),
    .CLK(net42),
    .Q(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2932_ (.D(_0000_),
    .Q(\p_shaping_I.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2933_ (.D(\p_shaping_I.bit_in_1 ),
    .RN(net58),
    .CLK(net43),
    .Q(\p_shaping_I.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2934_ (.D(_0023_),
    .RN(net52),
    .CLK(clknet_1_0__leaf_CLK),
    .Q(\bit2symb.regi ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2935_ (.D(\Reg_Delay_Q.Out ),
    .RN(net49),
    .CLK(_0005_),
    .Q(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__latrnq_1 _2936_ (.D(_0002_),
    .Q(\p_shaping_Q.ctl_1 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2937_ (.D(\p_shaping_Q.bit_in_1 ),
    .RN(net49),
    .CLK(_0005_),
    .Q(\p_shaping_Q.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2938_ (.D(_0024_),
    .RN(net57),
    .CLK(net43),
    .Q(\p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 _2939_ (.D(_0025_),
    .RN(net57),
    .CLK(net43),
    .Q(\p_shaping_I.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input1 (.I(BitIn),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input2 (.I(EN),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(RST),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output4 (.I(net4),
    .Z(I[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output5 (.I(net5),
    .Z(I[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output6 (.I(net6),
    .Z(I[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output7 (.I(net7),
    .Z(I[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output8 (.I(net8),
    .Z(I[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output9 (.I(net9),
    .Z(I[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output10 (.I(net10),
    .Z(I[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(I[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(I[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net13),
    .Z(I[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(I[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(I[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(I[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(Q[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net18),
    .Z(Q[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(Q[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(Q[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(Q[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(Q[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(Q[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(Q[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(Q[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net26),
    .Z(Q[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(Q[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(Q[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(Q[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(addI[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(addI[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(addI[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(addI[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(addI[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(addI[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(addQ[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(addQ[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(addQ[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(addQ[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(addQ[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(addQ[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout42 (.I(_0004_),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout43 (.I(_0004_),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout44 (.I(net41),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout45 (.I(net40),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout46 (.I(net36),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout47 (.I(net35),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout48 (.I(net50),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout49 (.I(net50),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout50 (.I(net59),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout51 (.I(net53),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout53 (.I(net56),
    .Z(net53));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout54 (.I(net56),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout55 (.I(net56),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout56 (.I(net58),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout57 (.I(net58),
    .Z(net57));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout58 (.I(net59),
    .Z(net58));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout59 (.I(net3),
    .Z(net59));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_CLK (.I(CLK),
    .Z(clknet_0_CLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_0__f_CLK (.I(clknet_0_CLK),
    .Z(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_1_1__f_CLK (.I(clknet_0_CLK),
    .Z(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(BitIn));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_CLK_I (.I(CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(EN));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(RST));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2874__A1 (.I(\Reg_Delay_Q.In ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__I1 (.I(\Reg_Delay_Q.In ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__D (.I(\Reg_Delay_Q.Out ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2021__B (.I(\Reg_Delay_Q.Out ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1988__I (.I(\Reg_Delay_Q.Out ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1527__I (.I(\Reg_Delay_Q.Out ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout43_I (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout42_I (.I(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__CLK (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2935__CLK (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__CLK (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__CLK (.I(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__D (.I(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__D (.I(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__D (.I(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__D (.I(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__D (.I(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__D (.I(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__D (.I(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__D (.I(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__D (.I(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__D (.I(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__D (.I(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__D (.I(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__D (.I(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__D (.I(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__D (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2908__A1 (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2180__A1 (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2119__A1 (.I(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__D (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2913__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2824__A1 (.I(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A1 (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2616__I (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__B (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A1 (.I(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A3 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A3 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2617__A2 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A2 (.I(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A1 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__A1 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A1 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__B2 (.I(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A2 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__A1 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A1 (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2371__C (.I(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A2 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2001__A2 (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1778__I (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A2 (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1463__I (.I(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A1 (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__B (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A1 (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2373__I (.I(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A3 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2495__A1 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__B2 (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2375__I (.I(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A3 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2662__A3 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A2 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__A2 (.I(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__B (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2380__B (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A2 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2401__A1 (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__B (.I(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A3 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A3 (.I(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A1 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A2 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A1 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A1 (.I(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__B1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A1 (.I(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__A1 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A1 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A2 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__A1 (.I(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2566__I (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A1 (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A1 (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A1 (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2674__I (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A2 (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__B (.I(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A2 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A2 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__A2 (.I(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A2 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2392__A3 (.I(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A1 (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1552__I (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1480__I (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1465__I (.I(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A2 (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__B (.I(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__B2 (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2395__A2 (.I(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2880__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A2 (.I(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2550__A2 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2548__A2 (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__B (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__B (.I(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2718__I (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__B (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__C (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A2 (.I(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A3 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A2 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__A2 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A2 (.I(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2476__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A3 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__B (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2412__A1 (.I(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A3 (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2413__A2 (.I(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A1 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2670__I (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__B (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2419__B (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A2 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A2 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A2 (.I(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__B1 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A2 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__B1 (.I(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A4 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A3 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A2 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2428__A1 (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__B2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__B1 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2500__A2 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A3 (.I(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A3 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2531__A3 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2489__A3 (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2430__I (.I(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__B2 (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2659__I (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__C (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__A1 (.I(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__A1 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__B2 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A3 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A1 (.I(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__B (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2436__A2 (.I(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2588__I (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A1 (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__C (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A1 (.I(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A3 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A2 (.I(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A3 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2537__A3 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A1 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2441__A3 (.I(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A1 (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1821__B (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__B (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1473__A2 (.I(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A1 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A1 (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2446__I (.I(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A2 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A2 (.I(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A1 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2632__I (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A1 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2449__A2 (.I(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2571__C (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2509__B (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2451__A2 (.I(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__B (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1568__I (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1546__I (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1471__I (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__A2 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A1 (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__B (.I(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A3 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__B (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__A2 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A2 (.I(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A2 (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__A2 (.I(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2520__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2463__A2 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A3 (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__B (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2464__A4 (.I(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2470__I (.I(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A1 (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A1 (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__A1 (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2473__A1 (.I(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A1 (.I(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A2 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A1 (.I(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__B (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__A2 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A3 (.I(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A3 (.I(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1474__A2 (.I(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A2 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A2 (.I(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__A2 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__A2 (.I(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2758__A3 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A2 (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__B (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2486__B (.I(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2624__A3 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2488__A3 (.I(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A1 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A1 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__A1 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2490__A1 (.I(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A2 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A2 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__A2 (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1806__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1783__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1510__A1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A1 (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2544__I (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A1 (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A1 (.I(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A2 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2497__I (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2581__A1 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2572__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2508__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2504__A2 (.I(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__B (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__A2 (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__B (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1587__I (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1478__A1 (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2555__A3 (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2503__I (.I(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A3 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A3 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A4 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2511__A4 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2510__B2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1632__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A2 (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1477__I (.I(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2515__B (.I(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__A1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__A1 (.I(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__A2 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__B1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2678__A2 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__B1 (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A3 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2599__A3 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2521__A1 (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2523__B (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2522__A4 (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2806__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__B (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2529__A1 (.I(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__C (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__C (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__B2 (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1479__I (.I(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A1 (.I(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__B (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A3 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__A2 (.I(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2735__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2541__A1 (.I(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__C (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__B (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__B (.I(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__A2 (.I(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1925__I (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__C (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__B (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A1 (.I(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2626__A3 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2586__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2543__A2 (.I(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A2 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2579__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2552__A1 (.I(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__A2 (.I(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__A2 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A3 (.I(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A1 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2558__A2 (.I(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2630__C (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2610__A1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2577__B (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__B2 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2776__I (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A1 (.I(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A2 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2621__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1766__I (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A1 (.I(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__A2 (.I(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2768__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2570__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2592__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2567__A1 (.I(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A2 (.I(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2684__C (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2633__B (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2629__A2 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2582__A3 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__B (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A1 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1484__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__B (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2729__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2584__A1 (.I(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__A3 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A3 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2587__A3 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2696__I (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A1 (.I(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__B1 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__A2 (.I(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A1 (.I(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2679__B (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2666__I (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2642__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2597__C (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2644__A4 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2600__A1 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2649__B (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A4 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A3 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2601__A3 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A3 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A2 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1486__I (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2705__A3 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2607__A2 (.I(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2609__I (.I(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2712__A1 (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__B (.I(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__A1 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1670__I (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A2 (.I(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A1 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A2 (.I(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2739__I (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A1 (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__B (.I(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2731__I (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2638__C (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A1 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2620__A1 (.I(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__B1 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2619__A2 (.I(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A3 (.I(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2672__A4 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2658__A4 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2631__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2627__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A1 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__B (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1489__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2848__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2691__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2687__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A1 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2820__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2634__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2819__I (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2693__A1 (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2636__B (.I(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2711__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2710__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2706__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2637__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A1 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1490__A3 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2780__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2694__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2646__A1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2707__I (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__A2 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2647__A3 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1508__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2653__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2655__B (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2827__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A3 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2669__A2 (.I(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2778__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__C (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2660__A2 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1602__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A1 (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1492__I (.I(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__B (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2698__C (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2695__I (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A1 (.I(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__C (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__B (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2700__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2667__C (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2671__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2668__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1713__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__A1 (.I(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2730__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2689__A2 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2673__A3 (.I(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A1 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__C (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__B (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__B (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1494__I (.I(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2685__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2683__A2 (.I(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__B (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__C (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__A2 (.I(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2809__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A1 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2701__B2 (.I(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A3 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1731__A2 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1608__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1496__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2717__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2703__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2716__I (.I(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A3 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A4 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2726__A1 (.I(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A2 (.I(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2877__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A1 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2764__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2728__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2727__A2 (.I(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2801__I (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2767__B (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2734__B (.I(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2737__A2 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__A3 (.I(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2781__B2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2775__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2740__A1 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__C (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1718__I (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1506__B (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1500__B (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2886__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2872__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2743__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__B (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2746__A3 (.I(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1721__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1501__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2754__I (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2761__A1 (.I(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2763__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A2 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A2 (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__B (.I(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1597__A1 (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1503__I (.I(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__A1 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__B2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2894__B (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__B2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2777__B (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2796__B1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2783__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2793__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2785__A2 (.I(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2791__I (.I(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A1 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__A2 (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1505__I (.I(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A3 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2797__A2 (.I(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A2 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2888__B (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2803__B (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2805__A3 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2804__A2 (.I(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2833__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2812__A2 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1507__A2 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__B1 (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2823__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2864__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A1 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2843__A3 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2829__A2 (.I(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2850__A2 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2831__I (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2852__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2835__A2 (.I(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2857__A1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2853__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2841__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2842__I (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2847__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2846__A2 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2855__I (.I(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__B1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__B1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__A2 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2798__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2762__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__B (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A1 (.I(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2909__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2744__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2448__A1 (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1516__I (.I(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__S (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1534__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1524__A2 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1523__A1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2811__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2455__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1522__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__C (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1857__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1533__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2875__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2128__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1728__A1 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1531__A2 (.I(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2085__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1562__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1539__I (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__B (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1620__A1 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1541__I (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1875__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A1 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1759__A1 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1625__A2 (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1594__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1545__I (.I(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1574__A2 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1549__A1 (.I(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1792__A3 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A1 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1555__A2 (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1548__I (.I(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1841__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1668__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A1 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1551__A2 (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__B1 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1654__A3 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__A3 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1754__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A2 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B1 (.I(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__C (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A1 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1556__B2 (.I(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1583__A2 (.I(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A2 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__B (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A1 (.I(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__C (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A2 (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1560__I (.I(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A1 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__B (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1607__I (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1561__A2 (.I(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__B (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1687__I (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1565__I (.I(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1949__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__B (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1753__B2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1566__B (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__B (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__I1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A1 (.I(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1717__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1570__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1651__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A1 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A2 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A3 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1573__I (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1874__I (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1610__A3 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1870__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1650__I (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__B (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1576__C (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A1 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1627__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1801__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1644__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1580__A2 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__B (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1763__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1581__I (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__B1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__B2 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1582__B (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1958__A1 (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1639__I (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1586__I (.I(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__C (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A1 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__B (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1674__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1588__I (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1757__A2 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A3 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1621__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1590__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1892__B (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__C (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1593__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1986__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__C2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__B1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2039__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1888__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1598__B2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1656__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1599__A2 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1815__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1715__A1 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1601__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1847__B (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1603__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A2 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1814__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1605__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2083__A1 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1606__A3 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1619__B1 (.I(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__B (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A1 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1655__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1611__A2 (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__B (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1867__B (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__B (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1614__I (.I(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A1 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1817__A2 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1712__I (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__I0 (.I(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1694__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1669__B (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1631__A1 (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1616__I (.I(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__B (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1617__A2 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__A2 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1618__S (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__C (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1638__A2 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2161__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1626__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1755__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1647__I (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1628__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1623__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1737__I (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1624__A4 (.I(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1982__I (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1852__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1680__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__A2 (.I(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__B (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1630__B (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__A2 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__B2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2059__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__B (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__B1 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__B (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A3 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1960__A3 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1634__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1850__A1 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__B (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1635__B2 (.I(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1640__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1636__A2 (.I(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2057__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A1 (.I(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__A2 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1897__B (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1748__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1665__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1642__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2020__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1885__I (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1744__I (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1643__I (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__B (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1664__I (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__B1 (.I(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A1 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A2 (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1685__I (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1645__I (.I(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2015__C (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2005__C (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1915__B (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1646__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1785__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1761__A1 (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1649__I (.I(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1851__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1652__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__A2 (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__C (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1653__B (.I(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__C (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1725__A2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1658__B2 (.I(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1661__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2159__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__C (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2053__B2 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1702__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__B2 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A1 (.I(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2013__A3 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A3 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1673__A2 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1984__A2 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1709__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2075__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1965__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1672__A2 (.I(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2072__I (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__B2 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1675__A1 (.I(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1916__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__A2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1890__B (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1707__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1677__I (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A1 (.I(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A1 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1679__A2 (.I(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1802__A1 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__A2 (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1849__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A1 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__S0 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1682__I (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2905__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__B (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A1 (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1684__B (.I(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1690__B1 (.I(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A1 (.I(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1774__I (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1735__I (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1688__A1 (.I(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__A3 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1689__A2 (.I(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1752__A2 (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1691__B (.I(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1739__I (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1695__A2 (.I(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__B2 (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1697__B (.I(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__B1 (.I(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A1 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1699__A2 (.I(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2073__B (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__B1 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1700__B2 (.I(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A2 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1701__A3 (.I(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__C (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__C (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1930__A1 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1704__I (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__B2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__B2 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A1 (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__C (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__C (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__B (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1706__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2077__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2011__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1711__A1 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1907__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1768__A1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1708__B1 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2903__A1 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1710__A2 (.I(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1808__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1723__A2 (.I(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__C (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A2 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A1 (.I(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2062__A1 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A3 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1906__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1720__A2 (.I(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__B (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1716__I (.I(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1797__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__B (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__A2 (.I(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1979__I (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1791__A1 (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1719__B (.I(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__B1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1722__A1 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A1 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1736__I0 (.I(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A1 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1835__B (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1834__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1732__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1966__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1853__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A1 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1734__A2 (.I(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1741__A2 (.I(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1961__A2 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1887__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__A1 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1740__A2 (.I(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1751__A3 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__B (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1743__A3 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__B (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1862__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1745__I (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2071__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1746__A1 (.I(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__C (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1749__I (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2907__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1750__A1 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2000__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A1 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__A2 (.I(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1948__A2 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1756__A1 (.I(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2061__A2 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__B1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__B1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__B (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1771__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1758__C (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1839__B (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1765__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1760__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__B (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1762__A1 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A3 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__A3 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1845__A3 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1764__A2 (.I(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1904__I (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1819__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1767__A1 (.I(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2076__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1901__A3 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1869__A2 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1770__A3 (.I(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A2 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1781__B1 (.I(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1873__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A1 (.I(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1899__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1789__B (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A1 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A2 (.I(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1963__A1 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__B (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1787__I (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1776__A3 (.I(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1803__A3 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1777__A2 (.I(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2898__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2897__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1900__A2 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1779__A1 (.I(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1877__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1780__B1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__B (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1973__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1784__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__C (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1974__A1 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__B2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__A2 (.I(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__B (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1818__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1790__A1 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__A2 (.I(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1978__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__A1 (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1788__C (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2904__A1 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__B (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A1 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1793__C (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1794__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1910__A1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A2 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__B1 (.I(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1858__A1 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1796__B2 (.I(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2046__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1813__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1800__A2 (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1928__A3 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1926__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1799__A2 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A1 (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1805__I (.I(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2051__C (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2009__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A1 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1807__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2118__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2080__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A1 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A3 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__A2 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1809__A4 (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1832__A4 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1811__A4 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1810__B2 (.I(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2084__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A1 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1816__A3 (.I(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2003__A3 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A1 (.I(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2014__A3 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__B1 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1822__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1863__A3 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1824__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1833__A3 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1826__B (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1825__A4 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1831__I (.I(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1914__A4 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1848__A4 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1838__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2040__B (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1840__A2 (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A3 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A1 (.I(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1980__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1946__A3 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1843__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1844__C (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1895__A4 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1886__A4 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1846__A1 (.I(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1861__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1860__A2 (.I(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1855__A2 (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2048__A1 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1854__A2 (.I(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1898__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1859__B1 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1856__A2 (.I(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2900__B2 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A1 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2012__A3 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1866__A3 (.I(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1913__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__B1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1959__B (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1952__A2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1868__B2 (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2010__A2 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__B1 (.I(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2114__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2087__A1 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1902__A2 (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1872__C (.I(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2899__B1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2022__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1912__A2 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1876__A1 (.I(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1989__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1931__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1878__A2 (.I(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1883__A4 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1879__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1882__I (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A1 (.I(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1891__B2 (.I(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1956__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1896__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1893__A2 (.I(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A1 (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1944__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1921__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1920__A2 (.I(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1903__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A2 (.I(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1924__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1923__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1905__A1 (.I(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2089__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1908__A2 (.I(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1918__A3 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1909__A3 (.I(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__I0 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1919__A1 (.I(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__A2 (.I(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2060__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2042__B2 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1929__A1 (.I(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1945__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1933__A2 (.I(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1942__I (.I(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1947__A2 (.I(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2120__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2006__A2 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A1 (.I(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1950__A2 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2136__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1951__A2 (.I(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__B2 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1968__A1 (.I(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2115__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2088__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1964__A3 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A3 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1967__B2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1971__A3 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1970__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1969__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1997__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1976__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1975__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2901__B2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__C (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__B2 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1981__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2113__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2074__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1983__A2 (.I(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2135__B (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2024__A2 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1985__B (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1987__B (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2029__B (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1998__A3 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1992__A3 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2121__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2047__A2 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2038__B (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2002__A4 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2055__I (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2008__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2036__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2019__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2018__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2017__S (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2143__B2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2127__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2025__A2 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2035__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2043__B (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2045__A2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2044__A3 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2049__A2 (.I(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2050__A2 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__B (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2056__A1 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2070__I (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2058__A3 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2063__A2 (.I(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2069__I (.I(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2139__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2095__C (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2078__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2079__S (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2906__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2160__B (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2126__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2086__A1 (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2091__A2 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2090__C (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2110__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2099__A2 (.I(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2117__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2116__A2 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2124__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2123__A2 (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2147__A2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2129__A3 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2134__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2138__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2137__A2 (.I(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2141__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2140__A2 (.I(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2178__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2168__A1 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2156__A2 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2142__A2 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2166__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2165__A1 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2157__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2144__A2 (.I(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2170__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2148__A2 (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2163__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2162__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2173__I (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2181__B (.I(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A2 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2192__A1 (.I(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A1 (.I(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A4 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A3 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2191__A2 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2549__B (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2329__I (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A2 (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2195__I (.I(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2513__B (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__C (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A1 (.I(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2202__I (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2200__A1 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2379__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2260__I (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2388__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1446__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2203__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2564__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A2 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A3 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2208__A3 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2893__A4 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2733__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2641__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A1 (.I(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2562__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2478__A1 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2207__A2 (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2501__B (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2426__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A1 (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2210__I (.I(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2559__I (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2554__S (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A1 (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2211__B (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2454__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2239__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2545__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2185__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2596__I (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2540__B (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2409__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A1 (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2774__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2393__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2381__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2372__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2249__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2216__I (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2613__I (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2460__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__B (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__A1 (.I(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2389__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2273__I (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2219__A2 (.I(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2404__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2331__I (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2236__A1 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A2 (.I(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A4 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__B2 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2244__B (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2225__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2266__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2254__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2228__I (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2224__A1 (.I(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2794__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A4 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__B1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__B1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A2 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2316__I (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2234__A1 (.I(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2538__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A1 (.I(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2484__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2233__A2 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2352__I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A2 (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1449__I (.I(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2680__B2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__A1 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2391__A2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2235__B2 (.I(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2518__C (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2429__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2237__I (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2682__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2590__B (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2477__A1 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2238__B2 (.I(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2411__A2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2307__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2339__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2336__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2283__I (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A1 (.I(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2865__B2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2849__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2747__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2306__A1 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2612__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2517__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__B (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2347__B (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A1 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2247__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2546__A1 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__B2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2400__C (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2248__B (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2766__A1 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__A2 (.I(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__B (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__B (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__B (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2250__I (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2516__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2362__I (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2443__A3 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2421__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2253__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2288__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2255__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2697__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__A2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A3 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__B2 (.I(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2676__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2561__B (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2369__I (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2257__C (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A2 (.I(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2442__A3 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__B (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2263__B (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2259__I (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2594__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2367__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A1 (.I(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2665__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2384__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2365__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2264__A2 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2271__I (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2262__A1 (.I(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2385__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2261__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2184__I (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A1 (.I(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2333__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__A3 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2425__B (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2298__A1 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2278__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2268__A3 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2825__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2639__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2311__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2269__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2563__A1 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2270__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2355__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2282__B1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2721__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__B (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2315__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2274__A2 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2741__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2732__A1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2568__A2 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2281__B1 (.I(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2458__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2376__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2317__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2277__I (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A3 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2512__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A1 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__A2 (.I(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2420__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2390__B (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A1 (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2280__B (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2258__I (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2204__A1 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2190__B (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1456__A2 (.I(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2450__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2382__C (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A1 (.I(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2499__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2435__B (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2427__A3 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A1 (.I(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2485__I (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A1 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2294__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2287__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2595__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A1 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__A2 (.I(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2722__A3 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__B1 (.I(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2589__A1 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2560__I (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2290__A2 (.I(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2720__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2498__A2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2408__A1 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2291__B2 (.I(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A1 (.I(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2481__B (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2403__B (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2340__I (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__A2 (.I(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2593__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2327__I (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2296__A2 (.I(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2487__C (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__A1 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__A3 (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2759__A1 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__B2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2299__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2514__C (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2433__A1 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2354__B (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2301__B2 (.I(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__B (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2302__B (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A1 (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2303__I (.I(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__B2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2305__A2 (.I(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2308__I (.I(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2799__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2765__C (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2611__A1 (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2310__I (.I(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2648__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2465__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2416__A1 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__A2 (.I(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2757__B (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2573__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2496__B (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2334__A1 (.I(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2891__A4 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2724__A3 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2214__A2 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1457__A4 (.I(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2439__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2407__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A1 (.I(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2351__A1 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2350__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2314__A2 (.I(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2494__A2 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2459__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2319__A1 (.I(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2681__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2675__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2618__A1 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A2 (.I(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2885__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2821__C (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2661__A1 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2318__A3 (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2479__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A1 (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2322__I (.I(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2493__A1 (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2444__B (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1515__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1458__I (.I(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2614__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2565__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2457__A1 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2323__A2 (.I(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2591__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2533__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2422__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2326__A2 (.I(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2547__A3 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2539__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2480__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2328__A2 (.I(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2622__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2536__A2 (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__B (.I(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2663__I (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2640__B (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2553__B (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2330__C (.I(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2868__A2 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2519__A1 (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1459__I (.I(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2492__A1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2394__A2 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2335__B1 (.I(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2828__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2770__B (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2654__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2397__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2736__B (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2688__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2585__B (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2535__B (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2461__C (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2445__B2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2341__I (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2845__B2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2822__A1 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2795__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__A2 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2690__A1 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2656__I (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2532__B (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2344__C (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2357__A1 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2773__A1 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2699__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2346__A2 (.I(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2664__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2423__A1 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2348__B (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2551__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2502__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2364__I (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2353__B (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2625__A2 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2356__I (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2396__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2358__A2 (.I(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2475__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2456__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2402__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2360__A2 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2760__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2719__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2483__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2363__A2 (.I(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1837__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1696__A2 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1557__A1 (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1462__I (.I(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__D (.I(\p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2447__A1 (.I(\p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1517__I (.I(\p_shaping_I.bit_in ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__D (.I(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2580__C (.I(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1512__I (.I(\p_shaping_I.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2912__A2 (.I(\p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2338__I (.I(\p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2241__A2 (.I(\p_shaping_I.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2937__D (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1917__B (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1724__I (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1525__I (.I(\p_shaping_Q.bit_in_1 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2082__I (.I(\p_shaping_Q.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1692__I (.I(\p_shaping_Q.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1666__I (.I(\p_shaping_Q.bit_in_2 ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2910__I1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2870__I0 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2890__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2882__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2876__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout59_I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output8_I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output17_I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output18_I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output19_I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output20_I (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2196__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1444__I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2223__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1450__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2220__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2198__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1454__I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2267__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1452__I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2265__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2193__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1448__I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout47_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout46_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1622__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1464__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1495__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1470__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1563__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1467__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout45_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout44_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__CLK (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2889__A2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2881__B1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2869__A2 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__CLK (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1589__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1579__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A2 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1476__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1577__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1559__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1498__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1475__I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1571__A2 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1543__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1487__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1460__I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1530__A1 (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1520__I (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2930__RN (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2929__RN (.I(net48));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout48_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout49_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__RN (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout54_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout55_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout53_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2931__RN (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2939__RN (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2938__RN (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1521__A2 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2933__RN (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout57_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout56_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout58_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout50_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2915__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2916__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2923__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2924__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2925__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2926__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2927__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2934__CLK (.I(clknet_1_0__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2914__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2917__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2918__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2919__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2920__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2921__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2922__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__2928__CLK (.I(clknet_1_1__leaf_CLK));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_507 ();
endmodule

