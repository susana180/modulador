magic
tech gf180mcuC
magscale 1 5
timestamp 1670198997
<< obsm1 >>
rect 672 1538 29839 28321
<< metal2 >>
rect 1344 29600 1400 29900
rect 4032 29600 4088 29900
rect 7056 29600 7112 29900
rect 9744 29600 9800 29900
rect 12768 29600 12824 29900
rect 15792 29600 15848 29900
rect 18480 29600 18536 29900
rect 21504 29600 21560 29900
rect 24192 29600 24248 29900
rect 27216 29600 27272 29900
rect 29904 29600 29960 29900
rect 0 100 56 400
rect 2688 100 2744 400
rect 5712 100 5768 400
rect 8400 100 8456 400
rect 11424 100 11480 400
rect 14112 100 14168 400
rect 17136 100 17192 400
rect 20160 100 20216 400
rect 22848 100 22904 400
rect 25872 100 25928 400
rect 28560 100 28616 400
<< obsm2 >>
rect 14 29570 1314 29600
rect 1430 29570 4002 29600
rect 4118 29570 7026 29600
rect 7142 29570 9714 29600
rect 9830 29570 12738 29600
rect 12854 29570 15762 29600
rect 15878 29570 18450 29600
rect 18566 29570 21474 29600
rect 21590 29570 24162 29600
rect 24278 29570 27186 29600
rect 27302 29570 29874 29600
rect 14 430 29946 29570
rect 86 350 2658 430
rect 2774 350 5682 430
rect 5798 350 8370 430
rect 8486 350 11394 430
rect 11510 350 14082 430
rect 14198 350 17106 430
rect 17222 350 20130 430
rect 20246 350 22818 430
rect 22934 350 25842 430
rect 25958 350 28530 430
rect 28646 350 29946 430
<< metal3 >>
rect 100 28560 400 28616
rect 29600 27216 29900 27272
rect 100 25872 400 25928
rect 29600 24192 29900 24248
rect 100 22848 400 22904
rect 29600 21504 29900 21560
rect 100 19824 400 19880
rect 29600 18480 29900 18536
rect 100 17136 400 17192
rect 29600 15792 29900 15848
rect 100 14112 400 14168
rect 29600 12768 29900 12824
rect 100 11424 400 11480
rect 29600 10080 29900 10136
rect 100 8400 400 8456
rect 29600 7056 29900 7112
rect 100 5712 400 5768
rect 29600 4032 29900 4088
rect 100 2688 400 2744
rect 29600 1344 29900 1400
<< obsm3 >>
rect 9 28530 70 28602
rect 430 28530 29951 28602
rect 9 27302 29951 28530
rect 9 27186 29570 27302
rect 29930 27186 29951 27302
rect 9 25958 29951 27186
rect 9 25842 70 25958
rect 430 25842 29951 25958
rect 9 24278 29951 25842
rect 9 24162 29570 24278
rect 29930 24162 29951 24278
rect 9 22934 29951 24162
rect 9 22818 70 22934
rect 430 22818 29951 22934
rect 9 21590 29951 22818
rect 9 21474 29570 21590
rect 29930 21474 29951 21590
rect 9 19910 29951 21474
rect 9 19794 70 19910
rect 430 19794 29951 19910
rect 9 18566 29951 19794
rect 9 18450 29570 18566
rect 29930 18450 29951 18566
rect 9 17222 29951 18450
rect 9 17106 70 17222
rect 430 17106 29951 17222
rect 9 15878 29951 17106
rect 9 15762 29570 15878
rect 29930 15762 29951 15878
rect 9 14198 29951 15762
rect 9 14082 70 14198
rect 430 14082 29951 14198
rect 9 12854 29951 14082
rect 9 12738 29570 12854
rect 29930 12738 29951 12854
rect 9 11510 29951 12738
rect 9 11394 70 11510
rect 430 11394 29951 11510
rect 9 10166 29951 11394
rect 9 10050 29570 10166
rect 29930 10050 29951 10166
rect 9 8486 29951 10050
rect 9 8370 70 8486
rect 430 8370 29951 8486
rect 9 7142 29951 8370
rect 9 7026 29570 7142
rect 29930 7026 29951 7142
rect 9 5798 29951 7026
rect 9 5682 70 5798
rect 430 5682 29951 5798
rect 9 4118 29951 5682
rect 9 4002 29570 4118
rect 29930 4002 29951 4118
rect 9 2774 29951 4002
rect 9 2658 70 2774
rect 430 2658 29951 2774
rect 9 1430 29951 2658
rect 9 1314 29570 1430
rect 29930 1314 29951 1430
rect 9 630 29951 1314
<< metal4 >>
rect 2224 1538 2384 28254
rect 9904 1538 10064 28254
rect 17584 1538 17744 28254
rect 25264 1538 25424 28254
<< obsm4 >>
rect 1022 1508 2194 27991
rect 2414 1508 9874 27991
rect 10094 1508 17554 27991
rect 17774 1508 25234 27991
rect 25454 1508 28882 27991
rect 1022 737 28882 1508
<< labels >>
rlabel metal3 s 100 8400 400 8456 6 BitIn
port 1 nsew signal input
rlabel metal2 s 22848 100 22904 400 6 CLK
port 2 nsew signal input
rlabel metal2 s 15792 29600 15848 29900 6 EN
port 3 nsew signal input
rlabel metal3 s 100 22848 400 22904 6 I[0]
port 4 nsew signal output
rlabel metal2 s 28560 100 28616 400 6 I[10]
port 5 nsew signal output
rlabel metal3 s 29600 1344 29900 1400 6 I[11]
port 6 nsew signal output
rlabel metal3 s 29600 18480 29900 18536 6 I[12]
port 7 nsew signal output
rlabel metal2 s 1344 29600 1400 29900 6 I[1]
port 8 nsew signal output
rlabel metal3 s 100 25872 400 25928 6 I[2]
port 9 nsew signal output
rlabel metal2 s 24192 29600 24248 29900 6 I[3]
port 10 nsew signal output
rlabel metal2 s 17136 100 17192 400 6 I[4]
port 11 nsew signal output
rlabel metal3 s 29600 21504 29900 21560 6 I[5]
port 12 nsew signal output
rlabel metal3 s 29600 4032 29900 4088 6 I[6]
port 13 nsew signal output
rlabel metal2 s 5712 100 5768 400 6 I[7]
port 14 nsew signal output
rlabel metal3 s 100 19824 400 19880 6 I[8]
port 15 nsew signal output
rlabel metal3 s 100 14112 400 14168 6 I[9]
port 16 nsew signal output
rlabel metal2 s 18480 29600 18536 29900 6 Q[0]
port 17 nsew signal output
rlabel metal2 s 27216 29600 27272 29900 6 Q[10]
port 18 nsew signal output
rlabel metal3 s 100 17136 400 17192 6 Q[11]
port 19 nsew signal output
rlabel metal3 s 29600 24192 29900 24248 6 Q[12]
port 20 nsew signal output
rlabel metal2 s 7056 29600 7112 29900 6 Q[1]
port 21 nsew signal output
rlabel metal2 s 0 100 56 400 6 Q[2]
port 22 nsew signal output
rlabel metal3 s 100 5712 400 5768 6 Q[3]
port 23 nsew signal output
rlabel metal3 s 29600 15792 29900 15848 6 Q[4]
port 24 nsew signal output
rlabel metal2 s 4032 29600 4088 29900 6 Q[5]
port 25 nsew signal output
rlabel metal3 s 100 2688 400 2744 6 Q[6]
port 26 nsew signal output
rlabel metal2 s 25872 100 25928 400 6 Q[7]
port 27 nsew signal output
rlabel metal2 s 21504 29600 21560 29900 6 Q[8]
port 28 nsew signal output
rlabel metal3 s 29600 7056 29900 7112 6 Q[9]
port 29 nsew signal output
rlabel metal2 s 2688 100 2744 400 6 RST
port 30 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 addI[0]
port 31 nsew signal output
rlabel metal2 s 11424 100 11480 400 6 addI[1]
port 32 nsew signal output
rlabel metal3 s 29600 10080 29900 10136 6 addI[2]
port 33 nsew signal output
rlabel metal2 s 14112 100 14168 400 6 addI[3]
port 34 nsew signal output
rlabel metal3 s 29600 27216 29900 27272 6 addI[4]
port 35 nsew signal output
rlabel metal2 s 29904 29600 29960 29900 6 addI[5]
port 36 nsew signal output
rlabel metal2 s 9744 29600 9800 29900 6 addQ[0]
port 37 nsew signal output
rlabel metal2 s 12768 29600 12824 29900 6 addQ[1]
port 38 nsew signal output
rlabel metal2 s 20160 100 20216 400 6 addQ[2]
port 39 nsew signal output
rlabel metal3 s 100 11424 400 11480 6 addQ[3]
port 40 nsew signal output
rlabel metal3 s 100 28560 400 28616 6 addQ[4]
port 41 nsew signal output
rlabel metal3 s 29600 12768 29900 12824 6 addQ[5]
port 42 nsew signal output
rlabel metal4 s 2224 1538 2384 28254 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 28254 6 vdd
port 43 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 28254 6 vss
port 44 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 28254 6 vss
port 44 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3990718
string GDS_FILE /home/urielcho/Proyectos_caravel/gf180nm/modulador/openlane/modulador/runs/22_12_04_18_07/results/signoff/OQPSK_PS_RCOSINE2.magic.gds
string GDS_START 359124
<< end >>

