* NGSPICE file created from OQPSK_PS_RCOSINE2.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffrnq_1 D RN CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__latrnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__latrnq_1 D E RN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

.subckt OQPSK_PS_RCOSINE2 BitIn CLK EN I[0] I[10] I[11] I[12] I[1] I[2] I[3] I[4]
+ I[5] I[6] I[7] I[8] I[9] Q[0] Q[10] Q[11] Q[12] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7]
+ Q[8] Q[9] RST addI[0] addI[1] addI[2] addI[3] addI[4] addI[5] addQ[0] addQ[1] addQ[2]
+ addQ[3] addQ[4] addQ[5] vdd vss
XTAP_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2106_ _1174_ _1175_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA_fanout56_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2037_ _1095_ _1100_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2939_ _0025_ net57 net43 p_shaping_I.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1757__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2706__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1479__I _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1942__I _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1920__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2881__B1 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2724_ _0418_ _0034_ _1389_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2655_ _0325_ _0335_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1606_ _0681_ _0683_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2586_ _0211_ _0222_ _0266_ _0268_ _0269_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_1537_ _0617_ _1537_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1468_ _0091_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1675__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1902__A2 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2593__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1969__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2394__A2 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2440_ _0110_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2371_ _0027_ _0029_ _0032_ _0033_ _0034_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2621__A3 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2909__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2707_ _0335_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2137__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2638_ _0272_ _0298_ _0095_ _0042_ _0302_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_59_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2569_ _0246_ _0247_ _0250_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1896__A1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2845__B1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2376__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1492__I _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2588__I _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1887__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1940_ _1013_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1811__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1871_ _0707_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2367__A2 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2423_ _1427_ _0090_ _0092_ _1319_ _0072_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_2354_ _1272_ _1328_ _1377_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2285_ _1258_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1802__B2 _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1577__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1802__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2358__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2076__C _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1487__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2070_ _1131_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1923_ _0981_ _0791_ _0919_ _0839_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1796__B1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1854_ _0814_ _0929_ _0930_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1785_ _0728_ _0649_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2760__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2406_ _1300_ _1265_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2337_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2512__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2268_ _1340_ _1300_ _1341_ _1323_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_65_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2199_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2640__B _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2200__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2019__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1490__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1570_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2776__I _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1848__A4 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2122_ _1160_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2053_ _1118_ _1119_ _1124_ _0744_ _1126_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_34_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2886_ _0439_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1906_ _0683_ _0793_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1837_ _0728_ _1443_ _0644_ _0406_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1768_ _0786_ _0844_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2733__A2 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1699_ _0659_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1590__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2421__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2724__A2 _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput20 net20 Q[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput7 net7 I[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput31 net31 addI[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2488__A1 _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2596__I _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2264__C _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2660__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2740_ _0435_ _0090_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2412__A1 _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2671_ _0349_ _0357_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2280__B _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1622_ net37 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1553_ _0632_ _0308_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1484_ _0243_ _0265_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2479__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2105_ _1140_ _1176_ _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2036_ _0828_ _1083_ _1092_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_fanout49_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2938_ _0024_ net57 net43 p_shaping_I.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2403__A1 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2190__B _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2921__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2869_ _0603_ net42 _0568_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2706__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2642__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1495__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2881__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1684__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2723_ _0365_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2654_ _1417_ _0318_ _0322_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2585_ _0211_ _0222_ _1419_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1605_ _0650_ _0684_ _0655_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1536_ _0604_ _0554_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1467_ net39 _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2872__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1675__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2624__A1 _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2019_ _0665_ _1083_ _1092_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1711__C _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2091__A2 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2370_ _1410_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_49_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2733__B _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2706_ _0317_ _0324_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_9_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2637_ _0317_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1593__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2568_ _0249_ _1350_ _1396_ _1421_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2499_ _0051_ _0159_ _1360_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1896__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1519_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2845__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2845__B2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2781__B1 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1887__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2553__B _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1870_ _0655_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2422_ _1391_ _1404_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2353_ _1430_ _1431_ _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1878__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2284_ _1296_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2827__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1999_ _1072_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1566__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1869__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2294__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2046__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1557__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2809__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1922_ _0962_ _0997_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1796__B2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1796__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1853_ _0729_ _0812_ _0854_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1784_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2405_ _0072_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2336_ _1311_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1720__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2267_ net33 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2198_ net32 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1588__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1711__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2019__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1498__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1490__A3 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1950__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1702__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2121_ _1191_ _1076_ _0762_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2052_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2885_ _1395_ _0579_ _0581_ _0217_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1905_ _0981_ _0838_ _0948_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1836_ _0912_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1767_ _0845_ _0810_ _0730_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1698_ _0427_ _0671_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2319_ _1392_ _1393_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2421__A2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput10 net10 I[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput21 net21 Q[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput8 net8 I[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2724__A3 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput32 net32 addI[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2488__A2 _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2660__A2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2561__B _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2670_ _0087_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1621_ _0669_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1552_ _0058_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1923__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1483_ _0254_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input3_I RST vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2479__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2104_ _1111_ _1138_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2736__B _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2035_ _1109_ net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2937_ p_shaping_Q.bit_in_1 net49 _0005_ p_shaping_Q.bit_in_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2868_ bit2symb.regi _1411_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2799_ _1386_ _0462_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1819_ _0845_ _0680_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1914__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1815__B _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1905__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2881__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2397__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2722_ _0026_ _0415_ _1364_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2653_ _0342_ net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2584_ _0267_ _0253_ _0258_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1604_ _0080_ _0674_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1535_ _0616_ _1535_/Z vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2310__I _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1466_ _0069_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2872__A2 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2018_ _0744_ _1083_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2624__A2 _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2220__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2095__C _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2890__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2379__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2551__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2705_ _0288_ _0286_ _0292_ _0336_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_2636_ _1416_ _0318_ _0322_ _0323_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1593__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2567_ _0248_ _0026_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2498_ _1364_ _1366_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1518_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1449_ _1302_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2845__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2781__B2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2934__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2421_ _1301_ _1325_ _0066_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2352_ _1302_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2283_ _1311_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1913__B _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2035__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1998_ _1051_ _1052_ _1067_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__1874__I _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2763__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2619_ _0303_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2638__C _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1784__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1557__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1921_ _0971_ _0974_ _0987_ _0996_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__1796__A2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1852_ _0696_ _0708_ _0693_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1783_ _0167_ _0544_ _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2404_ _1291_ _1260_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2335_ _1310_ _1387_ _1383_ _1414_ _1382_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2266_ _1293_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1720__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2197_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1484__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__B _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__B _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1950__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2120_ _0749_ _1024_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2051_ _0873_ _0975_ _0803_ _0885_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_13_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1904_ _0845_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2884_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2741__C _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1835_ _0688_ _0651_ _0810_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1766_ _0243_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1697_ _0297_ _0705_ _0775_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2318_ _1345_ _1394_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2249_ _1284_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1457__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2223__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2185__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput9 net9 I[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput22 net22 Q[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 addI[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput11 net11 I[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2379__B _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2488__A3 _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2660__A3 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1620__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1620_ _0620_ _0427_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1551_ _0351_ _0630_ _0406_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__1923__A2 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1482_ _0091_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2103_ _1111_ _1138_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2034_ _1102_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2308__I _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2936_ _0002_ _2936_/E _2936_/RN p_shaping_Q.ctl_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2867_ _0567_ net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1611__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1818_ _0865_ _0896_ _0714_ _0210_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2798_ _0586_ _0496_ _0267_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1749_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1882__I _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1850__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1602__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1905__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1669__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1841__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2721_ _1348_ _1336_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2652_ _0336_ _0340_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2583_ _0224_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1603_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1534_ _0604_ _0599_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1465_ _0058_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2747__B _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout54_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2872__A3 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2017_ _1047_ _1084_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2624__A3 _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1832__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2919_ _0011_ net54 clknet_1_1__leaf_CLK net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1826__B _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1899__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1787__I _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2379__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2000__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1814__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2704_ _0344_ _0397_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2635_ _1312_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2566_ _0053_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2497_ _0172_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1517_ p_shaping_I.bit_in _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1448_ net34 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2058__A1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2533__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2049__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1811__A4 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2420_ _1354_ _1267_ _0070_ _1292_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2351_ _1391_ _1327_ _1321_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2282_ _1278_ _1330_ _1338_ _1344_ _1356_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_37_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2316__I _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2460__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1997_ _1034_ _1050_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2763__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2618_ _1394_ _1365_ _0094_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2549_ _0227_ _0228_ _1261_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2690__A1 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1920_ _0971_ _0974_ _0987_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2442__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1851_ _0729_ _0502_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1782_ _0610_ _0613_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2403_ _1305_ _0070_ _1369_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2334_ _1388_ _1397_ _1409_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2265_ net34 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2196_ net30 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1484__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2433__A1 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1885__I _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2924__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2921__D _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1818__C _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2736__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1834__B _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2672__A1 _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2727__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2050_ _1082_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1903_ _0976_ _0977_ _0978_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2883_ _0278_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1834_ _0232_ _0810_ _0644_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1765_ _0243_ _0838_ _0645_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1696_ _0727_ _1443_ _0620_ _0688_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2317_ _1351_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2248_ _1317_ _1251_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2916__D _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2654__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2179_ _1235_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1457__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput34 net34 addI[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput12 net12 I[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 Q[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__1696__A2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2893__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1550_ _0623_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_1481_ _0232_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1923__A3 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2102_ _1102_ _1139_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2033_ _1103_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_47_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2935_ Reg_Delay_Q.Out net49 _0005_ p_shaping_Q.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2866_ _1415_ _0082_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1611__A2 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1817_ _0047_ _0694_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2797_ _0238_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_7_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1748_ _0721_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1679_ _0756_ _0757_ _0638_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2875__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2627__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__A1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1841__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2720_ _1364_ _1366_ _0249_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2651_ _0286_ _0293_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1602_ _0351_ _0406_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2582_ _0169_ _0261_ _0263_ _0264_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1533_ _0609_ _0554_ _0615_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1464_ net37 _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2857__A1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2016_ _1086_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA_fanout47_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2918_ _0010_ net53 clknet_1_1__leaf_CLK net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2849_ _1315_ _0462_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__1899__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2848__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2076__A2 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2000__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2551__A3 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1978__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1814__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2703_ _0386_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_9_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2634_ _0320_ _0321_ _0315_ _0316_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2565_ _1345_ _1401_ _0073_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1516_ _0592_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1750__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2496_ _0170_ _0171_ _1388_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1447_ net47 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2924__D _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1837__B _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__B1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2049__A2 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1980__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1732__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2350_ _1299_ _1391_ _1429_ _1353_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2281_ _1345_ _1349_ _1350_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2288__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1799__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2460__A2 _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1996_ _1071_ net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1971__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2617_ _0038_ _0030_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1723__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2548_ _0037_ _0066_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2919__D _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2479_ _1399_ _1254_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2451__A2 _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2203__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2442__A2 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2580__C p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1850_ _0714_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1781_ _0687_ _0847_ _0849_ _0856_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2402_ _1250_ _1440_ _1331_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2333_ _1412_ _1338_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2264_ _1332_ _1333_ _1336_ _1337_ _1262_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_2195_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2681__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2327__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2433__A2 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1979_ _0797_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2736__A3 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1944__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2237__I _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2700__I _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2360__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1902_ _0276_ _0949_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2882_ _0418_ net2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1833_ _0824_ _0889_ _0903_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1926__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1764_ _0831_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1695_ _0635_ _0773_ _0178_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2351__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2316_ _1297_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2247_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2178_ _1211_ _1234_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1917__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput13 net13 I[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2590__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 Q[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 addI[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1908__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2430__I _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2581__A1 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1480_ _0058_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2101_ _1103_ _1107_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2032_ _1069_ _1105_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2914__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2934_ _0023_ net52 clknet_1_0__leaf_CLK bit2symb.regi vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_15_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2865_ _0559_ _0563_ _0566_ _0520_ _1315_ net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1816_ _0618_ _0893_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2796_ _0412_ _0228_ _0480_ _0475_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__2572__A1 _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1747_ _0742_ _0822_ _0825_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2340__I _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1914__A4 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1678_ _0731_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2496__B _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2927__D _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2563__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2250__I _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2315__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2937__CLK _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__A2 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2650_ _0208_ _0337_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_12_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1601_ _0675_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2581_ _0173_ _0180_ _0184_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1532_ _0554_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1463_ _0036_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2306__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input1_I BitIn vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2015_ _1087_ _1088_ _1089_ _0725_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2917_ _0009_ net54 clknet_1_1__leaf_CLK net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2848_ _0320_ _0549_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2070__I _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2545__A1 _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2779_ _0078_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2775__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2702_ _0387_ _0394_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2633_ _0578_ _0255_ _0263_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2564_ _0026_ _1271_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1515_ _1400_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2495_ _0039_ _0041_ _0037_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1446_ _1269_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2058__A3 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_1_1__f_CLK clknet_0_CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2766__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__A1 _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1741__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2757__A1 _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1980__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1732__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2280_ _1334_ _1352_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1799__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1995_ _1068_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2613__I _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2616_ _0028_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1971__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2547_ _1399_ _1297_ _1406_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2478_ _1274_ _0090_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1723__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2935__D Reg_Delay_Q.Out vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2203__A3 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2679__B _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1478__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2690__A3 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2442__A3 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1780_ _0818_ _0846_ _0858_ _0661_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_2401_ _0043_ _1257_ _0067_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2332_ _1410_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2263_ _1250_ _1287_ _1331_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_1_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2194_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1512__I p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1978_ _0866_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1944__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2499__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2121__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1699__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2360__A2 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1623__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2881_ _0248_ _0576_ net42 _0577_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_1901_ _0746_ _0683_ _0848_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1832_ _0828_ _0843_ _0875_ _0888_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_30_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1763_ _0660_ _0832_ _0837_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1694_ _0695_ _0652_ _0692_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1926__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2351__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2315_ _1253_ _1348_ _1347_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2246_ _1346_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2338__I p_shaping_I.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2177_ _1243_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1457__A4 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1862__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1618__S _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1917__A2 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2801__I _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput25 net25 Q[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput14 net14 I[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2590__A2 _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2022__B _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput36 net36 addQ[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2893__A3 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1853__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1605__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1908__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2333__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2100_ _1144_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_39_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2031_ _1073_ _1104_ _1021_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1844__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2933_ p_shaping_I.bit_in_1 net58 net43 p_shaping_I.bit_in_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2864_ _0529_ _0564_ _0565_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1946__B _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1815_ _0622_ _0680_ _0667_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_30_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2795_ _1405_ _1422_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1746_ _0824_ _0806_ _0821_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2572__A2 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1677_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1780__B1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2777__B _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2229_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2088__A1 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2012__A1 _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2563__A2 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2315__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2618__A3 _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1826__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1600_ _0628_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2003__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2580_ _0034_ _0234_ _0262_ p_shaping_I.bit_in_1 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1531_ _0604_ _0612_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1462_ _1443_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1817__A1 _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2014_ _0797_ _1059_ _0900_ _1088_ _1087_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__2616__I _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2490__A1 _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1832__A4 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1520__I net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2916_ _0008_ net52 clknet_1_0__leaf_CLK Reg_Delay_Q.Out vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2847_ _0321_ _0547_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2793__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2778_ _0348_ _0472_ _0473_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__2545__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1729_ _0481_ _0502_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1753__B1 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1808__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A1 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2233__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2261__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2224__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2701_ _0348_ _0226_ _0392_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2632_ _0120_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2563_ _1343_ _0244_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1514_ _0578_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2494_ _1297_ _1392_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1515__I _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1445_ _1258_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout52_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2927__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2766__A2 _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2684__C _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2930__RN net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2454__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2757__A2 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2693__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2445__B2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2445__A1 _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1994_ _1011_ _1017_ _1069_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2615_ _1402_ _1405_ _1421_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1971__A3 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1708__B1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2546_ _1319_ _0225_ _0110_ _0131_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2477_ _1308_ _0150_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_18_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2436__A1 _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2427__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2442__A4 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1758__C _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2400_ _1317_ _0065_ _0066_ _1319_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2331_ _1291_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2262_ _1334_ _1270_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2193_ net34 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2681__A4 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1977_ _1051_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1684__B _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2529_ _0206_ _0165_ _0183_ _0186_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_0_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2672__A4 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2409__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1632__A2 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1699__A2 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2648__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2820__A1 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2880_ _0574_ _0065_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1900_ _0756_ _0857_ _0712_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1831_ _0909_ net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1762_ _0839_ _0639_ _0748_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__1926__A3 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1693_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2314_ _1390_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2245_ _1266_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2639__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2176_ _1225_ _1226_ _1237_ _1239_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_38_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__B _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2811__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput15 net15 I[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput37 net37 addQ[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput26 net26 Q[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2893__A4 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1853__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1605__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1608__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2869__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2030_ _1021_ _1073_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2932_ _0000_ _2932_/E _2932_/RN p_shaping_I.ctl_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__latrnq_1
X_2863_ _0532_ _0551_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1814_ _0265_ _0684_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2794_ _1295_ _1326_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1745_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1676_ _0727_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1780__B2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1780__A1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2228_ _1293_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2088__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2159_ _0743_ _1126_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1599__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2796__B1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2259__I _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1523__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1762__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1530_ net48 p_shaping_Q.ctl_1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1461_ _1432_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2597__C _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1817__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2013_ _0667_ _0792_ _0748_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2915_ _0007_ net52 clknet_1_0__leaf_CLK Reg_Delay_Q.In vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2632__I _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2846_ _0049_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2777_ _0241_ _0474_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1753__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1728_ _0612_ _0664_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1753__B2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1659_ _0718_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1808__A2 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2481__A2 _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2233__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1867__B _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2536__A3 _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2698__B _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2700_ _0356_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1983__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2631_ _0310_ _0313_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2562_ _1274_ _0225_ _0111_ _0242_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1513_ _0570_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_2493_ _1400_ _0119_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_4_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1444_ net30 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2160__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout45_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2463__A2 _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2362__I _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1974__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2829_ _0525_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1706__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__B _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout50 net59 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1717__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2390__A1 _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1616__I _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2142__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1993_ _0961_ _1010_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1956__A1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2614_ _1401_ _0298_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XANTENNA__1708__B2 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2545_ _0053_ _1280_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2476_ _0075_ _0149_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2436__A2 _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1947__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2675__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2267__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2427__A2 _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1635__B1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2363__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2330_ _1402_ _1405_ _1407_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1790__B _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2261_ _1335_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2917__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2115__B2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2115__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2192_ _1251_ _1257_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1976_ _1034_ _1050_ _0723_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1965__B _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1929__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2528_ _0148_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2459_ _1392_ _0131_ _0042_ _0073_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_56_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1859__C _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2648__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2820__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2281__B1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1830_ _0826_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2584__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1761_ _0728_ _0319_ _0287_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1692_ p_shaping_Q.bit_in_2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2313_ _1289_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2639__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2244_ _1253_ _1270_ _1292_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2175_ _1225_ _1226_ _1237_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__B1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__B _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1959_ _0813_ _0876_ _0945_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput38 net38 addQ[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 Q[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput16 net16 I[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2869__A2 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2931_ p_shaping_I.bit_in net57 net42 p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_15_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2862_ _0532_ _0551_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2793_ _0471_ _0484_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1813_ _0833_ _0876_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1744_ _0722_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1675_ _0753_ _0672_ _0619_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2227_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2158_ _1225_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2089_ _0777_ _0984_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1599__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2796__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2796__B2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2548__A1 _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2012__A3 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1872__C _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1444__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2720__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2539__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2003__A3 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1762__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1460_ net46 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2711__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2894__B _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2012_ _0047_ _0730_ _0943_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_23_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2778__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2914_ _0006_ net53 clknet_1_1__leaf_CLK p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_12_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2845_ _0475_ _1375_ _0304_ _1422_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2776_ _0240_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1727_ _0781_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1753__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1658_ _0719_ _0720_ _0723_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1589_ net44 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2698__C _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2630_ _1359_ _0314_ _0315_ _0316_ _0239_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__1983__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1793__B _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2561_ _0241_ _0040_ _1329_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1512_ p_shaping_I.bit_in_1 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2492_ _1414_ _0059_ _0060_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_4_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2160__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2828_ _1417_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2759_ _1375_ _0390_ _0455_ _0388_ _0356_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_2_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output19_I net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout51 net53 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1965__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1717__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2390__A2 _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2142__A2 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1788__B _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1653__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1992_ _1021_ _1053_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_20_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1956__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1807__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2613_ _1286_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2544_ _0169_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1708__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2905__A1 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2381__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2475_ _1440_ _1303_ _1403_ _0039_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_55_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2373__I _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1947__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2124__A2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1452__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2675__A3 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1883__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2427__A3 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1635__B2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2283__I _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2060__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2899__B1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2363__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2260_ _1267_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_34_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2115__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2191_ _1253_ _1254_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2910__I1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1626__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__B _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2193__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1975_ _1034_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2051__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2527_ _0205_ net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2354__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2458_ _1301_ _1351_ _1353_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_29_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2389_ _0053_ _1287_ _0054_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_28_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1617__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2831__I _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2042__A1 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2042__B2 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2278__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2648__A3 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1856__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1760_ _0766_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1691_ _0745_ _0720_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2312_ _1324_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2243_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2174_ _1218_ _1223_ _1238_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2137__B _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__B _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2024__B2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1958_ _0665_ _1030_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1889_ _0893_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput28 net28 Q[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput17 net17 Q[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput39 net39 addQ[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_29_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1838__A1 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2318__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2930_ _0022_ net48 _0005_ p_shaping_Q.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2254__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2861_ _0561_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2006__A1 _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2792_ _0463_ _0467_ _0468_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_7_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1812_ _0664_ _0820_ _0611_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1743_ _0743_ _0806_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1674_ _0667_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2226_ _1346_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2157_ _1212_ _1213_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2493__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2088_ _0762_ _1039_ _1157_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_34_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2796__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2548__A2 _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2330__B _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2720__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2484__A1 _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1460__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2236__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2539__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1762__A3 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2711__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2011_ _0785_ _1085_ _0619_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2475__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2475__B2 _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2913_ _0025_ _0600_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2844_ _0530_ _0532_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2775_ _0435_ _0388_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1726_ _0802_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1545__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1657_ _0726_ _0733_ _0734_ _0735_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_1588_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2209_ net47 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1992__A3 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2933__RN net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2457__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1680__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1793__C _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2560_ _1365_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2491_ _0118_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1511_ _0554_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2448__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2196__I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2620__A1 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2827_ _0345_ _0501_ _0526_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2758_ _0389_ _0153_ _0160_ _0279_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1709_ _0749_ _0633_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2689_ _0360_ _0363_ _0361_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2687__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2439__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout52 net53 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2678__A1 _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2850__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1653__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1788__C _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1991_ _1063_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2612_ _1317_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2543_ _0211_ _0222_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2474_ p_shaping_I.counter\[1\] _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2381__A3 _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2669__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout50_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1580__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2427__A4 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1635__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2513__B _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2899__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1571__A1 _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1643__I _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2739__I _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2190_ _1269_ _1255_ _1357_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1799__B _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1974_ _0863_ _1045_ _1046_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2526_ _0147_ _0203_ _0204_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__1562__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2457_ _1401_ _1393_ _0129_ _0104_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2388_ _1269_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1617__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2290__A2 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2042__A2 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1891__C _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2559__I _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1463__I _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2648__A4 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1856__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2805__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1792__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1690_ _0752_ _0754_ _0763_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2311_ _1313_ _1342_ _1281_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2242_ _1312_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2173_ _1241_ net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1847__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2024__A2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1548__I _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1957_ _0745_ _0972_ _1031_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1888_ _0178_ _0677_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1783__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput18 net18 Q[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput29 net29 Q[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2509_ _0184_ _0118_ _0122_ _0185_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1838__A2 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2263__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2842__I _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1458__I _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2318__A3 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2860_ _0546_ _0560_ _0555_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1811_ _0666_ _0843_ _0875_ _0888_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_30_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2791_ _0490_ net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2006__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1765__A1 _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1742_ _0807_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1673_ _0746_ _0748_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2190__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1831__I _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2225_ _1292_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2156_ _1208_ _1211_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2493__A2 _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2087_ _0949_ _1159_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1987__B _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__B _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1756__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__A1 _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2330__C _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2484__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1897__B _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2236__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1651__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2010_ _0656_ _0947_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2912_ _0206_ p_shaping_I.counter\[0\] _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1986__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2843_ _0025_ _0524_ _0529_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2774_ _0393_ _1283_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1725_ _0803_ _0737_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1656_ _0673_ _0678_ _0668_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1587_ _0178_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2163__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1910__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2208_ _1262_ _1267_ _1271_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_26_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2139_ _1145_ _0672_ _1160_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_14_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1901__A1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1471__I _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1968__A1 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2490_ _0163_ _0164_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1510_ _0167_ _0544_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2448__A2 _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2826_ _0501_ _0526_ _0425_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2384__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2757_ _0105_ _0195_ _1388_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2688_ _1419_ _0359_ _0364_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1708_ _0629_ _0631_ _0786_ _0746_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_1639_ _0665_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2136__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2136__B2 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2439__A2 _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout53 net56 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xfanout42 _0004_ net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2611__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2127__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2678__A2 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2850__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1990_ _1064_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2611_ _1386_ _0260_ _0285_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2542_ _0214_ _0215_ _0220_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2473_ _0144_ _0126_ _0137_ _0146_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2118__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2669__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout43_I _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2841__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2670__I _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2809_ _0393_ _0472_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2357__A1 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1580__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1868__B1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2348__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2899__A2 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1571__A2 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1859__B1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2823__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1973_ _0862_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2525_ _0083_ _0142_ _0140_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2456_ _1440_ _1325_ _1318_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1562__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2387_ _1252_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__B _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1744__I _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2502__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2310_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2741__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2241_ _1311_ p_shaping_I.counter\[0\] _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2172_ _1238_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2485__I _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2930__CLK _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1956_ _0964_ _0969_ _0772_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1887_ _0690_ _0818_ _0660_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput19 net19 Q[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_2508_ _0169_ _0173_ _0180_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2732__A1 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2439_ _1390_ _0109_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2799__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2344__B _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1739__I _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1649__I _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1810_ _0666_ _0843_ _0875_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2790_ _0486_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1741_ _0764_ _0815_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1765__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1672_ _0749_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2224_ _1293_ _1263_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2155_ _1224_ net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2086_ _1158_ _1121_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1939_ _1014_ _0907_ _1012_ _0957_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__2705__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1508__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2074__B _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2911_ _0598_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2842_ _0543_ net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2773_ _1425_ _0303_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1724_ p_shaping_Q.bit_in_1 _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1655_ _0687_ _0690_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1586_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2163__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2207_ _1273_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_66_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2138_ _1084_ _1206_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2069_ _1142_ net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1901__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2532__B _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2393__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1959__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2825_ _0503_ _1342_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2908__A1 _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2756_ _0452_ _0443_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2687_ _0320_ _0376_ _0378_ _0266_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1707_ _0755_ _0649_ _0319_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2384__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1638_ _0666_ _0699_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2136__A2 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1569_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout43 _0004_ net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout54 net56 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2611__A3 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2678__A3 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1638__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2063__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1810__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1810__B2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2610_ _0239_ _0259_ _0206_ _0223_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2541_ _0216_ _0219_ _0028_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2472_ _0101_ _0103_ _0123_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_5_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1877__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1801__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2808_ _0473_ _0476_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2739_ _0299_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1868__B2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1868__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1883__A4 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2347__B _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2045__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1477__I _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2348__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1556__B1 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1859__B2 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2520__A2 _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2036__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1972_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2587__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2524_ _0201_ _0202_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2455_ _0603_ _0127_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2386_ _0051_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__2511__A2 _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2805__A3 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2018__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1792__A3 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2540__B _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2741__A2 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2240_ p_shaping_I.counter\[1\] _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2171_ _1218_ _1223_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1670__I _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2257__B2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2009__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1955_ _1023_ _1027_ _1028_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1886_ _0716_ _0779_ _0842_ _0922_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2507_ _0570_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2732__A2 _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2438_ _1361_ _1255_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2369_ _1329_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2248__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2799__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2344__C _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2420__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2420__B2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2487__A1 _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2239__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2535__B _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_7_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1740_ _0817_ _0818_ _0221_ _0635_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1665__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1671_ _0705_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2223_ net31 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2478__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2154_ _1218_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2085_ _0618_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1938_ _0830_ _0904_ _0905_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1869_ _0675_ _0848_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2641__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2090__B _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2920__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2910_ bit2symb.regi net1 _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2841_ _0538_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2772_ _0463_ _0469_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2396__B1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1723_ _0783_ _0790_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1654_ _0646_ _0629_ _0631_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1585_ p_shaping_Q.counter\[1\] _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2206_ _1256_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2137_ _1084_ _1206_ _0823_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2068_ _1139_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2918__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1901__A3 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2614__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2393__A3 _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1656__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2824_ _0025_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2755_ _0424_ _0433_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2686_ _0235_ _0236_ _0377_ _0184_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1706_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1637_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1568_ _0124_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1499_ _0427_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1895__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2633__B _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout55 net56 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout44 net41 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1886__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1638__A2 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2063__A2 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2540_ _1347_ _0218_ _1282_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2471_ _1314_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1574__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1801__A2 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2807_ _0500_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2738_ _0424_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2669_ _0345_ _0347_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1868__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__A2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1707__B _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1556__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1556__B2 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1859__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2257__C _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2036__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1668__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1971_ _0883_ _0933_ _1044_ _0608_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__2587__A3 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2523_ _0144_ _0187_ _0188_ _0199_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2454_ _1279_ _1309_ _0077_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2385_ _1335_ _1290_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2511__A3 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 BitIn net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2630__C _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2202__I _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2077__C _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2018__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1777__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2821__B _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2170_ _1214_ _1217_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2257__A2 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1900__B _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1954_ _0963_ _0970_ _1029_ _0772_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1768__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1885_ _0722_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2506_ _0166_ _0168_ _0181_ _0182_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2437_ _1353_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2368_ _0031_ _1393_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2299_ _1362_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2248__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1759__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2420__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2641__B _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1771__I _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2411__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1670_ _0297_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2478__A2 _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2222_ _1290_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2153_ _1173_ _1179_ _1219_ _1221_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1630__B _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2084_ _0894_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1937_ _0742_ _0822_ _0825_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2402__A2 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1868_ _0866_ _0676_ _0944_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2705__A3 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2166__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1799_ _0729_ _0877_ _0853_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2636__B _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1766__I _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2090__C _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2546__B _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2880__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2840_ _0486_ _0489_ _0515_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_2771_ _0467_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2396__B2 _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1722_ _0799_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1653_ _0647_ _0697_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2699__A2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1584_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2205_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2456__B _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout59_I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2136_ _0687_ _1026_ _1205_ _0783_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2067_ _1102_ _1108_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1586__I _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2139__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2210__I _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2614__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1496__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2302__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1736__S0 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2853__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2823_ _0520_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2754_ _0451_ net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1705_ _0761_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2685_ _0370_ _0374_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1636_ _0706_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1567_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2541__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1498_ net45 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1895__A3 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2119_ _0022_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout56 net58 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xfanout45 net40 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2780__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1583__A2 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2532__A1 _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1886__A3 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2835__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2470_ _0143_ net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1574__A2 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2523__A1 _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2933__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2734__B _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1801__A3 _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2806_ _0206_ _0505_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2737_ _0425_ _0431_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2762__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2668_ _0349_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1619_ _0668_ _0679_ _0686_ _0691_ _0698_ _0673_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_4
XANTENNA__2514__B2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2514__A1 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2599_ _0127_ _0136_ _0197_ _0602_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_59_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2695__I _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1774__I _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1970_ _0994_ _1044_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2522_ _1312_ _0187_ _0188_ _0199_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__2744__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2453_ _0101_ _0103_ _0123_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2384_ _1333_ _1271_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2511__A4 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 EN net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_56_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2680__B1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1594__I _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2735__A1 _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1710__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1474__A1 _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__B1 _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1777__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2821__C _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2726__B2 _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2726__A1 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__B _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1953_ _1023_ _1027_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1884_ _0939_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2303__I _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2505_ _0578_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2436_ _0105_ _0106_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2459__B _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2367_ _1332_ _0030_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2298_ _1341_ _1302_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1456__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1589__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1931__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1695__A1 _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2221_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2152_ _1181_ _1182_ _1200_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2083_ _0685_ _0795_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1989__A2 _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1936_ _1012_ _0957_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2461__C _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1610__A1 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1867_ _0747_ _0416_ _0693_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
X_1798_ _0634_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1913__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2419_ _1381_ _1437_ _0087_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1821__B _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2371__C _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1601__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2157__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2770_ _0360_ _0465_ _1417_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2396__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1721_ _0764_ _0449_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1652_ _0729_ _0730_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__2148__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1583_ _0619_ _0636_ _0642_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__1692__I p_shaping_Q.bit_in_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2204_ _1357_ _1302_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2135_ _0746_ _0817_ _1060_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2066_ _1074_ _1101_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2084__A1 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1919_ _0988_ _0887_ _0994_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2899_ _0756_ _0576_ _0952_ _0590_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2139__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2311__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2382__B _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2870__I0 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1822__A1 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2550__A2 _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2302__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__A1 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1687__I _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2822_ _1422_ _0305_ _0521_ _0240_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2753_ _0447_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1704_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2684_ _0182_ _0255_ _0375_ _0263_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1635_ _0707_ _0710_ _0711_ _0712_ _0714_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1566_ _0243_ _0628_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1497_ _0406_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1895__A4 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2118_ _0886_ _1188_ _1126_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2049_ _0894_ _1120_ _1122_ _1055_ _0782_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__2057__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout46 net36 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout57 net58 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_13_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1886__A4 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2296__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2048__A1 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2599__A2 _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2805_ _0345_ _0501_ _0504_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2736_ _0345_ _0347_ _0431_ _1419_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2762__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2667_ _0352_ _0354_ _0355_ _0356_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1618_ _0694_ _0647_ _0697_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__2514__A2 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2598_ _0275_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1549_ _0625_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2216__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2450__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1556__A3 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2441__A1 _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2521_ _0197_ _0198_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2452_ _0101_ _0103_ _0123_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2383_ _0570_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput3 RST net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2680__B2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1875__I _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1808__C _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2719_ _0299_ _1442_ _0195_ _0105_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_10_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2655__B _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2671__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1474__A2 _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2423__B2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2423__A1 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2390__B _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2923__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1701__A3 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2565__B _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__A1 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1952_ _0734_ _0945_ _0640_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1883_ _0823_ _0938_ _0939_ _0956_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2717__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2504_ _0169_ _0173_ _0180_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2435_ _1250_ _0074_ _1360_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2459__C _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2366_ _1304_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2297_ _1281_ _1339_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1456__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1695__A2 _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1998__A3 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2939__RN net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2220_ net32 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2151_ _1202_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2082_ p_shaping_Q.bit_in_2 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_19_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1935_ _0911_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1866_ _0845_ _0047_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1797_ _0755_ _0796_ _0265_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2418_ _0086_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2874__A1 Reg_Delay_Q.In vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2349_ _1361_ _1255_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1601__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2865__B2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1840__A2 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2134__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1720_ _0791_ _0793_ _0795_ _0798_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_1651_ _0650_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1582_ _0647_ _0656_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2203_ _1268_ _1270_ _1254_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2134_ _1204_ net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2065_ _1111_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1918_ _0886_ _0980_ _0985_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2898_ _0857_ _0590_ _0591_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1849_ _0760_ _0330_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1898__A2 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2847__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2075__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2382__C _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2870__I1 Reg_Delay_Q.In vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1822__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1510__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1813__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2821_ _0389_ _1251_ _0353_ _1395_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2752_ _0398_ _0409_ _0448_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1703_ _0764_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1917__B p_shaping_Q.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2683_ _0370_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1634_ _0630_ _0713_ _0254_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1565_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1496_ _0395_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2117_ _0874_ _1186_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2048_ _0929_ _0833_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2914__D _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout47 net35 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
Xfanout58 net59 net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_13_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1740__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2296__A2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2048__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2599__A3 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1559__A1 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2287__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2039__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2804_ _0501_ _0504_ _0425_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2322__I _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2735_ _0216_ _0328_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2666_ _0281_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1617_ _0362_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2597_ _0033_ _0277_ _0280_ _0281_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1548_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1722__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1479_ _0210_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1789__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2450__A2 _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1713__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2269__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__A2 _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2520_ _0127_ _0136_ _0602_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2451_ _0121_ _0122_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2382_ _0035_ _0046_ _0586_ _1358_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2901__B1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2317__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2718_ _0073_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_10_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2649_ _0144_ _0260_ _0270_ _0285_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2499__A2 _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1840__B _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2120__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2671__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2423__A2 _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1951_ _0661_ _1026_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1882_ _0959_ net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2178__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2503_ _0179_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2434_ _1431_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2365_ _0028_ _1333_ _1271_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2350__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2296_ _1264_ _1372_ _1321_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2922__D _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1835__B _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1916__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A2 _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1907__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2580__A1 _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2150_ _1181_ _1182_ _1200_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2081_ _0962_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1843__B1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1934_ _0961_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1865_ _0899_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1610__A3 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1796_ _0860_ _0863_ _0873_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2417_ p_shaping_I.bit_in_2 _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2323__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2486__B _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2348_ _1399_ _1426_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2917__D _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2279_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2562__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2314__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2617__A2 _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1650_ _0655_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1581_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2553__A1 _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2305__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2202_ _1264_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2133_ _1201_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2064_ _1132_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_19_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2897_ _0857_ _0587_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1917_ _0860_ _0993_ p_shaping_Q.bit_in_1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_8_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1848_ _0760_ _0871_ _0925_ _0915_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_1779_ _0857_ _0724_ _0156_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2847__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2820_ _0120_ _0321_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2751_ _0344_ _0397_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_12_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1702_ _0744_ _0770_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2682_ _1308_ _0371_ _0372_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__2774__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1633_ _0632_ _0648_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1564_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1495_ net38 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2829__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1501__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2116_ _1048_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout57_I net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2047_ _0866_ _1076_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2055__I _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout48 net50 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xfanout59 net3 net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2930__D _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2765__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2517__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1740__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1559__A2 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2508__A1 _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1731__A2 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1979__I _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2803_ _0472_ _0350_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2747__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2734_ _0426_ _0428_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2665_ _1333_ _0133_ _0352_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1970__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1616_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2596_ _1282_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1547_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1478_ _0178_ _0200_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_39_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2925__D _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1789__A2 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1961__A2 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1713__A2 _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2441__A3 _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2729__A1 _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2450_ _1358_ _0035_ _0046_ _0578_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_5_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1952__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2381_ _1412_ _1283_ _0045_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2901__A1 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2901__B2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2717_ _0386_ _0396_ _0380_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2648_ _1387_ _0260_ _0270_ _0285_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2579_ _0226_ _0229_ _0231_ _1410_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_19_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2120__A2 _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1631__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2662__A3 _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1950_ _1024_ _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1881_ _0911_ _0957_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_41_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2502_ _1433_ _0174_ _0175_ _0177_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2433_ _1377_ _0043_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__1689__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2364_ _1433_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2350__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2295_ _1298_ _1323_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2638__B1 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1861__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output20_I net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1852__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2644__A3 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2080_ _0886_ _1152_ _1126_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1843__A1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1933_ _0999_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1864_ _0611_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1795_ _0803_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2020__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2416_ _1387_ _0063_ _0081_ _0084_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2767__B _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2323__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2486__C _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2347_ _1252_ _1264_ _1318_ _1266_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2278_ _1341_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2087__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2626__A3 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2933__D p_shaping_I.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1598__B1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2011__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2314__A2 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2078__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1825__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1580_ _0658_ _0659_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__2553__A2 _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2305__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2079__S _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2201_ _1252_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2132_ _1173_ _1179_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2063_ _1096_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_19_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1816__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2241__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2896_ _0584_ _0571_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1916_ _0754_ _0990_ _0991_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1847_ _0628_ _0652_ _0682_ _0621_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2341__I _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1778_ _0036_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2928__D _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2480__A1 _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2783__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2535__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2299__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2750_ _0445_ _0446_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2681_ _0365_ _1394_ _0278_ _1295_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__2774__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1701_ _0772_ _0717_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1632_ _0427_ _0189_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1563_ net39 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1494_ _0373_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1505__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2115_ _0851_ _1039_ _1168_ _0783_ _1185_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_2046_ _0868_ _0876_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2336__I _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_10_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2214__A1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2879_ _0574_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2517__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1843__C _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2926__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2508__A2 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2444__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2802_ _0426_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2733_ _1273_ _0415_ _0356_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2664_ _0353_ _1426_ _0092_ _0095_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1615_ _0626_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2595_ _1363_ _0279_ _0176_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1546_ _0124_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2759__C _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1477_ _0189_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2683__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2029_ _1051_ _1052_ _1067_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2426__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2380_ _0038_ _0040_ _0042_ _0044_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2901__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2595__B _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2665__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1640__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2716_ _0410_ net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2647_ _0296_ _0325_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_2578_ _0184_ _0118_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1529_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2408__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1631__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1603__I _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1880_ _0826_ _0908_ _0906_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2501_ _0129_ _0176_ _1277_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2432_ _0088_ _0100_ _1416_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2335__B1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2886__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1689__A2 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2363_ _1363_ _1442_ _0026_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2609__I _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2294_ _1296_ _1362_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_2_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2638__B2 _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2638__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1861__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1669__B _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2877__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2629__A1 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2644__A4 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1852__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1489__B _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1843__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1932_ _1007_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1863_ _0663_ _0820_ _0902_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1794_ _0619_ _0872_ _0799_ _0800_ _0699_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__2113__B _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2415_ _1439_ _0062_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1952__B _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2346_ _1299_ _1425_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2339__I _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2277_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1834__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1598__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1598__B2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2562__A3 _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1770__A1 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1522__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2249__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2078__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2002__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1761__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2200_ _1264_ _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2131_ _1144_ _1172_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2062_ _0793_ _1133_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1915_ _0714_ _0927_ _0725_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2241__A2 p_shaping_I.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2895_ _0585_ _0588_ _0589_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1846_ _0922_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1777_ _0851_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__1752__A1 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2069__I _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2329_ _1261_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2480__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__C _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1743__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2299__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2707__I _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2680_ _0365_ _0278_ _1295_ _1305_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1700_ _0670_ _0774_ _0767_ _0776_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_1631_ _0695_ _0676_ _0373_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1734__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1562_ _0618_ _0449_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1493_ _0102_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2114_ _0949_ _0685_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_27_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2045_ _0988_ _1117_ _0862_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2214__A2 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2352__I _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1973__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2878_ _0575_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1829_ _0906_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2939__D _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2211__B _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2444__A2 _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2801_ _0429_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2732_ _1350_ _0092_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2663_ _1408_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1707__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1614_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2594_ _1332_ _0278_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1545_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1516__I _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2121__B _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1476_ net44 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2683__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1891__B1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2028_ _1013_ _1011_ _1016_ _1068_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_54_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2435__A2 _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2082__I p_shaping_Q.bit_in_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1946__A1 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2015__C _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2371__B2 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2123__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2114__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2665__A2 _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1928__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2715_ _0398_ _0409_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2646_ _0332_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2577_ _1359_ _0223_ _0239_ _0259_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1528_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2916__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1459_ _1411_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2408__A2 _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1919__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2592__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2344__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1855__B1 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2500_ _1260_ _0095_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2431_ _0088_ _0100_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2335__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2939__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2335__B2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2362_ _1322_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2293_ _1340_ _1300_ _1368_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2638__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2629_ _0120_ _0263_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2326__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1704__I _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2629__A2 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2868__A2 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1614__I _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1931_ _0941_ _0955_ _0611_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1862_ _0823_ _0938_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1793_ _0867_ _0869_ _0870_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2113__C _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2414_ _1415_ _0082_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_57_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2345_ _1296_ _1379_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1531__A2 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2276_ _1289_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1598__A2 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2547__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1770__A2 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2078__A3 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2265__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2235__B1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2538__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2002__A3 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1761__A2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2710__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2130_ _1183_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2061_ _0700_ _0835_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1816__A3 _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1914_ _0785_ _0871_ _0925_ _0915_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2777__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2894_ _0474_ _0581_ _0475_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2529__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1845_ _0717_ _0779_ _0842_ _0771_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1776_ _0809_ _0852_ _0853_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__1752__A2 _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2701__B2 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2701__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2328_ _1354_ _1406_ _1328_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2259_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2085__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2759__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1630_ _0491_ _0708_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1734__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1561_ _0638_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1492_ _0351_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2113_ _0943_ _1058_ _0713_ _1054_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_54_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2044_ _0994_ _1045_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_50_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2877_ _0418_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1828_ _0904_ _0905_ _0830_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1725__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1759_ _0624_ _0688_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__1489__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1712__I _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2029__B _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1964__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2913__A1 _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2141__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1622__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2718__I _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1652__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2800_ _0497_ _0498_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2731_ _0302_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2662_ _0033_ _0350_ _0040_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1613_ _0692_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2402__B _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2593_ _1372_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1544_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1707__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2904__A1 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2380__A2 _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1475_ net45 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout55_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1891__A1 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2027_ _1074_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1891__B2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2929_ _0021_ net48 _0005_ p_shaping_Q.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1946__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2123__A2 _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2426__A3 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1634__A1 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2273__I _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2114__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1873__A1 _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2822__B1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1928__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2714_ _0399_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2050__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2645_ _0601_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1527__I Reg_Delay_Q.Out vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2576_ _0224_ _0253_ _0258_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_59_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1527_ Reg_Delay_Q.Out _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_1458_ _1400_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2408__A3 _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1919__A2 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2592__A2 _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2344__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2647__A3 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1855__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2280__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2731__I _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2430_ _0099_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2335__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2361_ _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2292_ net47 _1339_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1846__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__B _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2628_ _0049_ _0236_ _0235_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2326__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2559_ _1278_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1837__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A1 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2014__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2565__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2253__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1930_ _0782_ _1001_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1861_ _0827_ _0924_ _0936_ _0937_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_42_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1792_ _0470_ _0692_ _0627_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_6_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2413_ _0064_ _0081_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1805__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2344_ _1367_ _1422_ _1378_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_2275_ _1288_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1819__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2492__A1 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2244__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1696__B _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2795__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2547__A2 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1770__A3 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1450__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2483__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1825__A4 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2929__CLK _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2235__B2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2235__A1 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2002__A4 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1761__A3 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2710__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2060_ _1002_ _0880_ _1078_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1913_ _0989_ _0944_ _0647_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2777__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2893_ _0393_ _0587_ _0030_ _1273_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2529__A2 _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2124__C _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1844_ _0660_ _0914_ _0916_ _0918_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_1775_ _0145_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2327_ _1372_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2701__A2 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2258_ _1357_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2465__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2189_ _1368_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2768__A2 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1743__A3 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2456__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2208__A1 _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1560_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1491_ _0069_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2112_ _0962_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2447__A1 p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2043_ _0765_ _1115_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2135__B _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2876_ net2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1827_ _0830_ _0904_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1758_ _0621_ _0833_ _0835_ _0775_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_1689_ _0765_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2914__RN net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2045__B _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2610__A1 _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1964__A3 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2429__A1 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2730_ _0087_ _0363_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2661_ _1395_ _0160_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1612_ _0643_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2592_ _0248_ _0213_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1543_ net46 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1474_ _0047_ _0156_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2668__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout48_I net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2026_ _1095_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2928_ _0020_ net55 clknet_1_1__leaf_CLK net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__1946__A3 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2859_ _0546_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2819__I _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output29_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1634__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1598__C _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2898__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1789__B _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2822__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2822__B2 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1625__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2713_ _0296_ _0402_ _0403_ _0407_ _0339_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__1928__A3 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2050__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2644_ _0127_ _0136_ _0197_ _0283_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_2575_ _0168_ _0255_ _0257_ _0182_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2889__B2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1526_ _0608_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1561__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1543__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1457_ _1280_ _1291_ _1313_ _1389_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__2510__B1 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2009_ _0885_ _1047_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1718__I _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2323__B _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1855__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2280__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1791__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2360_ _1390_ _1440_ _1290_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2291_ _1360_ _1363_ _1364_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2099__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2627_ _0310_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2558_ _0224_ _0238_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2489_ _1381_ _1437_ _0099_ _0086_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2369__I _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1509_ _0533_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1837__A2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2262__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1876__C _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1448__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1892__B _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2253__A2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1860_ _0827_ _0924_ _0936_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_14_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1791_ _0797_ _0788_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2412_ _0077_ _0079_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2343_ p_shaping_I.bit_in_2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2274_ _1347_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1819__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2492__A2 _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2244__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2795__A3 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2547__A3 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1989_ _0941_ _0955_ _1007_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__1755__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2180__A1 _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2483__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1887__B _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1746__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1797__B _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1912_ _0731_ _0952_ _0948_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2892_ _0584_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1985__A1 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1843_ _0919_ _0920_ _0835_ _0637_ _0639_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_30_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2529__A3 _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1774_ _0766_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2421__B _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2326_ _1352_ _1404_ _1286_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2257_ _1316_ _1320_ _1326_ _1328_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_65_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2188_ _1379_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1500__B _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1976__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1728__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1900__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2456__A2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1967__B2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1967__A1 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1719__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2392__A1 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1490_ _0276_ _0297_ _0330_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_3_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2111_ _1181_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2042_ _0276_ _0710_ _0880_ _1002_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1958__A1 _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2875_ _0612_ _0572_ _0573_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1826_ _0824_ _0889_ _0890_ _0903_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__1546__I _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1757_ _0657_ _0669_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1688_ _0766_ _0658_ _0652_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2919__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2135__A1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2309_ _1312_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2326__B _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1949__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2126__A1 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2660_ _0299_ _0348_ _0030_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1794__C _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1611_ _0687_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_5_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2591_ _0272_ _1404_ _0074_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2365__A1 _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1542_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1473_ _0080_ _0113_ _0145_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_4_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2117__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I EN vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2668__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2025_ _1096_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2927_ _0019_ net52 clknet_1_0__leaf_CLK net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__1985__B _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2858_ _0552_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_2789_ _0487_ _0447_ _0488_ _0445_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1809_ _0609_ _0884_ _0886_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_49_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1619__C2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1619__B1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2595__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2712_ _0295_ _0337_ _0404_ _0405_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2586__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2643_ _0326_ _0327_ _0331_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_2574_ _0256_ _0251_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_1525_ p_shaping_Q.bit_in_1 _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2889__A2 net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1561__A2 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1456_ _1335_ _1357_ _1379_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2510__B2 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2008_ _1081_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2501__A1 _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2804__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1791__A2 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1644__I _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2740__A1 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2290_ _1318_ _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2626_ _0311_ _0312_ _0222_ _0087_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2557_ _0237_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1534__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2488_ _0151_ _0157_ _0162_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_1508_ _0221_ _0341_ _0459_ _0522_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2798__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2014__A3 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1464__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2509__B _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2244__B _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1639__I _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1790_ _0865_ _0868_ _0784_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1764__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2411_ _0078_ _1310_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2342_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2273_ _1287_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2419__B _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1988_ Reg_Delay_Q.Out _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2609_ _0294_ net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1507__A2 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1459__I _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2891_ _0418_ _0503_ _0584_ _1389_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_30_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1911_ _0608_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1842_ _0692_ _0689_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_30_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2529__A4 _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1773_ _0747_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2162__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2325_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2256_ _1313_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2187_ _1252_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1673__A1 _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2663__I _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1976__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1900__A2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2208__A3 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1967__A2 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1719__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2144__A2 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2110_ _1165_ _1171_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2041_ _1055_ _1113_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1655__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2080__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2874_ Reg_Delay_Q.In _0572_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1825_ _0743_ _0889_ _0890_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XANTENNA__2907__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1756_ _0834_ _0816_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_7_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1687_ _0644_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2135__A2 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2308_ _1385_ net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2239_ _1279_ _1309_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2071__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1737__I _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2126__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2601__A3 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2062__A1 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1647__I _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1610_ _0265_ _0689_ _0653_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2590_ _0272_ _0273_ _1308_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2365__A2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1541_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1472_ _0135_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_5_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2117__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1876__A1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1628__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2024_ _0783_ _1060_ _1098_ _0661_ _1035_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2053__B2 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2926_ _0018_ net51 clknet_1_0__leaf_CLK net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2857_ _0542_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1808_ _0765_ _0790_ _0801_ _0737_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2788_ _0448_ _0446_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1739_ _0773_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1506__B _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2388__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1467__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2347__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1858__A1 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2711_ _0317_ _0324_ _0401_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2586__A2 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1794__B1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2642_ _0281_ _0329_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2573_ _1388_ _0244_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1524_ _0586_ _0599_ _0607_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1455_ _1368_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1849__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2510__A2 _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout53_I net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2007_ _0963_ _0970_ _1029_ _0771_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_63_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2909_ _0592_ _0572_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2501__A2 _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2514__C _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2568__A2 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1925__I _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_0_CLK CLK clknet_0_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__2740__A2 _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1700__B1 _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2008__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2625_ _1380_ _1436_ _0099_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2556_ _0235_ _0236_ _0570_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2487_ _0052_ _0158_ _0161_ _1374_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1507_ _0200_ _0513_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2495__A1 _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1570__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2666__I _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2798__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1758__B1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1745__I _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2722__A2 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2486__A1 _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1480__I _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2238__B2 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2238__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2017__S _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2410_ _0601_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2341_ _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2272_ _1285_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2477__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2435__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1987_ _0765_ _1057_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2401__A1 _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1755__A3 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1565__I _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2608_ _0286_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2539_ _1270_ _1406_ _0217_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_28_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1691__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1475__I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2459__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2631__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2890_ net2 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1910_ _0873_ _0975_ _0986_ _0803_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_1841_ _0630_ _0491_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_8_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1772_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2324_ _1324_ _1263_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2255_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2186_ _1324_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1673__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2622__A1 _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1736__I0 _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2803__B _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2392__A3 _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_12_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2040_ _0818_ _1059_ _0917_ _1055_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_47_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1655__A2 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2873_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1824_ _0891_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1755_ _0702_ _1432_ _0395_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_1686_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_38_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2307_ _1310_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2238_ _1282_ _1283_ _1306_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__2674__I _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2169_ _1227_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2843__A1 _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1646__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1582__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1540_ _0091_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2365__A3 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1471_ _0124_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1876__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2023_ _1056_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2825__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2925_ _0017_ net51 clknet_1_0__leaf_CLK net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2856_ _0537_ _0553_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1800__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1807_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2787_ _0399_ _0408_ _0398_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1738_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1669_ _0470_ _0747_ _0695_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1573__I _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1506__C _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1748__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2353__B _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1555__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1858__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2263__B _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2710_ _0317_ _0324_ _0401_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2641_ _1273_ _0050_ _0154_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2572_ _0117_ _0173_ _0180_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1523_ _0599_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1454_ net32 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1849__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2006_ _1002_ _1024_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_fanout46_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2274__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1568__I _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2908_ _0022_ _0596_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1785__A1 _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2839_ _0516_ _0539_ _0540_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2348__B _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__A1 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1700__B2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1700__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2008__A2 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1767__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2624_ _0151_ _0157_ _0162_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_2555_ _0117_ _0172_ _0179_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__2192__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1506_ _0481_ _0502_ _0438_ _0384_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_2486_ _0052_ _0159_ _0160_ _0108_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_46_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1758__B2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2722__A3 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1930__A1 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2486__A2 _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2238__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1997__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2541__B _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2340_ _1369_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__1921__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2271_ _1334_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1986_ _0673_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2607_ _0288_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2165__A1 _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2538_ _1299_ _1303_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1581__I _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2469_ _0083_ _0142_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2626__B _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2640__A2 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2156__A1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2459__A2 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1840_ _0864_ _0917_ _0836_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_8_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2395__A1 _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1771_ _0836_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1666__I p_shaping_Q.bit_in_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2497__I _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2323_ _1334_ _1401_ _1348_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2254_ _1293_ _1258_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2185_ _1250_ _1280_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1658__B1 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2622__A2 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2181__B _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1969_ _0988_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2689__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1486__I _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2301__B2 _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2852__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2872_ _0439_ _0415_ _0412_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1823_ _0892_ _0895_ _0897_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_30_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1754_ _0627_ _0633_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_1685_ _0724_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2306_ _1315_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2237_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2168_ _1211_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2099_ _1165_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1582__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1470_ net38 _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2022_ _0757_ _0952_ _0709_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2825__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2589__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2924_ _0016_ net51 clknet_1_0__leaf_CLK net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2855_ _0557_ net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1806_ _0167_ _0533_ _0861_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_2786_ _0453_ _0485_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1737_ _0703_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2761__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1668_ _0630_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1599_ _0673_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2044__A3 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1555__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2504__A1 _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1618__I0 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2640_ _0038_ _0298_ _1408_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1794__A2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2571_ _0049_ _0236_ _0252_ _0122_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__1674__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2743__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1522_ _0603_ _0604_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1453_ _1346_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1623__B _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2005_ _1075_ _1077_ _1079_ _0725_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2454__B _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2907_ _0828_ p_shaping_Q.counter\[0\] _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1785__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2838_ _0493_ _0514_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2769_ _0425_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1776__A2 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1494__I _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2539__B _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1767__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2623_ _0300_ _0301_ _0306_ _0309_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_2554_ _0233_ _0234_ _1278_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_1505_ _0491_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2485_ _1362_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_55_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1579__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1758__A2 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__1694__A1 _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1997__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1921__A2 _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2270_ _1277_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1985_ _0839_ _1059_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2606_ _0289_ _0141_ _0290_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2537_ _0108_ _0055_ _0111_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2468_ _0140_ _0141_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1912__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2399_ _1370_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2156__A2 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1903__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1770_ _0812_ _0384_ _0848_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__2395__A2 _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2147__A2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1682__I _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2322_ _1399_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2253_ _1322_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1658__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2184_ _1335_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1658__B2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1631__B _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2083__A1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2622__A3 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1968_ _1035_ _1038_ _1040_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1899_ _0852_ _0732_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2138__A2 _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2074__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2091__C _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1888__A1 _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2871_ _0569_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1677__I _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1822_ _0898_ _0900_ _0794_ _0850_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1753_ _0625_ _0287_ _0631_ _0645_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_7_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1684_ _0758_ _0759_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2305_ _1358_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2540__A2 _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2236_ _1291_ _1261_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2457__B _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2843__A3 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2167_ _1234_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2098_ _1166_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2056__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1587__I _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2047__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2021_ _1063_ _1065_ Reg_Delay_Q.Out _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_35_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2791__I _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2589__A2 _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2923_ _0015_ net51 clknet_1_0__leaf_CLK net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2854_ _0553_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2785_ _0471_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_1805_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1736_ _0808_ _0654_ _0811_ _0813_ _0760_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_1667_ _0730_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1598_ _0675_ _0297_ _0676_ _0677_ _0670_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2513__A2 _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1870__I _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2219_ _1268_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2504__A2 _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2876__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1618__I1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2570_ _0240_ _0245_ _0251_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2743__A2 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1521_ p_shaping_I.ctl_1 net57 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1452_ net33 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2004_ _1075_ _1078_ _1077_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2906_ _1158_ _0595_ _0594_ _0712_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2837_ _0493_ _0514_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2768_ _0360_ _0245_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1719_ _0756_ _0796_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2699_ _0388_ _1425_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2696__I _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2498__A1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1473__A2 _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2422__A1 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1776__A3 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2380__B _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1700__A3 _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1685__I _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2922__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2622_ _0302_ _1407_ _0307_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_2553_ _0194_ _0056_ _1408_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_1504_ _0135_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2484_ _0053_ _1301_ _1303_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2465__B _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2404__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1694__A2 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2891__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1719__B _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_0_CLK_I CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2938__RN net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2882__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2634__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1984_ _0668_ _0749_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2605_ _0085_ _0138_ _0139_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2929__RN net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2536_ _1410_ _1407_ _0105_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2467_ _0138_ _0139_ _0085_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2398_ _1294_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2625__A1 _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2864__A1 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2321_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2252_ _1298_ _1323_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2183_ _0826_ _1249_ net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1658__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2607__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1967_ _0694_ _0877_ _1041_ _1042_ _0210_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_1898_ _0884_ _0933_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2519_ _1411_ _0193_ _0196_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XANTENNA__1822__B _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2074__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2129__A3 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1888__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2301__A3 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2870_ net1 Reg_Delay_Q.In _0599_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1821_ _0674_ _0899_ _0113_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__A1 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1752_ _0720_ _0769_ _0745_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1683_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1879__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2304_ _1359_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2828__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2235_ _1286_ _1288_ _1295_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2166_ _1213_ _1233_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2457__C _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1500__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2097_ _1167_ _1168_ _1169_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2056__A2 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1803__A2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2531__A3 _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1778__I _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2047__A2 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2020_ _0722_ _1093_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_47_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2922_ _0014_ net54 clknet_1_1__leaf_CLK net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XANTENNA__2589__A3 _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1797__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2853_ _0538_ _0542_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1549__A1 _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1804_ _0707_ _0879_ _0881_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_2784_ _0478_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1735_ _0766_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1666_ p_shaping_Q.bit_in_2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1597_ _0470_ _0145_ _0373_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2218_ _1379_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2149_ _1201_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1788__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1960__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1779__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__2743__A3 _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1951__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1520_ net48 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1451_ _1324_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2900__B1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2003_ _0622_ _0761_ _0898_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2905_ _0762_ _0594_ _0595_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2836_ _0537_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__2719__B1 _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2767_ _0426_ _0230_ _0429_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_2_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1718_ _0438_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2698_ _0389_ _0390_ _0213_ _0353_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_1649_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_58_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2498__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2422__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1740__B _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2661__A2 _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2413__A2 _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2621_ _0241_ _1336_ _0213_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2552_ _0226_ _0229_ _0231_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1503_ _0470_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1915__B _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1924__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1924__B2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2483_ _1322_ _1442_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_fanout44_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2481__B _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2168__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2819_ _0323_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1915__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2891__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2159__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1906__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2882__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2634__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1983_ _0650_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2604_ _0147_ _0201_ _0202_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2570__A1 _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2535_ _0212_ _0213_ _1420_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2466_ _0085_ _0138_ _0139_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2397_ _1417_ _1418_ _1439_ _0062_ _0063_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_56_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2625__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2389__A1 _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2561__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2552__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2320_ _1263_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2251_ _1368_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2182_ _0822_ _0825_ _0742_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2296__B _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2607__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1966_ _0481_ _0812_ _0696_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1897_ _0745_ _0972_ _0973_ _0721_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2543__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2518_ _0194_ _0065_ _0195_ _0038_ _1307_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2449_ _0118_ _0120_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2935__CLK _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2846__A2 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1820_ _0626_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1751_ _0743_ _0806_ _0821_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_7_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1576__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2773__A1 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1682_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1907__C _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2303_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1923__B _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2234_ _1297_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2165_ _1213_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1500__A2 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2096_ _1064_ _0544_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1803__A3 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2920__D _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1949_ _0645_ _0816_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2764__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2522__A4 _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2921_ _0013_ net55 clknet_1_1__leaf_CLK net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1797__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2852_ _0534_ _0536_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1803_ _0850_ _0849_ _0855_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_2783_ _0479_ _0480_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2746__A1 _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1734_ _0809_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1665_ _0721_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1596_ _0632_ _0308_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1653__B _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1721__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2217_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2148_ _1214_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2079_ _0988_ _1048_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1788__A2 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2503__I _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2268__A3 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2394__B _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1779__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2743__A4 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1450_ net31 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1951__A2 _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2900__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2900__B2 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2002_ _0761_ _0796_ _0713_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__2664__B1 _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2904_ _0870_ _0572_ _0587_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2835_ _0534_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_31_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2719__B2 _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2719__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2766_ _1320_ _0042_ _0328_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1717_ _0319_ _0649_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_2697_ _0298_ _1328_ _0217_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1648_ _0727_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1579_ net44 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1630__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1933__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2389__B _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2489__A3 _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1697__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1740__C _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2110__A2 _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2571__C _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1621__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2620_ _0302_ _0305_ _1412_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__1982__I _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2551_ _1433_ _0115_ _0230_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_1502_ _0069_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2482_ _0152_ _0155_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1688__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2818_ _0519_ net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2749_ _0443_ _0444_ _0411_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1679__A1 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2228__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1851__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1906__A2 _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2095__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2095__B2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1982_ _0708_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2603_ _1415_ _0082_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2534_ _1337_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2465_ _1387_ _0125_ _0126_ _0137_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__2570__A2 _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2396_ _1359_ _1438_ _0048_ _0061_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2757__B _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2086__A1 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2625__A3 _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1833__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2923__D _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2389__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2010__A1 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2561__A2 _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2077__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1746__B _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2250_ _1321_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2577__B _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2181_ _1242_ _1245_ _1247_ _1248_ net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1815__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1965_ _0854_ _0750_ _0693_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1896_ _0964_ _0969_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2331__I _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2543__A2 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2517_ _1317_ _0065_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_2448_ _0592_ _0119_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__2918__D _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2379_ _1253_ _1267_ _0043_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2059__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1806__A1 _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1566__B _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2298__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1750_ _0828_ _0770_ _0780_ _0805_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_7_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1681_ _0657_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2773__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2302_ _1367_ _1369_ _1378_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2233_ _1299_ _1301_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2164_ _1228_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2095_ _0981_ _0945_ _1003_ _1054_ _1145_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_61_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2461__A1 _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2770__B _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1948_ _0113_ _0834_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1879_ _0940_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2764__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2516__A2 _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2204__A1 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2691__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2443__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2920_ _0012_ net54 clknet_1_1__leaf_CLK net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffrnq_1
X_2851_ _0546_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2590__B _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2925__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1802_ _0759_ _0878_ _0880_ _0210_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_2782_ _0078_ _0477_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1733_ _0747_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_1664_ _0723_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1595_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2216_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2765__B _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2147_ _1215_ _1199_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__2682__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2078_ _1145_ _0638_ _1042_ _1146_ _1150_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_34_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2931__D p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2737__A2 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1960__A3 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2425__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1779__A3 _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2728__A2 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2900__A2 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2585__B _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2001_ _0481_ _0036_ _0854_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2664__B2 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2664__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2416__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output8_I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2903_ _0788_ _0593_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2834_ _0500_ _0507_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2719__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2765_ _0267_ _0461_ _0462_ _1386_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_2696_ _0272_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1716_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1647_ _0702_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_1578_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2495__B _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2926__D _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2407__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__1839__B _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1630__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2894__A1 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2646__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2550_ _1285_ _0066_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2481_ _0153_ _0154_ _1369_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1501_ _0200_ _0449_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1688__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2885__A1 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2637__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1503__I _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1860__A2 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2817_ _0515_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2748_ _0411_ _0443_ _0444_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2679_ _0368_ _0369_ _0281_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1679__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2891__A4 _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2619__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2095__A2 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1981_ _1054_ _0757_ _1055_ _0867_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2602_ _0146_ _0138_ _0203_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2533_ _1347_ _1404_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2464_ _1314_ _0125_ _0126_ _0137_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_2395_ _0048_ _0061_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_3_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2329__I _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1530__A1 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1597__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2010__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2849__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1852__B _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2667__C _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1824__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2001__A2 _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1760__A1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2180_ _0022_ _1084_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1988__I Reg_Delay_Q.Out vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1815__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1964_ _0640_ _0849_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2612__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1895_ _0717_ _0779_ _0842_ _0922_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2516_ _1322_ _0074_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1751__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2447_ p_shaping_I.bit_in _0605_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__2487__C _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2378_ _1339_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_44_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2059__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1847__B _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1582__B _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2298__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1680_ _0502_ _0708_ _0384_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__1981__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2301_ _1371_ _1373_ _1374_ _1376_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_2232_ _1265_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2163_ _0874_ _1230_ _1231_ _0863_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2094_ _1063_ _1065_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2461__A2 _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1947_ _0851_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1878_ _0942_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_0_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2204__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1963__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1715__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2140__A1 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2850_ _0529_ _0531_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_1801_ _0625_ _0659_ _0156_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2781_ _1345_ _0300_ _0273_ _0435_ _0426_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__2746__A3 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1732_ _0809_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1663_ _0718_ _0741_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1594_ _0624_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2215_ _1346_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2765__C _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2146_ _1190_ _1195_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2077_ _0785_ _1147_ _1149_ _0782_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_41_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2072__I _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2005__C _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1844__C _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2021__B Reg_Delay_Q.Out vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2247__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2113__A1 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2000_ _0330_ _0833_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2664__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__B1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2902_ _0584_ _0571_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_2833_ _0508_ _0512_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2764_ _0238_ _0421_ _0422_ _0224_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1715_ _0680_ _0653_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2695_ _0353_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1646_ _0725_ _0672_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1577_ net45 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1680__B _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2655__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2129_ _1190_ _1195_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2407__A2 _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1839__C _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1918__A1 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2591__A1 _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2915__CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1765__B _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1909__A1 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2582__A1 _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1500_ _0362_ _0384_ _0416_ _0438_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2480_ _0037_ _1406_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2334__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1688__A3 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2637__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2816_ _0516_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2747_ _1315_ _0434_ _0442_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2573__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2678_ _0028_ _0195_ _0131_ _0367_ _0366_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_1629_ _0632_ _0648_ _0102_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2938__CLK net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2937__D p_shaping_Q.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2260__I _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2619__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1980_ _0753_ _0920_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2601_ _0208_ _0271_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_9_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2555__A1 _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2532_ _0163_ _0209_ _1423_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__2307__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2463_ _0128_ _0136_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2394_ _0049_ _1414_ _0059_ _0060_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout42_I _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1833__A3 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2794__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2546__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2849__A2 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1521__A2 net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2255__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2537__A1 _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1760__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1963_ _0853_ _0816_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1894_ _0772_ _0963_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2515_ _0190_ _0191_ _0192_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2446_ _0117_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2377_ _0041_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2519__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1981__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2300_ _1281_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2231_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_31_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2162_ _1048_ _1230_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_2093_ _1064_ _0544_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1946_ _0808_ _0750_ _0920_ _0690_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1877_ _0858_ _0951_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2429_ _1307_ _0089_ _0093_ _0098_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_28_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1715__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2140__A2 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2443__A3 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1800_ _0868_ _0876_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2780_ _0332_ _0333_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1731_ _0623_ _0395_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_11_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1662_ _0664_ _0739_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2903__A1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1593_ _0670_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2214_ _1262_ _1389_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2145_ _1190_ _1195_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2076_ _0953_ _0848_ _1148_ _0681_ _0784_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2554__S _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1642__A1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1929_ _1002_ _1004_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__1945__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2302__B _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2673__A3 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1607__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2113__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__A1 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2416__A3 _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1624__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2901_ _1024_ _0788_ _0590_ _0576_ _1054_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_16_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2173__I _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2832_ _0530_ _0532_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2763_ _0238_ _0458_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_1714_ _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2694_ _0332_ _0333_ _0601_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1645_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1517__I p_shaping_I.bit_in vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1576_ _0650_ _0653_ _0654_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2128_ _0612_ _1197_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2059_ _0709_ _0712_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1918__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2040__A1 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2591__A2 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2258__I _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1909__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2270__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2815_ _0486_ _0489_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_2746_ _0144_ _0434_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_11_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2022__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2573__A2 _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2677_ _0366_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1628_ _0702_ _1432_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1781__B1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1691__B _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1559_ net45 net44 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2089__A1 _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2564__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2697__B _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2716__I _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2600_ _0283_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_2531_ _1381_ _1437_ _0099_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__2555__A2 _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2462_ _0130_ _0132_ _0134_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_2393_ _1412_ _1283_ _0045_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2400__B _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1818__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2729_ _0267_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_59_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1809__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2234__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2785__A2 _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2271__I _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2537__A2 _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__A1 _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2446__I _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2225__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2928__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1962_ _1036_ _1037_ _0850_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1893_ _0964_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_2514_ _0043_ _0129_ _1441_ _1375_ _1377_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1751__A3 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1525__I p_shaping_Q.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2445_ _0104_ _0107_ _0112_ _1420_ _0116_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_56_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2376_ _1351_ _1327_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2356__I _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2767__A2 _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2040__B _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2931__RN net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2266__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2455__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2207__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2758__A2 _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2230_ _1258_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_2161_ _0701_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2694__A1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2092_ _1154_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1945_ _1019_ _1009_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1876_ _0952_ _0638_ _0795_ _0953_ _0221_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_2428_ _0094_ _0052_ _0096_ _0097_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__2685__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2359_ _1398_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2912__A2 p_shaping_I.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2676__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__A1 _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1730_ _0080_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2600__A1 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1661_ _0740_ net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1592_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2213_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2144_ _1212_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2075_ _0948_ _0750_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__1959__B _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1928_ _0791_ _0684_ _0877_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1859_ _0884_ _0887_ _0933_ _0863_ _0609_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_30_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2658__A1 _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2544__I _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2897__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2649__A1 _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1872__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2900_ _0834_ _0817_ _0590_ _0576_ _0943_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_43_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1624__A2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2831_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2762_ _0586_ _0458_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2403__B _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1713_ _0362_ _0036_ _0416_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2693_ _0323_ _0380_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_6_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1644_ _0659_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2888__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1575_ _0621_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2127_ _1096_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2058_ _0723_ _1127_ _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__2364__I _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1918__A3 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2591__A3 _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1551__A1 _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1854__A2 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__A2 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1909__A3 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2582__A3 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1790__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1845__A2 _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2184__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2270__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2814_ _0452_ _0443_ _0485_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2745_ _0387_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2022__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2676_ _0248_ _1329_ _0109_ _0094_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_1627_ _0658_ _0189_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__1781__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1558_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1533__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1489_ _0319_ _0145_ _0113_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2089__A2 _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2043__B _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1524__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2530_ _0207_ _0201_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2555__A3 _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2888__B _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1763__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2461_ _0111_ _0133_ _0031_ _1420_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2400__C _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2392_ _0033_ _0050_ _0056_ _0057_ _1421_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_3_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2798__B _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2728_ _0237_ _0421_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__1754__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2659_ _0104_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2038__B _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1690__B1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2537__A3 _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2501__B _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1961_ _0814_ _0817_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1892_ _0966_ _0968_ _0670_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2513_ _1336_ _0131_ _1262_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2444_ _1374_ _0114_ _0115_ _1400_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_2375_ _0039_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2161__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1541__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1697__B _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2372__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1716__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2207__A2 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2758__A3 _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__A1 _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2885__C _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2143__B2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2160_ _1145_ _1025_ _1158_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2091_ _1155_ _1161_ _1163_ _0744_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_1944_ _0971_ _0974_ _0987_ _0996_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_9_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1875_ _0622_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__1709__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2382__A1 _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2427_ _1268_ _0054_ _1360_ _1254_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2358_ _1419_ _1438_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__2685__A2 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2289_ _1340_ _1265_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1948__A1 _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1446__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1890__B _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2918__CLK clknet_1_1__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2676__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2277__I _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2428__A2 _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1660_ _0664_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_1591_ _0069_ _0308_ _0102_ _0648_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2212_ net47 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2143_ _1064_ _0522_ _1196_ _1096_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_38_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2074_ _0757_ _1058_ _0865_ _0953_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_46_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1927_ _0953_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1858_ _0874_ _0873_ _0934_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__2355__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1789_ _0809_ _0696_ _0852_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__B1 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2560__I _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2594__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2346__A1 _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1904__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A2 _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2282__B1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1624__A3 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2821__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2830_ _0078_ _0476_ _0509_ _0387_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2761_ _0454_ _0456_ _0457_ _0388_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__2470__I _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2585__A1 _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2692_ _0381_ _0382_ _0383_ _0266_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1712_ _0694_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_1643_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1574_ _0362_ _0625_ _0416_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout58_I net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2126_ _1158_ _0341_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__1863__A3 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2057_ _0719_ _1128_ _1130_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2812__A2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2328__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__1724__I p_shaping_Q.bit_in_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1551__A2 _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1606__A3 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2567__A1 _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2319__A1 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1845__A3 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2813_ _0493_ _0514_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_31_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2744_ _0592_ _0437_ _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2675_ _0365_ _1394_ _1352_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1626_ _0701_ _0704_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1557_ _1443_ _0491_ _0254_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__2730__A1 _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1488_ _0308_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2109_ _1154_ _1164_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2375__I _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2797__A1 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2013__A3 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1524__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1454__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2721__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2460_ _1286_ _0092_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__2712__A1 _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2391_ _0034_ _1305_ _1355_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_3_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2195__I _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2079__I0 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1967__C _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1539__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2727_ _0182_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1754__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2658_ _0163_ _0209_ _0346_ _0310_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_59_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1609_ _0232_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_2589_ _1365_ _0094_ _0039_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_59_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__A3 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2038__C _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1449__I _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2170__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2473__A3 _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_1960_ _0675_ _0814_ _0713_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1891_ _0786_ _0844_ _0900_ _0967_ _0438_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__1984__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2512_ _1332_ _1352_ _0160_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2443_ _1280_ _1285_ _1325_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_2374_ _1298_ _1361_ _1323_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_24_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1672__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2653__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1975__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1966__A2 _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2512__B _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2391__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2090_ _1155_ _1162_ _1129_ _1161_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_46_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1943_ _0962_ _0997_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1874_ _0653_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2906__A1 _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1709__A2 _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2141__C _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2906__B2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2426_ _1277_ _1313_ _0095_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_2357_ _1424_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__1552__I _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2288_ _1290_ _1327_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1893__A1 _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__1948__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2051__C _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1462__I _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2676__A3 _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1636__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1590_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2116__A2 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2211_ _1259_ _1276_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2142_ _1208_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_2073_ _0759_ _0795_ _0778_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1627__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1926_ _0683_ _0877_ _0793_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_1857_ _0609_ _0884_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1788_ _0852_ _0865_ _0796_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_1_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2409_ _1282_ _0068_ _0071_ _0076_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__1866__A1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2291__B2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2043__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2346__A2 _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2649__A3 _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1857__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2282__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1624__A4 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2760_ _1274_ _1442_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2585__A2 _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2691_ _0320_ _0376_ _0378_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_1711_ _0785_ _0787_ _0789_ _0732_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_1642_ _0721_ p_shaping_Q.counter\[0\] _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1573_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2198__I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__1848__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2125_ _0459_ _0522_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2056_ _1129_ _1123_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2025__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1909_ _0885_ _0980_ _0985_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_2889_ _0574_ net42 _0581_ _0474_ _0583_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2328__A2 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2610__B _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2500__A2 _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2264__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput4 net4 I[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1650__I _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2812_ _0508_ _0512_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__2558__A2 _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2743_ _0439_ _0241_ _0040_ _0412_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_2674_ _0054_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1625_ _0232_ _0624_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_1556_ _0622_ _0629_ _0631_ _0633_ _0635_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2730__A2 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1487_ net46 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2494__A1 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2656__I _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1560__I _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2108_ _1180_ net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2039_ _0681_ _0677_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2797__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2549__A2 _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1735__I _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2566__I _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1470__I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2515__B _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1645__I _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2390_ _0052_ _0055_ _1354_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2476__A1 _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2425__B _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2400__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2726_ _0412_ _0413_ _0414_ _0104_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_2657_ _0214_ _0215_ _0220_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2160__B _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1608_ _0395_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__2703__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2588_ _0108_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1539_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_47_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1809__A4 _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2219__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1690__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1465__I _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2458__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1890_ _0674_ _0899_ _0755_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_2511_ _0148_ _0165_ _0183_ _0186_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_2442_ _1268_ _0054_ _1331_ _1292_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__2697__A1 _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2373_ _0037_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2464__A4 _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1672__A2 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2870__S _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2621__A1 _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2709_ _0400_ _0401_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__2688__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2049__C _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2754__I _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_1942_ _1018_ net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1873_ _0851_ _0946_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2425_ _1269_ _1255_ _1341_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_2356_ _1436_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2287_ _1266_ _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__1893__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2676__A4 _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1636__A2 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2523__B _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2061__A2 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_2210_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2141_ _1155_ _1209_ _1210_ _0666_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_38_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2072_ _0753_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2824__A1 _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1627__A2 _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1925_ _0221_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1856_ _0862_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1787_ _0853_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__2659__I _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1563__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2408_ _1366_ _0073_ _0075_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__2658__A4 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2339_ _1311_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1866__A2 _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2291__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2806__A1 _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2282__A2 _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2690_ _1423_ _0358_ _0347_ _0148_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_1710_ _0668_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_1641_ p_shaping_Q.counter\[1\] _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1572_ _0651_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_2124_ _1155_ _1193_ _1194_ _0827_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__1848__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_2055_ _1082_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2025__A2 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2888_ _0439_ _0580_ _0503_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1908_ _0754_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_1839_ _0080_ _0899_ _0838_ _0373_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2328__A3 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2264__A2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2073__B _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput5 net5 I[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput40 net40 addQ[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2248__B _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_1_0__f_CLK clknet_0_CLK clknet_1_0__leaf_CLK vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2811_ _0603_ _0510_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2742_ _0389_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2673_ _0360_ _0361_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_1624_ _0620_ _0658_ _0669_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_1555_ _0351_ _0627_ _0634_ _0254_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__2191__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_1486_ _0287_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__2494__A2 _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2107_ _1173_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_2038_ _0731_ _1058_ _1076_ _0791_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1920__A1 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1661__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__1987__A1 _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2400__A2 _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2441__B _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2725_ _0155_ _0417_ _0419_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_2656_ _1423_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1607_ _0640_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_2587_ _1314_ _0260_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_1538_ _0200_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_1469_ _0102_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2219__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2351__B _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1902__A1 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2458__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__1969__A1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2510_ _0148_ _0165_ _0183_ _0186_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_2441_ _0108_ _0055_ _0111_ _0106_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__2697__A2 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2372_ _1284_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__1605__B _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__2449__A2 _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2708_ _0400_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__2385__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2639_ _0240_ _1342_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1476__I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2376__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2128__A1 _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1654__A3 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1941_ _1011_ _1017_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_1872_ _0330_ _0929_ _0947_ _0948_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__2367__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2119__A1 _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2424_ _1429_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_2355_ _1344_ _1428_ _1434_ _1435_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_29_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2286_ _1340_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_37_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2358__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2855__I _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__2833__A2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__2597__A1 _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2521__A1 _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2140_ _1129_ _1209_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2071_ _0824_ _1127_ _1137_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_46_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1924_ _0981_ _0965_ _1000_ _0753_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_1855_ _0724_ _0926_ _0928_ _0778_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_1786_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2760__A1 _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_2407_ _1390_ _0074_ _1321_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__2512__A1 _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2338_ p_shaping_I.counter\[0\] _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__1866__A3 _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2269_ _1339_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2579__A1 _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__2931__CLK net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2518__C _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__1490__A1 _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2282__A3 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_1640_ _0706_ _0715_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_1571_ _0058_ net46 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__1664__I _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2123_ _1129_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2054_ _1118_ _1119_ _1125_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__2444__B _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2163__C _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_2887_ _0582_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_1907_ _0786_ _0982_ _0983_ _0784_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_1838_ _0871_ _0915_ _0705_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_1769_ _0689_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__2733__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__1749__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__2354__B _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput6 net6 I[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__2724__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput30 net30 addI[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 addQ[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2810_ _0387_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_2741_ _0435_ _1350_ _0436_ _0348_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_2672_ _0163_ _0209_ _0346_ _0310_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_1623_ _0702_ _0623_ _0124_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_1554_ _1432_ _0135_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__2191__A2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_1485_ _0091_ _0135_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

