magic
tech gf180mcuC
magscale 1 10
timestamp 1670198993
<< metal1 >>
rect 36978 56590 36990 56642
rect 37042 56639 37054 56642
rect 37874 56639 37886 56642
rect 37042 56593 37886 56639
rect 37042 56590 37054 56593
rect 37874 56590 37886 56593
rect 37938 56590 37950 56642
rect 1344 56474 58576 56508
rect 1344 56422 19838 56474
rect 19890 56422 19942 56474
rect 19994 56422 20046 56474
rect 20098 56422 50558 56474
rect 50610 56422 50662 56474
rect 50714 56422 50766 56474
rect 50818 56422 58576 56474
rect 1344 56388 58576 56422
rect 4734 56306 4786 56318
rect 4734 56242 4786 56254
rect 54238 56194 54290 56206
rect 3042 56142 3054 56194
rect 3106 56142 3118 56194
rect 19506 56142 19518 56194
rect 19570 56142 19582 56194
rect 25890 56142 25902 56194
rect 25954 56142 25966 56194
rect 57810 56142 57822 56194
rect 57874 56142 57886 56194
rect 54238 56130 54290 56142
rect 21422 56082 21474 56094
rect 40910 56082 40962 56094
rect 4162 56030 4174 56082
rect 4226 56030 4238 56082
rect 8866 56030 8878 56082
rect 8930 56030 8942 56082
rect 14354 56030 14366 56082
rect 14418 56030 14430 56082
rect 20626 56030 20638 56082
rect 20690 56030 20702 56082
rect 27010 56030 27022 56082
rect 27074 56030 27086 56082
rect 37202 56030 37214 56082
rect 37266 56030 37278 56082
rect 21422 56018 21474 56030
rect 40910 56018 40962 56030
rect 41246 56082 41298 56094
rect 41246 56018 41298 56030
rect 41582 56082 41634 56094
rect 42914 56030 42926 56082
rect 42978 56030 42990 56082
rect 48850 56030 48862 56082
rect 48914 56030 48926 56082
rect 54674 56030 54686 56082
rect 54738 56030 54750 56082
rect 56690 56030 56702 56082
rect 56754 56030 56766 56082
rect 41582 56018 41634 56030
rect 13918 55970 13970 55982
rect 27582 55970 27634 55982
rect 8082 55918 8094 55970
rect 8146 55918 8158 55970
rect 15138 55918 15150 55970
rect 15202 55918 15214 55970
rect 13918 55906 13970 55918
rect 27582 55906 27634 55918
rect 36430 55970 36482 55982
rect 41134 55970 41186 55982
rect 37874 55918 37886 55970
rect 37938 55918 37950 55970
rect 36430 55906 36482 55918
rect 41134 55906 41186 55918
rect 42478 55970 42530 55982
rect 43698 55918 43710 55970
rect 43762 55918 43774 55970
rect 49522 55918 49534 55970
rect 49586 55918 49598 55970
rect 55458 55918 55470 55970
rect 55522 55918 55534 55970
rect 42478 55906 42530 55918
rect 1344 55690 58576 55724
rect 1344 55638 4478 55690
rect 4530 55638 4582 55690
rect 4634 55638 4686 55690
rect 4738 55638 35198 55690
rect 35250 55638 35302 55690
rect 35354 55638 35406 55690
rect 35458 55638 58576 55690
rect 1344 55604 58576 55638
rect 31390 55410 31442 55422
rect 1922 55358 1934 55410
rect 1986 55358 1998 55410
rect 31390 55346 31442 55358
rect 40238 55298 40290 55310
rect 54350 55298 54402 55310
rect 3042 55246 3054 55298
rect 3106 55246 3118 55298
rect 37762 55246 37774 55298
rect 37826 55246 37838 55298
rect 39778 55246 39790 55298
rect 39842 55246 39854 55298
rect 42578 55246 42590 55298
rect 42642 55246 42654 55298
rect 43698 55246 43710 55298
rect 43762 55246 43774 55298
rect 55122 55246 55134 55298
rect 55186 55246 55198 55298
rect 40238 55234 40290 55246
rect 54350 55234 54402 55246
rect 23326 55186 23378 55198
rect 23326 55122 23378 55134
rect 23662 55186 23714 55198
rect 23662 55122 23714 55134
rect 26798 55186 26850 55198
rect 26798 55122 26850 55134
rect 27134 55186 27186 55198
rect 27134 55122 27186 55134
rect 29598 55186 29650 55198
rect 29598 55122 29650 55134
rect 29934 55186 29986 55198
rect 37550 55186 37602 55198
rect 31938 55134 31950 55186
rect 32002 55134 32014 55186
rect 29934 55122 29986 55134
rect 37550 55122 37602 55134
rect 39342 55186 39394 55198
rect 44158 55186 44210 55198
rect 42242 55134 42254 55186
rect 42306 55134 42318 55186
rect 39342 55122 39394 55134
rect 44158 55122 44210 55134
rect 46622 55186 46674 55198
rect 46622 55122 46674 55134
rect 46958 55186 47010 55198
rect 56018 55134 56030 55186
rect 56082 55134 56094 55186
rect 46958 55122 47010 55134
rect 3502 55074 3554 55086
rect 3502 55010 3554 55022
rect 22878 55074 22930 55086
rect 22878 55010 22930 55022
rect 34414 55074 34466 55086
rect 34414 55010 34466 55022
rect 56590 55074 56642 55086
rect 56590 55010 56642 55022
rect 1344 54906 58576 54940
rect 1344 54854 19838 54906
rect 19890 54854 19942 54906
rect 19994 54854 20046 54906
rect 20098 54854 50558 54906
rect 50610 54854 50662 54906
rect 50714 54854 50766 54906
rect 50818 54854 58576 54906
rect 1344 54820 58576 54854
rect 40574 54738 40626 54750
rect 39666 54686 39678 54738
rect 39730 54686 39742 54738
rect 40574 54674 40626 54686
rect 37550 54626 37602 54638
rect 37550 54562 37602 54574
rect 42142 54626 42194 54638
rect 42142 54562 42194 54574
rect 42478 54514 42530 54526
rect 38210 54462 38222 54514
rect 38274 54462 38286 54514
rect 40786 54462 40798 54514
rect 40850 54462 40862 54514
rect 42478 54450 42530 54462
rect 42702 54514 42754 54526
rect 43710 54514 43762 54526
rect 43250 54462 43262 54514
rect 43314 54462 43326 54514
rect 42702 54450 42754 54462
rect 43710 54450 43762 54462
rect 43822 54514 43874 54526
rect 43822 54450 43874 54462
rect 43934 54514 43986 54526
rect 43934 54450 43986 54462
rect 39118 54402 39170 54414
rect 38434 54350 38446 54402
rect 38498 54350 38510 54402
rect 39118 54338 39170 54350
rect 39342 54402 39394 54414
rect 39342 54338 39394 54350
rect 40462 54402 40514 54414
rect 40462 54338 40514 54350
rect 42254 54402 42306 54414
rect 42254 54338 42306 54350
rect 1344 54122 58576 54156
rect 1344 54070 4478 54122
rect 4530 54070 4582 54122
rect 4634 54070 4686 54122
rect 4738 54070 35198 54122
rect 35250 54070 35302 54122
rect 35354 54070 35406 54122
rect 35458 54070 58576 54122
rect 1344 54036 58576 54070
rect 42814 53842 42866 53854
rect 40450 53790 40462 53842
rect 40514 53790 40526 53842
rect 42814 53778 42866 53790
rect 39006 53730 39058 53742
rect 39006 53666 39058 53678
rect 39342 53730 39394 53742
rect 43486 53730 43538 53742
rect 40338 53678 40350 53730
rect 40402 53678 40414 53730
rect 41570 53678 41582 53730
rect 41634 53678 41646 53730
rect 43138 53678 43150 53730
rect 43202 53678 43214 53730
rect 39342 53666 39394 53678
rect 43486 53666 43538 53678
rect 2718 53618 2770 53630
rect 2718 53554 2770 53566
rect 3166 53618 3218 53630
rect 40450 53566 40462 53618
rect 40514 53566 40526 53618
rect 41682 53566 41694 53618
rect 41746 53566 41758 53618
rect 3166 53554 3218 53566
rect 2382 53506 2434 53518
rect 2382 53442 2434 53454
rect 39118 53506 39170 53518
rect 39118 53442 39170 53454
rect 42478 53506 42530 53518
rect 42478 53442 42530 53454
rect 42926 53506 42978 53518
rect 42926 53442 42978 53454
rect 43934 53506 43986 53518
rect 43934 53442 43986 53454
rect 44382 53506 44434 53518
rect 44382 53442 44434 53454
rect 1344 53338 58576 53372
rect 1344 53286 19838 53338
rect 19890 53286 19942 53338
rect 19994 53286 20046 53338
rect 20098 53286 50558 53338
rect 50610 53286 50662 53338
rect 50714 53286 50766 53338
rect 50818 53286 58576 53338
rect 1344 53252 58576 53286
rect 35086 53170 35138 53182
rect 35086 53106 35138 53118
rect 35982 53170 36034 53182
rect 35982 53106 36034 53118
rect 40910 53170 40962 53182
rect 40910 53106 40962 53118
rect 42030 53170 42082 53182
rect 42030 53106 42082 53118
rect 42814 53170 42866 53182
rect 42814 53106 42866 53118
rect 47070 53170 47122 53182
rect 47070 53106 47122 53118
rect 38894 53058 38946 53070
rect 38894 52994 38946 53006
rect 40686 53058 40738 53070
rect 40686 52994 40738 53006
rect 42590 53058 42642 53070
rect 42590 52994 42642 53006
rect 43038 53058 43090 53070
rect 43038 52994 43090 53006
rect 43598 53058 43650 53070
rect 43598 52994 43650 53006
rect 43822 53058 43874 53070
rect 43822 52994 43874 53006
rect 33630 52946 33682 52958
rect 33630 52882 33682 52894
rect 33966 52946 34018 52958
rect 33966 52882 34018 52894
rect 34190 52946 34242 52958
rect 34190 52882 34242 52894
rect 39230 52946 39282 52958
rect 39230 52882 39282 52894
rect 40574 52946 40626 52958
rect 40574 52882 40626 52894
rect 41470 52946 41522 52958
rect 44382 52946 44434 52958
rect 41794 52894 41806 52946
rect 41858 52894 41870 52946
rect 41470 52882 41522 52894
rect 44382 52882 44434 52894
rect 46846 52946 46898 52958
rect 46846 52882 46898 52894
rect 47182 52946 47234 52958
rect 47182 52882 47234 52894
rect 47406 52946 47458 52958
rect 47406 52882 47458 52894
rect 33742 52834 33794 52846
rect 33742 52770 33794 52782
rect 34750 52834 34802 52846
rect 34750 52770 34802 52782
rect 35646 52834 35698 52846
rect 35646 52770 35698 52782
rect 36542 52834 36594 52846
rect 36542 52770 36594 52782
rect 38334 52834 38386 52846
rect 38334 52770 38386 52782
rect 39790 52834 39842 52846
rect 39790 52770 39842 52782
rect 41694 52834 41746 52846
rect 41694 52770 41746 52782
rect 42702 52834 42754 52846
rect 42702 52770 42754 52782
rect 45054 52834 45106 52846
rect 45054 52770 45106 52782
rect 46398 52834 46450 52846
rect 46398 52770 46450 52782
rect 47966 52834 48018 52846
rect 47966 52770 48018 52782
rect 43710 52722 43762 52734
rect 43710 52658 43762 52670
rect 44158 52722 44210 52734
rect 44158 52658 44210 52670
rect 1344 52554 58576 52588
rect 1344 52502 4478 52554
rect 4530 52502 4582 52554
rect 4634 52502 4686 52554
rect 4738 52502 35198 52554
rect 35250 52502 35302 52554
rect 35354 52502 35406 52554
rect 35458 52502 58576 52554
rect 1344 52468 58576 52502
rect 34862 52386 34914 52398
rect 42030 52386 42082 52398
rect 38994 52334 39006 52386
rect 39058 52334 39070 52386
rect 40786 52334 40798 52386
rect 40850 52383 40862 52386
rect 41794 52383 41806 52386
rect 40850 52337 41806 52383
rect 40850 52334 40862 52337
rect 41794 52334 41806 52337
rect 41858 52334 41870 52386
rect 34862 52322 34914 52334
rect 42030 52322 42082 52334
rect 42814 52386 42866 52398
rect 42814 52322 42866 52334
rect 43262 52386 43314 52398
rect 43262 52322 43314 52334
rect 43934 52386 43986 52398
rect 43934 52322 43986 52334
rect 45950 52386 46002 52398
rect 45950 52322 46002 52334
rect 35086 52274 35138 52286
rect 35086 52210 35138 52222
rect 36654 52274 36706 52286
rect 36654 52210 36706 52222
rect 38334 52274 38386 52286
rect 38334 52210 38386 52222
rect 40462 52274 40514 52286
rect 40462 52210 40514 52222
rect 40910 52274 40962 52286
rect 43710 52274 43762 52286
rect 42466 52222 42478 52274
rect 42530 52222 42542 52274
rect 40910 52210 40962 52222
rect 43710 52210 43762 52222
rect 44158 52274 44210 52286
rect 44158 52210 44210 52222
rect 45390 52274 45442 52286
rect 49310 52274 49362 52286
rect 47058 52222 47070 52274
rect 47122 52222 47134 52274
rect 45390 52210 45442 52222
rect 49310 52210 49362 52222
rect 32510 52162 32562 52174
rect 36430 52162 36482 52174
rect 2818 52110 2830 52162
rect 2882 52110 2894 52162
rect 33170 52110 33182 52162
rect 33234 52110 33246 52162
rect 33842 52110 33854 52162
rect 33906 52110 33918 52162
rect 32510 52098 32562 52110
rect 36430 52098 36482 52110
rect 37438 52162 37490 52174
rect 37438 52098 37490 52110
rect 39118 52162 39170 52174
rect 41358 52162 41410 52174
rect 39778 52110 39790 52162
rect 39842 52110 39854 52162
rect 39118 52098 39170 52110
rect 41358 52098 41410 52110
rect 42254 52162 42306 52174
rect 42254 52098 42306 52110
rect 47630 52162 47682 52174
rect 47630 52098 47682 52110
rect 48750 52162 48802 52174
rect 48750 52098 48802 52110
rect 35870 52050 35922 52062
rect 1922 51998 1934 52050
rect 1986 51998 1998 52050
rect 32722 51998 32734 52050
rect 32786 51998 32798 52050
rect 34514 51998 34526 52050
rect 34578 51998 34590 52050
rect 35870 51986 35922 51998
rect 36094 52050 36146 52062
rect 36094 51986 36146 51998
rect 36206 52050 36258 52062
rect 36206 51986 36258 51998
rect 42590 52050 42642 52062
rect 42590 51986 42642 51998
rect 44382 52050 44434 52062
rect 44382 51986 44434 51998
rect 46510 52050 46562 52062
rect 46510 51986 46562 51998
rect 47518 52050 47570 52062
rect 47518 51986 47570 51998
rect 47742 52050 47794 52062
rect 47742 51986 47794 51998
rect 26798 51938 26850 51950
rect 26798 51874 26850 51886
rect 32622 51938 32674 51950
rect 32622 51874 32674 51886
rect 37886 51938 37938 51950
rect 37886 51874 37938 51886
rect 46062 51938 46114 51950
rect 46062 51874 46114 51886
rect 46286 51938 46338 51950
rect 46286 51874 46338 51886
rect 48414 51938 48466 51950
rect 48414 51874 48466 51886
rect 1344 51770 58576 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 58576 51770
rect 1344 51684 58576 51718
rect 23550 51602 23602 51614
rect 23550 51538 23602 51550
rect 24670 51602 24722 51614
rect 24670 51538 24722 51550
rect 38334 51602 38386 51614
rect 38334 51538 38386 51550
rect 43150 51602 43202 51614
rect 43150 51538 43202 51550
rect 49870 51602 49922 51614
rect 49870 51538 49922 51550
rect 26238 51490 26290 51502
rect 26238 51426 26290 51438
rect 28030 51490 28082 51502
rect 28030 51426 28082 51438
rect 40350 51490 40402 51502
rect 40350 51426 40402 51438
rect 41470 51490 41522 51502
rect 41470 51426 41522 51438
rect 43822 51490 43874 51502
rect 43822 51426 43874 51438
rect 23438 51378 23490 51390
rect 23438 51314 23490 51326
rect 23662 51378 23714 51390
rect 23662 51314 23714 51326
rect 24110 51378 24162 51390
rect 24110 51314 24162 51326
rect 24558 51378 24610 51390
rect 24558 51314 24610 51326
rect 24894 51378 24946 51390
rect 33742 51378 33794 51390
rect 35310 51378 35362 51390
rect 38334 51378 38386 51390
rect 27346 51326 27358 51378
rect 27410 51326 27422 51378
rect 32386 51326 32398 51378
rect 32450 51326 32462 51378
rect 34178 51326 34190 51378
rect 34242 51326 34254 51378
rect 36082 51326 36094 51378
rect 36146 51326 36158 51378
rect 37426 51326 37438 51378
rect 37490 51326 37502 51378
rect 24894 51314 24946 51326
rect 33742 51314 33794 51326
rect 35310 51314 35362 51326
rect 38334 51314 38386 51326
rect 40126 51378 40178 51390
rect 40126 51314 40178 51326
rect 40462 51378 40514 51390
rect 40462 51314 40514 51326
rect 43262 51378 43314 51390
rect 43262 51314 43314 51326
rect 47294 51378 47346 51390
rect 49534 51378 49586 51390
rect 47954 51326 47966 51378
rect 48018 51326 48030 51378
rect 47294 51314 47346 51326
rect 49534 51314 49586 51326
rect 49758 51378 49810 51390
rect 49758 51314 49810 51326
rect 50206 51378 50258 51390
rect 50206 51314 50258 51326
rect 21870 51266 21922 51278
rect 34638 51266 34690 51278
rect 39342 51266 39394 51278
rect 27682 51214 27694 51266
rect 27746 51214 27758 51266
rect 32274 51214 32286 51266
rect 32338 51214 32350 51266
rect 37538 51214 37550 51266
rect 37602 51214 37614 51266
rect 21870 51202 21922 51214
rect 34638 51202 34690 51214
rect 39342 51202 39394 51214
rect 39678 51266 39730 51278
rect 39678 51202 39730 51214
rect 42030 51266 42082 51278
rect 42030 51202 42082 51214
rect 42702 51266 42754 51278
rect 42702 51202 42754 51214
rect 44830 51266 44882 51278
rect 44830 51202 44882 51214
rect 45166 51266 45218 51278
rect 45166 51202 45218 51214
rect 45726 51266 45778 51278
rect 45726 51202 45778 51214
rect 46174 51266 46226 51278
rect 46174 51202 46226 51214
rect 46510 51266 46562 51278
rect 46510 51202 46562 51214
rect 48750 51266 48802 51278
rect 48750 51202 48802 51214
rect 50766 51266 50818 51278
rect 50766 51202 50818 51214
rect 26126 51154 26178 51166
rect 26126 51090 26178 51102
rect 26462 51154 26514 51166
rect 38446 51154 38498 51166
rect 32722 51102 32734 51154
rect 32786 51102 32798 51154
rect 26462 51090 26514 51102
rect 38446 51090 38498 51102
rect 38670 51154 38722 51166
rect 38670 51090 38722 51102
rect 43486 51154 43538 51166
rect 43486 51090 43538 51102
rect 44046 51154 44098 51166
rect 47506 51102 47518 51154
rect 47570 51102 47582 51154
rect 44046 51090 44098 51102
rect 1344 50986 58576 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 58576 50986
rect 1344 50900 58576 50934
rect 36318 50818 36370 50830
rect 40126 50818 40178 50830
rect 49198 50818 49250 50830
rect 37426 50766 37438 50818
rect 37490 50815 37502 50818
rect 37874 50815 37886 50818
rect 37490 50769 37886 50815
rect 37490 50766 37502 50769
rect 37874 50766 37886 50769
rect 37938 50815 37950 50818
rect 38434 50815 38446 50818
rect 37938 50769 38446 50815
rect 37938 50766 37950 50769
rect 38434 50766 38446 50769
rect 38498 50766 38510 50818
rect 47394 50766 47406 50818
rect 47458 50815 47470 50818
rect 48290 50815 48302 50818
rect 47458 50769 48302 50815
rect 47458 50766 47470 50769
rect 48290 50766 48302 50769
rect 48354 50766 48366 50818
rect 36318 50754 36370 50766
rect 40126 50754 40178 50766
rect 49198 50754 49250 50766
rect 49534 50818 49586 50830
rect 49534 50754 49586 50766
rect 50318 50818 50370 50830
rect 50754 50766 50766 50818
rect 50818 50815 50830 50818
rect 51314 50815 51326 50818
rect 50818 50769 51326 50815
rect 50818 50766 50830 50769
rect 51314 50766 51326 50769
rect 51378 50766 51390 50818
rect 50318 50754 50370 50766
rect 27470 50706 27522 50718
rect 24658 50654 24670 50706
rect 24722 50654 24734 50706
rect 27470 50642 27522 50654
rect 37438 50706 37490 50718
rect 37438 50642 37490 50654
rect 38334 50706 38386 50718
rect 48302 50706 48354 50718
rect 39778 50654 39790 50706
rect 39842 50654 39854 50706
rect 42466 50654 42478 50706
rect 42530 50654 42542 50706
rect 38334 50642 38386 50654
rect 48302 50642 48354 50654
rect 50430 50706 50482 50718
rect 50430 50642 50482 50654
rect 50878 50706 50930 50718
rect 50878 50642 50930 50654
rect 51326 50706 51378 50718
rect 51326 50642 51378 50654
rect 22542 50594 22594 50606
rect 22194 50542 22206 50594
rect 22258 50542 22270 50594
rect 22542 50530 22594 50542
rect 22766 50594 22818 50606
rect 26126 50594 26178 50606
rect 36094 50594 36146 50606
rect 24098 50542 24110 50594
rect 24162 50542 24174 50594
rect 26338 50542 26350 50594
rect 26402 50542 26414 50594
rect 22766 50530 22818 50542
rect 26126 50530 26178 50542
rect 36094 50530 36146 50542
rect 36542 50594 36594 50606
rect 36542 50530 36594 50542
rect 36766 50594 36818 50606
rect 36766 50530 36818 50542
rect 37886 50594 37938 50606
rect 41022 50594 41074 50606
rect 45390 50594 45442 50606
rect 38994 50542 39006 50594
rect 39058 50542 39070 50594
rect 42690 50542 42702 50594
rect 42754 50542 42766 50594
rect 43474 50542 43486 50594
rect 43538 50542 43550 50594
rect 44706 50542 44718 50594
rect 44770 50542 44782 50594
rect 37886 50530 37938 50542
rect 41022 50530 41074 50542
rect 45390 50530 45442 50542
rect 9214 50482 9266 50494
rect 9214 50418 9266 50430
rect 25006 50482 25058 50494
rect 25006 50418 25058 50430
rect 27022 50482 27074 50494
rect 27022 50418 27074 50430
rect 34750 50482 34802 50494
rect 34750 50418 34802 50430
rect 35198 50482 35250 50494
rect 35198 50418 35250 50430
rect 39230 50482 39282 50494
rect 39230 50418 39282 50430
rect 39902 50482 39954 50494
rect 39902 50418 39954 50430
rect 42030 50482 42082 50494
rect 45726 50482 45778 50494
rect 42578 50430 42590 50482
rect 42642 50430 42654 50482
rect 43362 50430 43374 50482
rect 43426 50430 43438 50482
rect 42030 50418 42082 50430
rect 45726 50418 45778 50430
rect 49758 50482 49810 50494
rect 49758 50418 49810 50430
rect 52110 50482 52162 50494
rect 52110 50418 52162 50430
rect 8878 50370 8930 50382
rect 8878 50306 8930 50318
rect 23214 50370 23266 50382
rect 23214 50306 23266 50318
rect 31838 50370 31890 50382
rect 31838 50306 31890 50318
rect 33070 50370 33122 50382
rect 33070 50306 33122 50318
rect 33518 50370 33570 50382
rect 33518 50306 33570 50318
rect 35646 50370 35698 50382
rect 41582 50370 41634 50382
rect 40674 50318 40686 50370
rect 40738 50318 40750 50370
rect 35646 50306 35698 50318
rect 41582 50306 41634 50318
rect 45614 50370 45666 50382
rect 45614 50306 45666 50318
rect 46174 50370 46226 50382
rect 46174 50306 46226 50318
rect 46846 50370 46898 50382
rect 47854 50370 47906 50382
rect 47170 50318 47182 50370
rect 47234 50318 47246 50370
rect 46846 50306 46898 50318
rect 47854 50306 47906 50318
rect 48638 50370 48690 50382
rect 48638 50306 48690 50318
rect 1344 50202 58576 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 58576 50202
rect 1344 50116 58576 50150
rect 40910 50034 40962 50046
rect 40910 49970 40962 49982
rect 42366 50034 42418 50046
rect 47518 50034 47570 50046
rect 43586 49982 43598 50034
rect 43650 49982 43662 50034
rect 42366 49970 42418 49982
rect 47518 49970 47570 49982
rect 9774 49922 9826 49934
rect 9774 49858 9826 49870
rect 24222 49922 24274 49934
rect 24222 49858 24274 49870
rect 26798 49922 26850 49934
rect 26798 49858 26850 49870
rect 28142 49922 28194 49934
rect 31614 49922 31666 49934
rect 30034 49870 30046 49922
rect 30098 49870 30110 49922
rect 28142 49858 28194 49870
rect 31614 49858 31666 49870
rect 36094 49922 36146 49934
rect 36094 49858 36146 49870
rect 42254 49922 42306 49934
rect 42254 49858 42306 49870
rect 13246 49810 13298 49822
rect 10434 49758 10446 49810
rect 10498 49758 10510 49810
rect 13246 49746 13298 49758
rect 13470 49810 13522 49822
rect 13470 49746 13522 49758
rect 13918 49810 13970 49822
rect 21534 49810 21586 49822
rect 22430 49810 22482 49822
rect 20626 49758 20638 49810
rect 20690 49758 20702 49810
rect 22194 49758 22206 49810
rect 22258 49758 22270 49810
rect 13918 49746 13970 49758
rect 21534 49746 21586 49758
rect 22430 49746 22482 49758
rect 23662 49810 23714 49822
rect 23662 49746 23714 49758
rect 23998 49810 24050 49822
rect 23998 49746 24050 49758
rect 26574 49810 26626 49822
rect 26574 49746 26626 49758
rect 26686 49810 26738 49822
rect 26686 49746 26738 49758
rect 27694 49810 27746 49822
rect 27694 49746 27746 49758
rect 28254 49810 28306 49822
rect 36206 49810 36258 49822
rect 46846 49810 46898 49822
rect 30258 49758 30270 49810
rect 30322 49758 30334 49810
rect 31154 49758 31166 49810
rect 31218 49758 31230 49810
rect 36418 49758 36430 49810
rect 36482 49758 36494 49810
rect 28254 49746 28306 49758
rect 36206 49746 36258 49758
rect 46846 49746 46898 49758
rect 13358 49698 13410 49710
rect 9986 49646 9998 49698
rect 10050 49646 10062 49698
rect 13358 49634 13410 49646
rect 19966 49698 20018 49710
rect 27918 49698 27970 49710
rect 21186 49646 21198 49698
rect 21250 49646 21262 49698
rect 19966 49634 20018 49646
rect 27918 49634 27970 49646
rect 32062 49698 32114 49710
rect 32062 49634 32114 49646
rect 32510 49698 32562 49710
rect 32510 49634 32562 49646
rect 34190 49698 34242 49710
rect 34190 49634 34242 49646
rect 36990 49698 37042 49710
rect 36990 49634 37042 49646
rect 37438 49698 37490 49710
rect 37438 49634 37490 49646
rect 38894 49698 38946 49710
rect 38894 49634 38946 49646
rect 39342 49698 39394 49710
rect 39342 49634 39394 49646
rect 39790 49698 39842 49710
rect 39790 49634 39842 49646
rect 40462 49698 40514 49710
rect 40462 49634 40514 49646
rect 41470 49698 41522 49710
rect 41470 49634 41522 49646
rect 42926 49698 42978 49710
rect 42926 49634 42978 49646
rect 44158 49698 44210 49710
rect 44158 49634 44210 49646
rect 44606 49698 44658 49710
rect 44606 49634 44658 49646
rect 45166 49698 45218 49710
rect 45166 49634 45218 49646
rect 45502 49698 45554 49710
rect 45502 49634 45554 49646
rect 46286 49698 46338 49710
rect 46286 49634 46338 49646
rect 47406 49698 47458 49710
rect 47406 49634 47458 49646
rect 47966 49698 48018 49710
rect 47966 49634 48018 49646
rect 48638 49698 48690 49710
rect 48638 49634 48690 49646
rect 49534 49698 49586 49710
rect 49534 49634 49586 49646
rect 49982 49698 50034 49710
rect 49982 49634 50034 49646
rect 50318 49698 50370 49710
rect 50318 49634 50370 49646
rect 50766 49698 50818 49710
rect 50766 49634 50818 49646
rect 51326 49698 51378 49710
rect 51326 49634 51378 49646
rect 51998 49698 52050 49710
rect 51998 49634 52050 49646
rect 52446 49698 52498 49710
rect 52446 49634 52498 49646
rect 52894 49698 52946 49710
rect 52894 49634 52946 49646
rect 53230 49698 53282 49710
rect 53230 49634 53282 49646
rect 53790 49698 53842 49710
rect 53790 49634 53842 49646
rect 54238 49698 54290 49710
rect 54238 49634 54290 49646
rect 54574 49698 54626 49710
rect 54574 49634 54626 49646
rect 55134 49698 55186 49710
rect 55134 49634 55186 49646
rect 55470 49698 55522 49710
rect 55470 49634 55522 49646
rect 22542 49586 22594 49598
rect 22542 49522 22594 49534
rect 23438 49586 23490 49598
rect 23438 49522 23490 49534
rect 24110 49586 24162 49598
rect 33966 49586 34018 49598
rect 40014 49586 40066 49598
rect 27234 49534 27246 49586
rect 27298 49534 27310 49586
rect 33618 49534 33630 49586
rect 33682 49534 33694 49586
rect 35634 49534 35646 49586
rect 35698 49534 35710 49586
rect 38994 49534 39006 49586
rect 39058 49583 39070 49586
rect 39554 49583 39566 49586
rect 39058 49537 39566 49583
rect 39058 49534 39070 49537
rect 39554 49534 39566 49537
rect 39618 49534 39630 49586
rect 24110 49522 24162 49534
rect 33966 49522 34018 49534
rect 40014 49522 40066 49534
rect 40238 49586 40290 49598
rect 40238 49522 40290 49534
rect 43934 49586 43986 49598
rect 49410 49534 49422 49586
rect 49474 49583 49486 49586
rect 50306 49583 50318 49586
rect 49474 49537 50318 49583
rect 49474 49534 49486 49537
rect 50306 49534 50318 49537
rect 50370 49534 50382 49586
rect 43934 49522 43986 49534
rect 1344 49418 58576 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 58576 49418
rect 1344 49332 58576 49366
rect 13918 49250 13970 49262
rect 13918 49186 13970 49198
rect 23438 49250 23490 49262
rect 23438 49186 23490 49198
rect 23774 49250 23826 49262
rect 32734 49250 32786 49262
rect 26114 49198 26126 49250
rect 26178 49198 26190 49250
rect 23774 49186 23826 49198
rect 32734 49186 32786 49198
rect 33294 49250 33346 49262
rect 33294 49186 33346 49198
rect 39902 49250 39954 49262
rect 39902 49186 39954 49198
rect 46174 49250 46226 49262
rect 46174 49186 46226 49198
rect 48078 49250 48130 49262
rect 48078 49186 48130 49198
rect 48190 49250 48242 49262
rect 48190 49186 48242 49198
rect 15822 49138 15874 49150
rect 15822 49074 15874 49086
rect 20862 49138 20914 49150
rect 33742 49138 33794 49150
rect 43710 49138 43762 49150
rect 46958 49138 47010 49150
rect 21746 49086 21758 49138
rect 21810 49086 21822 49138
rect 26786 49086 26798 49138
rect 26850 49086 26862 49138
rect 31266 49086 31278 49138
rect 31330 49086 31342 49138
rect 40114 49086 40126 49138
rect 40178 49086 40190 49138
rect 46386 49086 46398 49138
rect 46450 49086 46462 49138
rect 20862 49074 20914 49086
rect 33742 49074 33794 49086
rect 43710 49074 43762 49086
rect 46958 49074 47010 49086
rect 47742 49138 47794 49150
rect 51102 49138 51154 49150
rect 49970 49086 49982 49138
rect 50034 49086 50046 49138
rect 47742 49074 47794 49086
rect 51102 49074 51154 49086
rect 51998 49138 52050 49150
rect 51998 49074 52050 49086
rect 9662 49026 9714 49038
rect 9662 48962 9714 48974
rect 12798 49026 12850 49038
rect 14142 49026 14194 49038
rect 13682 48974 13694 49026
rect 13746 48974 13758 49026
rect 12798 48962 12850 48974
rect 14142 48962 14194 48974
rect 16046 49026 16098 49038
rect 16046 48962 16098 48974
rect 16942 49026 16994 49038
rect 30270 49026 30322 49038
rect 21634 48974 21646 49026
rect 21698 48974 21710 49026
rect 26898 48974 26910 49026
rect 26962 48974 26974 49026
rect 16942 48962 16994 48974
rect 30270 48962 30322 48974
rect 30606 49026 30658 49038
rect 30606 48962 30658 48974
rect 32398 49026 32450 49038
rect 32398 48962 32450 48974
rect 33518 49026 33570 49038
rect 33518 48962 33570 48974
rect 34190 49026 34242 49038
rect 34190 48962 34242 48974
rect 35086 49026 35138 49038
rect 37886 49026 37938 49038
rect 35522 48974 35534 49026
rect 35586 48974 35598 49026
rect 35086 48962 35138 48974
rect 37886 48962 37938 48974
rect 39230 49026 39282 49038
rect 39230 48962 39282 48974
rect 40014 49026 40066 49038
rect 40014 48962 40066 48974
rect 40462 49026 40514 49038
rect 40462 48962 40514 48974
rect 40686 49026 40738 49038
rect 40686 48962 40738 48974
rect 43934 49026 43986 49038
rect 43934 48962 43986 48974
rect 46734 49026 46786 49038
rect 46734 48962 46786 48974
rect 47854 49026 47906 49038
rect 47854 48962 47906 48974
rect 49534 49026 49586 49038
rect 50418 48974 50430 49026
rect 50482 48974 50494 49026
rect 55122 48974 55134 49026
rect 55186 48974 55198 49026
rect 49534 48962 49586 48974
rect 10110 48914 10162 48926
rect 10110 48850 10162 48862
rect 10334 48914 10386 48926
rect 10334 48850 10386 48862
rect 12462 48914 12514 48926
rect 12462 48850 12514 48862
rect 12686 48914 12738 48926
rect 12686 48850 12738 48862
rect 17054 48914 17106 48926
rect 17054 48850 17106 48862
rect 18958 48914 19010 48926
rect 18958 48850 19010 48862
rect 21982 48914 22034 48926
rect 21982 48850 22034 48862
rect 23662 48914 23714 48926
rect 23662 48850 23714 48862
rect 29598 48914 29650 48926
rect 29598 48850 29650 48862
rect 30046 48914 30098 48926
rect 30046 48850 30098 48862
rect 31614 48914 31666 48926
rect 31614 48850 31666 48862
rect 32174 48914 32226 48926
rect 32174 48850 32226 48862
rect 34862 48914 34914 48926
rect 34862 48850 34914 48862
rect 41694 48914 41746 48926
rect 41694 48850 41746 48862
rect 42478 48914 42530 48926
rect 42478 48850 42530 48862
rect 43374 48914 43426 48926
rect 43374 48850 43426 48862
rect 45390 48914 45442 48926
rect 45390 48850 45442 48862
rect 46398 48914 46450 48926
rect 46398 48850 46450 48862
rect 48638 48914 48690 48926
rect 56018 48862 56030 48914
rect 56082 48862 56094 48914
rect 48638 48850 48690 48862
rect 9998 48802 10050 48814
rect 9998 48738 10050 48750
rect 12910 48802 12962 48814
rect 12910 48738 12962 48750
rect 13806 48802 13858 48814
rect 17278 48802 17330 48814
rect 16370 48750 16382 48802
rect 16434 48750 16446 48802
rect 13806 48738 13858 48750
rect 17278 48738 17330 48750
rect 18734 48802 18786 48814
rect 18734 48738 18786 48750
rect 18846 48802 18898 48814
rect 18846 48738 18898 48750
rect 22430 48802 22482 48814
rect 22430 48738 22482 48750
rect 22878 48802 22930 48814
rect 22878 48738 22930 48750
rect 30270 48802 30322 48814
rect 30270 48738 30322 48750
rect 31390 48802 31442 48814
rect 31390 48738 31442 48750
rect 33966 48802 34018 48814
rect 33966 48738 34018 48750
rect 34078 48802 34130 48814
rect 34078 48738 34130 48750
rect 35198 48802 35250 48814
rect 35198 48738 35250 48750
rect 35310 48802 35362 48814
rect 35310 48738 35362 48750
rect 35982 48802 36034 48814
rect 35982 48738 36034 48750
rect 36654 48802 36706 48814
rect 36654 48738 36706 48750
rect 37550 48802 37602 48814
rect 37550 48738 37602 48750
rect 38334 48802 38386 48814
rect 38334 48738 38386 48750
rect 39342 48802 39394 48814
rect 39342 48738 39394 48750
rect 41246 48802 41298 48814
rect 41246 48738 41298 48750
rect 42814 48802 42866 48814
rect 42814 48738 42866 48750
rect 43598 48802 43650 48814
rect 43598 48738 43650 48750
rect 43822 48802 43874 48814
rect 43822 48738 43874 48750
rect 44494 48802 44546 48814
rect 44494 48738 44546 48750
rect 51550 48802 51602 48814
rect 51550 48738 51602 48750
rect 52782 48802 52834 48814
rect 52782 48738 52834 48750
rect 53454 48802 53506 48814
rect 53454 48738 53506 48750
rect 53902 48802 53954 48814
rect 53902 48738 53954 48750
rect 54350 48802 54402 48814
rect 54350 48738 54402 48750
rect 1344 48634 58576 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 58576 48634
rect 1344 48548 58576 48582
rect 3278 48466 3330 48478
rect 17726 48466 17778 48478
rect 9762 48414 9774 48466
rect 9826 48414 9838 48466
rect 3278 48402 3330 48414
rect 17726 48402 17778 48414
rect 17950 48466 18002 48478
rect 17950 48402 18002 48414
rect 21198 48466 21250 48478
rect 21198 48402 21250 48414
rect 21870 48466 21922 48478
rect 21870 48402 21922 48414
rect 31390 48466 31442 48478
rect 31390 48402 31442 48414
rect 32734 48466 32786 48478
rect 32734 48402 32786 48414
rect 34526 48466 34578 48478
rect 39566 48466 39618 48478
rect 47070 48466 47122 48478
rect 37314 48414 37326 48466
rect 37378 48414 37390 48466
rect 40786 48414 40798 48466
rect 40850 48414 40862 48466
rect 43138 48414 43150 48466
rect 43202 48414 43214 48466
rect 34526 48402 34578 48414
rect 39566 48402 39618 48414
rect 47070 48402 47122 48414
rect 47182 48466 47234 48478
rect 47182 48402 47234 48414
rect 48078 48466 48130 48478
rect 48078 48402 48130 48414
rect 51662 48466 51714 48478
rect 51662 48402 51714 48414
rect 52334 48466 52386 48478
rect 52334 48402 52386 48414
rect 54238 48466 54290 48478
rect 54238 48402 54290 48414
rect 2382 48354 2434 48366
rect 2382 48290 2434 48302
rect 2718 48354 2770 48366
rect 2718 48290 2770 48302
rect 10446 48354 10498 48366
rect 10446 48290 10498 48302
rect 11790 48354 11842 48366
rect 11790 48290 11842 48302
rect 12462 48354 12514 48366
rect 18174 48354 18226 48366
rect 21982 48354 22034 48366
rect 14130 48302 14142 48354
rect 14194 48302 14206 48354
rect 18946 48302 18958 48354
rect 19010 48302 19022 48354
rect 12462 48290 12514 48302
rect 18174 48290 18226 48302
rect 21982 48290 22034 48302
rect 24334 48354 24386 48366
rect 24334 48290 24386 48302
rect 27134 48354 27186 48366
rect 27134 48290 27186 48302
rect 27246 48354 27298 48366
rect 27246 48290 27298 48302
rect 30830 48354 30882 48366
rect 30830 48290 30882 48302
rect 35870 48354 35922 48366
rect 35870 48290 35922 48302
rect 48638 48354 48690 48366
rect 48638 48290 48690 48302
rect 51326 48354 51378 48366
rect 51326 48290 51378 48302
rect 52782 48354 52834 48366
rect 52782 48290 52834 48302
rect 9774 48242 9826 48254
rect 9774 48178 9826 48190
rect 9998 48242 10050 48254
rect 9998 48178 10050 48190
rect 10222 48242 10274 48254
rect 10222 48178 10274 48190
rect 11678 48242 11730 48254
rect 11678 48178 11730 48190
rect 12014 48242 12066 48254
rect 23438 48242 23490 48254
rect 13122 48190 13134 48242
rect 13186 48190 13198 48242
rect 13794 48190 13806 48242
rect 13858 48190 13870 48242
rect 16594 48190 16606 48242
rect 16658 48190 16670 48242
rect 18834 48190 18846 48242
rect 18898 48190 18910 48242
rect 19730 48190 19742 48242
rect 19794 48190 19806 48242
rect 23202 48190 23214 48242
rect 23266 48190 23278 48242
rect 12014 48178 12066 48190
rect 23438 48178 23490 48190
rect 24110 48242 24162 48254
rect 24110 48178 24162 48190
rect 24446 48242 24498 48254
rect 24446 48178 24498 48190
rect 26910 48242 26962 48254
rect 26910 48178 26962 48190
rect 29710 48242 29762 48254
rect 29710 48178 29762 48190
rect 30494 48242 30546 48254
rect 30494 48178 30546 48190
rect 31726 48242 31778 48254
rect 31726 48178 31778 48190
rect 35758 48242 35810 48254
rect 35758 48178 35810 48190
rect 36990 48242 37042 48254
rect 40126 48242 40178 48254
rect 39330 48190 39342 48242
rect 39394 48190 39406 48242
rect 36990 48178 37042 48190
rect 40126 48178 40178 48190
rect 40350 48242 40402 48254
rect 40350 48178 40402 48190
rect 40574 48242 40626 48254
rect 40574 48178 40626 48190
rect 40798 48242 40850 48254
rect 46958 48242 47010 48254
rect 47854 48242 47906 48254
rect 46722 48190 46734 48242
rect 46786 48190 46798 48242
rect 47394 48190 47406 48242
rect 47458 48190 47470 48242
rect 40798 48178 40850 48190
rect 46958 48178 47010 48190
rect 47854 48178 47906 48190
rect 48190 48242 48242 48254
rect 51550 48242 51602 48254
rect 50306 48190 50318 48242
rect 50370 48190 50382 48242
rect 48190 48178 48242 48190
rect 51550 48178 51602 48190
rect 51774 48242 51826 48254
rect 53442 48190 53454 48242
rect 53506 48190 53518 48242
rect 51774 48178 51826 48190
rect 15150 48130 15202 48142
rect 15150 48066 15202 48078
rect 15934 48130 15986 48142
rect 17838 48130 17890 48142
rect 23550 48130 23602 48142
rect 16258 48078 16270 48130
rect 16322 48078 16334 48130
rect 19506 48078 19518 48130
rect 19570 48078 19582 48130
rect 15934 48066 15986 48078
rect 17838 48066 17890 48078
rect 23550 48066 23602 48078
rect 24894 48130 24946 48142
rect 24894 48066 24946 48078
rect 26126 48130 26178 48142
rect 26126 48066 26178 48078
rect 29934 48130 29986 48142
rect 33630 48130 33682 48142
rect 32834 48078 32846 48130
rect 32898 48078 32910 48130
rect 29934 48066 29986 48078
rect 33630 48066 33682 48078
rect 34862 48130 34914 48142
rect 34862 48066 34914 48078
rect 38222 48130 38274 48142
rect 38222 48066 38274 48078
rect 38670 48130 38722 48142
rect 38670 48066 38722 48078
rect 41582 48130 41634 48142
rect 41582 48066 41634 48078
rect 41918 48130 41970 48142
rect 41918 48066 41970 48078
rect 42366 48130 42418 48142
rect 42366 48066 42418 48078
rect 43710 48130 43762 48142
rect 43710 48066 43762 48078
rect 44158 48130 44210 48142
rect 44158 48066 44210 48078
rect 44606 48130 44658 48142
rect 44606 48066 44658 48078
rect 45054 48130 45106 48142
rect 45054 48066 45106 48078
rect 45502 48130 45554 48142
rect 45502 48066 45554 48078
rect 46062 48130 46114 48142
rect 46062 48066 46114 48078
rect 49646 48130 49698 48142
rect 54798 48130 54850 48142
rect 49970 48078 49982 48130
rect 50034 48078 50046 48130
rect 53666 48078 53678 48130
rect 53730 48078 53742 48130
rect 49646 48066 49698 48078
rect 54798 48066 54850 48078
rect 55246 48130 55298 48142
rect 55246 48066 55298 48078
rect 55582 48130 55634 48142
rect 55582 48066 55634 48078
rect 56030 48130 56082 48142
rect 56030 48066 56082 48078
rect 56478 48130 56530 48142
rect 56478 48066 56530 48078
rect 57486 48130 57538 48142
rect 57486 48066 57538 48078
rect 21870 48018 21922 48030
rect 21870 47954 21922 47966
rect 26686 48018 26738 48030
rect 26686 47954 26738 47966
rect 27470 48018 27522 48030
rect 32510 48018 32562 48030
rect 29362 47966 29374 48018
rect 29426 47966 29438 48018
rect 27470 47954 27522 47966
rect 32510 47954 32562 47966
rect 33854 48018 33906 48030
rect 33854 47954 33906 47966
rect 34078 48018 34130 48030
rect 34078 47954 34130 47966
rect 35534 48018 35586 48030
rect 35534 47954 35586 47966
rect 36094 48018 36146 48030
rect 36094 47954 36146 47966
rect 36318 48018 36370 48030
rect 36318 47954 36370 47966
rect 43486 48018 43538 48030
rect 43486 47954 43538 47966
rect 1344 47850 58576 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 58576 47850
rect 1344 47764 58576 47798
rect 8990 47682 9042 47694
rect 8990 47618 9042 47630
rect 11454 47682 11506 47694
rect 22318 47682 22370 47694
rect 40238 47682 40290 47694
rect 14466 47630 14478 47682
rect 14530 47630 14542 47682
rect 16594 47630 16606 47682
rect 16658 47630 16670 47682
rect 19618 47630 19630 47682
rect 19682 47630 19694 47682
rect 34738 47630 34750 47682
rect 34802 47679 34814 47682
rect 35074 47679 35086 47682
rect 34802 47633 35086 47679
rect 34802 47630 34814 47633
rect 35074 47630 35086 47633
rect 35138 47630 35150 47682
rect 39106 47630 39118 47682
rect 39170 47630 39182 47682
rect 11454 47618 11506 47630
rect 22318 47618 22370 47630
rect 40238 47618 40290 47630
rect 54238 47682 54290 47694
rect 54238 47618 54290 47630
rect 8766 47570 8818 47582
rect 18286 47570 18338 47582
rect 22878 47570 22930 47582
rect 26462 47570 26514 47582
rect 10322 47518 10334 47570
rect 10386 47518 10398 47570
rect 16706 47518 16718 47570
rect 16770 47518 16782 47570
rect 19506 47518 19518 47570
rect 19570 47518 19582 47570
rect 25554 47518 25566 47570
rect 25618 47518 25630 47570
rect 8766 47506 8818 47518
rect 18286 47506 18338 47518
rect 22878 47506 22930 47518
rect 26462 47506 26514 47518
rect 33742 47570 33794 47582
rect 33742 47506 33794 47518
rect 34750 47570 34802 47582
rect 34750 47506 34802 47518
rect 35198 47570 35250 47582
rect 35198 47506 35250 47518
rect 36766 47570 36818 47582
rect 36766 47506 36818 47518
rect 41694 47570 41746 47582
rect 57038 47570 57090 47582
rect 51650 47518 51662 47570
rect 51714 47518 51726 47570
rect 41694 47506 41746 47518
rect 57038 47506 57090 47518
rect 57486 47570 57538 47582
rect 57486 47506 57538 47518
rect 57934 47570 57986 47582
rect 57934 47506 57986 47518
rect 12238 47458 12290 47470
rect 10434 47406 10446 47458
rect 10498 47406 10510 47458
rect 11442 47406 11454 47458
rect 11506 47406 11518 47458
rect 12238 47394 12290 47406
rect 12686 47458 12738 47470
rect 12686 47394 12738 47406
rect 12910 47458 12962 47470
rect 12910 47394 12962 47406
rect 13806 47458 13858 47470
rect 13806 47394 13858 47406
rect 14030 47458 14082 47470
rect 22654 47458 22706 47470
rect 16258 47406 16270 47458
rect 16322 47406 16334 47458
rect 19282 47406 19294 47458
rect 19346 47406 19358 47458
rect 14030 47394 14082 47406
rect 22654 47394 22706 47406
rect 23438 47458 23490 47470
rect 23438 47394 23490 47406
rect 23774 47458 23826 47470
rect 37550 47458 37602 47470
rect 39678 47458 39730 47470
rect 40910 47458 40962 47470
rect 26002 47406 26014 47458
rect 26066 47406 26078 47458
rect 30034 47406 30046 47458
rect 30098 47406 30110 47458
rect 31154 47406 31166 47458
rect 31218 47406 31230 47458
rect 33282 47406 33294 47458
rect 33346 47406 33358 47458
rect 37762 47406 37774 47458
rect 37826 47406 37838 47458
rect 37986 47406 37998 47458
rect 38050 47406 38062 47458
rect 39442 47406 39454 47458
rect 39506 47406 39518 47458
rect 40674 47406 40686 47458
rect 40738 47406 40750 47458
rect 23774 47394 23826 47406
rect 37550 47394 37602 47406
rect 39678 47394 39730 47406
rect 40910 47394 40962 47406
rect 41134 47458 41186 47470
rect 48862 47458 48914 47470
rect 51886 47458 51938 47470
rect 43026 47406 43038 47458
rect 43090 47406 43102 47458
rect 43474 47406 43486 47458
rect 43538 47406 43550 47458
rect 44034 47406 44046 47458
rect 44098 47406 44110 47458
rect 46498 47406 46510 47458
rect 46562 47406 46574 47458
rect 47842 47406 47854 47458
rect 47906 47406 47918 47458
rect 49634 47406 49646 47458
rect 49698 47406 49710 47458
rect 51538 47406 51550 47458
rect 51602 47406 51614 47458
rect 41134 47394 41186 47406
rect 48862 47394 48914 47406
rect 51886 47394 51938 47406
rect 53566 47458 53618 47470
rect 53566 47394 53618 47406
rect 54014 47458 54066 47470
rect 54014 47394 54066 47406
rect 9886 47346 9938 47358
rect 9886 47282 9938 47294
rect 11790 47346 11842 47358
rect 11790 47282 11842 47294
rect 13918 47346 13970 47358
rect 13918 47282 13970 47294
rect 23550 47346 23602 47358
rect 33630 47346 33682 47358
rect 30930 47294 30942 47346
rect 30994 47294 31006 47346
rect 23550 47282 23602 47294
rect 33630 47282 33682 47294
rect 33854 47346 33906 47358
rect 33854 47282 33906 47294
rect 34302 47346 34354 47358
rect 34302 47282 34354 47294
rect 41022 47346 41074 47358
rect 53454 47346 53506 47358
rect 43698 47294 43710 47346
rect 43762 47294 43774 47346
rect 44370 47294 44382 47346
rect 44434 47294 44446 47346
rect 46834 47294 46846 47346
rect 46898 47294 46910 47346
rect 41022 47282 41074 47294
rect 53454 47282 53506 47294
rect 53790 47346 53842 47358
rect 53790 47282 53842 47294
rect 54910 47346 54962 47358
rect 54910 47282 54962 47294
rect 55246 47346 55298 47358
rect 55246 47282 55298 47294
rect 12574 47234 12626 47246
rect 9314 47182 9326 47234
rect 9378 47182 9390 47234
rect 12574 47170 12626 47182
rect 14926 47234 14978 47246
rect 14926 47170 14978 47182
rect 17950 47234 18002 47246
rect 17950 47170 18002 47182
rect 18174 47234 18226 47246
rect 18174 47170 18226 47182
rect 18398 47234 18450 47246
rect 18398 47170 18450 47182
rect 24110 47234 24162 47246
rect 35646 47234 35698 47246
rect 30146 47182 30158 47234
rect 30210 47182 30222 47234
rect 24110 47170 24162 47182
rect 35646 47170 35698 47182
rect 36318 47234 36370 47246
rect 36318 47170 36370 47182
rect 42254 47234 42306 47246
rect 42254 47170 42306 47182
rect 45390 47234 45442 47246
rect 45390 47170 45442 47182
rect 46062 47234 46114 47246
rect 52558 47234 52610 47246
rect 51314 47182 51326 47234
rect 51378 47182 51390 47234
rect 46062 47170 46114 47182
rect 52558 47170 52610 47182
rect 55694 47234 55746 47246
rect 55694 47170 55746 47182
rect 56142 47234 56194 47246
rect 56142 47170 56194 47182
rect 56590 47234 56642 47246
rect 56590 47170 56642 47182
rect 1344 47066 58576 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 58576 47066
rect 1344 46980 58576 47014
rect 12798 46898 12850 46910
rect 16830 46898 16882 46910
rect 14354 46846 14366 46898
rect 14418 46846 14430 46898
rect 12798 46834 12850 46846
rect 16830 46834 16882 46846
rect 17054 46898 17106 46910
rect 17054 46834 17106 46846
rect 18286 46898 18338 46910
rect 18286 46834 18338 46846
rect 22654 46898 22706 46910
rect 22654 46834 22706 46846
rect 22878 46898 22930 46910
rect 22878 46834 22930 46846
rect 23214 46898 23266 46910
rect 23214 46834 23266 46846
rect 24894 46898 24946 46910
rect 24894 46834 24946 46846
rect 34862 46898 34914 46910
rect 34862 46834 34914 46846
rect 40462 46898 40514 46910
rect 40462 46834 40514 46846
rect 40686 46898 40738 46910
rect 40686 46834 40738 46846
rect 43262 46898 43314 46910
rect 43262 46834 43314 46846
rect 44270 46898 44322 46910
rect 44270 46834 44322 46846
rect 48302 46898 48354 46910
rect 48302 46834 48354 46846
rect 49870 46898 49922 46910
rect 55694 46898 55746 46910
rect 53554 46846 53566 46898
rect 53618 46846 53630 46898
rect 54450 46846 54462 46898
rect 54514 46846 54526 46898
rect 49870 46834 49922 46846
rect 55694 46834 55746 46846
rect 56142 46898 56194 46910
rect 56142 46834 56194 46846
rect 16718 46786 16770 46798
rect 16718 46722 16770 46734
rect 18510 46786 18562 46798
rect 18510 46722 18562 46734
rect 26910 46786 26962 46798
rect 26910 46722 26962 46734
rect 33742 46786 33794 46798
rect 33742 46722 33794 46734
rect 33966 46786 34018 46798
rect 33966 46722 34018 46734
rect 36878 46786 36930 46798
rect 36878 46722 36930 46734
rect 39566 46786 39618 46798
rect 45054 46786 45106 46798
rect 42914 46734 42926 46786
rect 42978 46734 42990 46786
rect 39566 46722 39618 46734
rect 45054 46722 45106 46734
rect 46734 46786 46786 46798
rect 46734 46722 46786 46734
rect 51998 46786 52050 46798
rect 51998 46722 52050 46734
rect 57822 46786 57874 46798
rect 57822 46722 57874 46734
rect 14030 46674 14082 46686
rect 10098 46622 10110 46674
rect 10162 46622 10174 46674
rect 14030 46610 14082 46622
rect 18622 46674 18674 46686
rect 22542 46674 22594 46686
rect 19618 46622 19630 46674
rect 19682 46622 19694 46674
rect 18622 46610 18674 46622
rect 22542 46610 22594 46622
rect 24222 46674 24274 46686
rect 24222 46610 24274 46622
rect 24670 46674 24722 46686
rect 34414 46674 34466 46686
rect 37774 46674 37826 46686
rect 40238 46674 40290 46686
rect 25890 46622 25902 46674
rect 25954 46622 25966 46674
rect 26114 46622 26126 46674
rect 26178 46622 26190 46674
rect 27234 46622 27246 46674
rect 27298 46622 27310 46674
rect 30258 46622 30270 46674
rect 30322 46622 30334 46674
rect 32386 46622 32398 46674
rect 32450 46622 32462 46674
rect 37538 46622 37550 46674
rect 37602 46622 37614 46674
rect 39330 46622 39342 46674
rect 39394 46622 39406 46674
rect 24670 46610 24722 46622
rect 34414 46610 34466 46622
rect 37774 46610 37826 46622
rect 40238 46610 40290 46622
rect 40350 46674 40402 46686
rect 40350 46610 40402 46622
rect 40574 46674 40626 46686
rect 43486 46674 43538 46686
rect 43026 46622 43038 46674
rect 43090 46622 43102 46674
rect 40574 46610 40626 46622
rect 43486 46610 43538 46622
rect 44046 46674 44098 46686
rect 48414 46674 48466 46686
rect 52894 46674 52946 46686
rect 44594 46622 44606 46674
rect 44658 46622 44670 46674
rect 47282 46622 47294 46674
rect 47346 46622 47358 46674
rect 48066 46622 48078 46674
rect 48130 46622 48142 46674
rect 49634 46622 49646 46674
rect 49698 46622 49710 46674
rect 52434 46622 52446 46674
rect 52498 46622 52510 46674
rect 44046 46610 44098 46622
rect 48414 46610 48466 46622
rect 52894 46610 52946 46622
rect 53902 46674 53954 46686
rect 54674 46622 54686 46674
rect 54738 46622 54750 46674
rect 53902 46610 53954 46622
rect 9102 46562 9154 46574
rect 10782 46562 10834 46574
rect 10322 46510 10334 46562
rect 10386 46510 10398 46562
rect 9102 46498 9154 46510
rect 10782 46498 10834 46510
rect 13246 46562 13298 46574
rect 13246 46498 13298 46510
rect 13806 46562 13858 46574
rect 24782 46562 24834 46574
rect 38334 46562 38386 46574
rect 19730 46510 19742 46562
rect 19794 46510 19806 46562
rect 26450 46510 26462 46562
rect 26514 46510 26526 46562
rect 27346 46510 27358 46562
rect 27410 46510 27422 46562
rect 30034 46510 30046 46562
rect 30098 46510 30110 46562
rect 32498 46510 32510 46562
rect 32562 46510 32574 46562
rect 33618 46510 33630 46562
rect 33682 46510 33694 46562
rect 13806 46498 13858 46510
rect 24782 46498 24834 46510
rect 38334 46498 38386 46510
rect 41470 46562 41522 46574
rect 41470 46498 41522 46510
rect 42254 46562 42306 46574
rect 44158 46562 44210 46574
rect 42690 46510 42702 46562
rect 42754 46510 42766 46562
rect 42254 46498 42306 46510
rect 44158 46498 44210 46510
rect 45614 46562 45666 46574
rect 45614 46498 45666 46510
rect 45950 46562 46002 46574
rect 50318 46562 50370 46574
rect 47394 46510 47406 46562
rect 47458 46510 47470 46562
rect 45950 46498 46002 46510
rect 50318 46498 50370 46510
rect 50878 46562 50930 46574
rect 50878 46498 50930 46510
rect 51214 46562 51266 46574
rect 51214 46498 51266 46510
rect 55358 46562 55410 46574
rect 55358 46498 55410 46510
rect 56590 46562 56642 46574
rect 56590 46498 56642 46510
rect 57374 46562 57426 46574
rect 57374 46498 57426 46510
rect 20178 46398 20190 46450
rect 20242 46398 20254 46450
rect 29922 46398 29934 46450
rect 29986 46398 29998 46450
rect 31826 46398 31838 46450
rect 31890 46398 31902 46450
rect 1344 46282 58576 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 58576 46282
rect 1344 46196 58576 46230
rect 12350 46114 12402 46126
rect 19182 46114 19234 46126
rect 52670 46114 52722 46126
rect 13682 46062 13694 46114
rect 13746 46062 13758 46114
rect 23314 46062 23326 46114
rect 23378 46062 23390 46114
rect 25442 46062 25454 46114
rect 25506 46062 25518 46114
rect 57250 46062 57262 46114
rect 57314 46111 57326 46114
rect 58034 46111 58046 46114
rect 57314 46065 58046 46111
rect 57314 46062 57326 46065
rect 58034 46062 58046 46065
rect 58098 46062 58110 46114
rect 12350 46050 12402 46062
rect 19182 46050 19234 46062
rect 52670 46050 52722 46062
rect 6414 46002 6466 46014
rect 27022 46002 27074 46014
rect 41694 46002 41746 46014
rect 10098 45950 10110 46002
rect 10162 45950 10174 46002
rect 22866 45950 22878 46002
rect 22930 45950 22942 46002
rect 26114 45950 26126 46002
rect 26178 45950 26190 46002
rect 29810 45950 29822 46002
rect 29874 45950 29886 46002
rect 35298 45950 35310 46002
rect 35362 45950 35374 46002
rect 6414 45938 6466 45950
rect 27022 45938 27074 45950
rect 41694 45938 41746 45950
rect 42926 46002 42978 46014
rect 48862 46002 48914 46014
rect 43698 45950 43710 46002
rect 43762 45950 43774 46002
rect 46946 45950 46958 46002
rect 47010 45950 47022 46002
rect 47170 45950 47182 46002
rect 47234 45950 47246 46002
rect 42926 45938 42978 45950
rect 48862 45938 48914 45950
rect 50318 46002 50370 46014
rect 50318 45938 50370 45950
rect 50766 46002 50818 46014
rect 50766 45938 50818 45950
rect 51214 46002 51266 46014
rect 51214 45938 51266 45950
rect 57262 46002 57314 46014
rect 57262 45938 57314 45950
rect 12686 45890 12738 45902
rect 2818 45838 2830 45890
rect 2882 45838 2894 45890
rect 12686 45826 12738 45838
rect 14030 45890 14082 45902
rect 14030 45826 14082 45838
rect 14254 45890 14306 45902
rect 24894 45890 24946 45902
rect 22978 45838 22990 45890
rect 23042 45838 23054 45890
rect 14254 45826 14306 45838
rect 24894 45826 24946 45838
rect 25118 45890 25170 45902
rect 28254 45890 28306 45902
rect 26562 45838 26574 45890
rect 26626 45838 26638 45890
rect 25118 45826 25170 45838
rect 28254 45826 28306 45838
rect 28478 45890 28530 45902
rect 28478 45826 28530 45838
rect 28926 45890 28978 45902
rect 37774 45890 37826 45902
rect 29922 45838 29934 45890
rect 29986 45838 29998 45890
rect 28926 45826 28978 45838
rect 37774 45826 37826 45838
rect 39118 45890 39170 45902
rect 48414 45890 48466 45902
rect 43474 45838 43486 45890
rect 43538 45838 43550 45890
rect 46610 45838 46622 45890
rect 46674 45838 46686 45890
rect 47506 45838 47518 45890
rect 47570 45838 47582 45890
rect 49746 45838 49758 45890
rect 49810 45838 49822 45890
rect 39118 45826 39170 45838
rect 48414 45826 48466 45838
rect 5854 45778 5906 45790
rect 1922 45726 1934 45778
rect 1986 45726 1998 45778
rect 5854 45714 5906 45726
rect 5966 45778 6018 45790
rect 12910 45778 12962 45790
rect 9090 45726 9102 45778
rect 9154 45726 9166 45778
rect 5966 45714 6018 45726
rect 12910 45714 12962 45726
rect 19518 45778 19570 45790
rect 19518 45714 19570 45726
rect 19966 45778 20018 45790
rect 19966 45714 20018 45726
rect 30606 45778 30658 45790
rect 40014 45778 40066 45790
rect 36642 45726 36654 45778
rect 36706 45726 36718 45778
rect 30606 45714 30658 45726
rect 40014 45714 40066 45726
rect 40350 45778 40402 45790
rect 40350 45714 40402 45726
rect 45726 45778 45778 45790
rect 45726 45714 45778 45726
rect 47966 45778 48018 45790
rect 52558 45778 52610 45790
rect 49522 45726 49534 45778
rect 49586 45726 49598 45778
rect 47966 45714 48018 45726
rect 52558 45714 52610 45726
rect 53454 45778 53506 45790
rect 53454 45714 53506 45726
rect 5630 45666 5682 45678
rect 5630 45602 5682 45614
rect 7310 45666 7362 45678
rect 7310 45602 7362 45614
rect 8206 45666 8258 45678
rect 8206 45602 8258 45614
rect 10558 45666 10610 45678
rect 10558 45602 10610 45614
rect 11118 45666 11170 45678
rect 11118 45602 11170 45614
rect 11790 45666 11842 45678
rect 11790 45602 11842 45614
rect 14702 45666 14754 45678
rect 14702 45602 14754 45614
rect 19294 45666 19346 45678
rect 19294 45602 19346 45614
rect 28366 45666 28418 45678
rect 28366 45602 28418 45614
rect 33070 45666 33122 45678
rect 33070 45602 33122 45614
rect 33630 45666 33682 45678
rect 33630 45602 33682 45614
rect 37438 45666 37490 45678
rect 37438 45602 37490 45614
rect 37662 45666 37714 45678
rect 37662 45602 37714 45614
rect 38222 45666 38274 45678
rect 38222 45602 38274 45614
rect 38782 45666 38834 45678
rect 38782 45602 38834 45614
rect 40798 45666 40850 45678
rect 40798 45602 40850 45614
rect 41246 45666 41298 45678
rect 41246 45602 41298 45614
rect 42254 45666 42306 45678
rect 42254 45602 42306 45614
rect 44382 45666 44434 45678
rect 44382 45602 44434 45614
rect 45614 45666 45666 45678
rect 45614 45602 45666 45614
rect 52110 45666 52162 45678
rect 54238 45666 54290 45678
rect 53778 45614 53790 45666
rect 53842 45614 53854 45666
rect 52110 45602 52162 45614
rect 54238 45602 54290 45614
rect 54798 45666 54850 45678
rect 54798 45602 54850 45614
rect 55246 45666 55298 45678
rect 55246 45602 55298 45614
rect 55806 45666 55858 45678
rect 55806 45602 55858 45614
rect 56254 45666 56306 45678
rect 56254 45602 56306 45614
rect 56590 45666 56642 45678
rect 56590 45602 56642 45614
rect 57598 45666 57650 45678
rect 57598 45602 57650 45614
rect 58046 45666 58098 45678
rect 58046 45602 58098 45614
rect 1344 45498 58576 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 58576 45498
rect 1344 45412 58576 45446
rect 2382 45330 2434 45342
rect 2382 45266 2434 45278
rect 3278 45330 3330 45342
rect 13022 45330 13074 45342
rect 8418 45278 8430 45330
rect 8482 45278 8494 45330
rect 3278 45266 3330 45278
rect 13022 45266 13074 45278
rect 13582 45330 13634 45342
rect 13582 45266 13634 45278
rect 19182 45330 19234 45342
rect 19182 45266 19234 45278
rect 19406 45330 19458 45342
rect 19406 45266 19458 45278
rect 20302 45330 20354 45342
rect 20302 45266 20354 45278
rect 23214 45330 23266 45342
rect 23214 45266 23266 45278
rect 26574 45330 26626 45342
rect 37214 45330 37266 45342
rect 30258 45278 30270 45330
rect 30322 45278 30334 45330
rect 26574 45266 26626 45278
rect 37214 45266 37266 45278
rect 42366 45330 42418 45342
rect 53230 45330 53282 45342
rect 47506 45278 47518 45330
rect 47570 45278 47582 45330
rect 52434 45278 52446 45330
rect 52498 45278 52510 45330
rect 42366 45266 42418 45278
rect 53230 45266 53282 45278
rect 2718 45218 2770 45230
rect 12014 45218 12066 45230
rect 9762 45166 9774 45218
rect 9826 45166 9838 45218
rect 2718 45154 2770 45166
rect 12014 45154 12066 45166
rect 12574 45218 12626 45230
rect 12574 45154 12626 45166
rect 13134 45218 13186 45230
rect 13134 45154 13186 45166
rect 16718 45218 16770 45230
rect 16718 45154 16770 45166
rect 22878 45218 22930 45230
rect 22878 45154 22930 45166
rect 22990 45218 23042 45230
rect 22990 45154 23042 45166
rect 25902 45218 25954 45230
rect 25902 45154 25954 45166
rect 29710 45218 29762 45230
rect 29710 45154 29762 45166
rect 36430 45218 36482 45230
rect 36430 45154 36482 45166
rect 40686 45218 40738 45230
rect 48078 45218 48130 45230
rect 43922 45166 43934 45218
rect 43986 45166 43998 45218
rect 44594 45166 44606 45218
rect 44658 45166 44670 45218
rect 45490 45166 45502 45218
rect 45554 45166 45566 45218
rect 40686 45154 40738 45166
rect 48078 45154 48130 45166
rect 54014 45218 54066 45230
rect 54014 45154 54066 45166
rect 57486 45218 57538 45230
rect 57486 45154 57538 45166
rect 57822 45218 57874 45230
rect 57822 45154 57874 45166
rect 10110 45106 10162 45118
rect 5394 45054 5406 45106
rect 5458 45054 5470 45106
rect 5842 45054 5854 45106
rect 5906 45054 5918 45106
rect 10110 45042 10162 45054
rect 12798 45106 12850 45118
rect 18510 45106 18562 45118
rect 16258 45054 16270 45106
rect 16322 45054 16334 45106
rect 12798 45042 12850 45054
rect 18510 45042 18562 45054
rect 19070 45106 19122 45118
rect 19070 45042 19122 45054
rect 19966 45106 20018 45118
rect 19966 45042 20018 45054
rect 29934 45106 29986 45118
rect 31726 45106 31778 45118
rect 33742 45106 33794 45118
rect 39566 45106 39618 45118
rect 46286 45106 46338 45118
rect 47966 45106 48018 45118
rect 30818 45054 30830 45106
rect 30882 45054 30894 45106
rect 32610 45054 32622 45106
rect 32674 45054 32686 45106
rect 34178 45054 34190 45106
rect 34242 45054 34254 45106
rect 40450 45054 40462 45106
rect 40514 45054 40526 45106
rect 42690 45054 42702 45106
rect 42754 45054 42766 45106
rect 43810 45054 43822 45106
rect 43874 45054 43886 45106
rect 44482 45054 44494 45106
rect 44546 45054 44558 45106
rect 45602 45054 45614 45106
rect 45666 45054 45678 45106
rect 46498 45054 46510 45106
rect 46562 45054 46574 45106
rect 29934 45042 29986 45054
rect 31726 45042 31778 45054
rect 33742 45042 33794 45054
rect 39566 45042 39618 45054
rect 46286 45042 46338 45054
rect 47966 45042 48018 45054
rect 48190 45106 48242 45118
rect 48190 45042 48242 45054
rect 49534 45106 49586 45118
rect 53790 45106 53842 45118
rect 50082 45054 50094 45106
rect 50146 45054 50158 45106
rect 49534 45042 49586 45054
rect 53790 45042 53842 45054
rect 54462 45106 54514 45118
rect 54462 45042 54514 45054
rect 10894 44994 10946 45006
rect 10894 44930 10946 44942
rect 11566 44994 11618 45006
rect 11566 44930 11618 44942
rect 14030 44994 14082 45006
rect 14030 44930 14082 44942
rect 15262 44994 15314 45006
rect 17726 44994 17778 45006
rect 15922 44942 15934 44994
rect 15986 44942 15998 44994
rect 15262 44930 15314 44942
rect 17726 44930 17778 44942
rect 18062 44994 18114 45006
rect 18062 44930 18114 44942
rect 20302 44994 20354 45006
rect 20302 44930 20354 44942
rect 20862 44994 20914 45006
rect 20862 44930 20914 44942
rect 26686 44994 26738 45006
rect 26686 44930 26738 44942
rect 31054 44994 31106 45006
rect 37662 44994 37714 45006
rect 32162 44942 32174 44994
rect 32226 44942 32238 44994
rect 31054 44930 31106 44942
rect 37662 44930 37714 44942
rect 38334 44994 38386 45006
rect 38334 44930 38386 44942
rect 38894 44994 38946 45006
rect 38894 44930 38946 44942
rect 41470 44994 41522 45006
rect 41470 44930 41522 44942
rect 41918 44994 41970 45006
rect 48750 44994 48802 45006
rect 45378 44942 45390 44994
rect 45442 44942 45454 44994
rect 41918 44930 41970 44942
rect 48750 44930 48802 44942
rect 55022 44994 55074 45006
rect 55022 44930 55074 44942
rect 55582 44994 55634 45006
rect 55582 44930 55634 44942
rect 55918 44994 55970 45006
rect 55918 44930 55970 44942
rect 56366 44994 56418 45006
rect 56366 44930 56418 44942
rect 8990 44882 9042 44894
rect 8990 44818 9042 44830
rect 20190 44882 20242 44894
rect 20190 44818 20242 44830
rect 25678 44882 25730 44894
rect 25678 44818 25730 44830
rect 26014 44882 26066 44894
rect 26014 44818 26066 44830
rect 31166 44882 31218 44894
rect 31166 44818 31218 44830
rect 53678 44882 53730 44894
rect 53678 44818 53730 44830
rect 54238 44882 54290 44894
rect 54238 44818 54290 44830
rect 1344 44714 58576 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 58576 44714
rect 1344 44628 58576 44662
rect 5966 44546 6018 44558
rect 5966 44482 6018 44494
rect 24222 44546 24274 44558
rect 24222 44482 24274 44494
rect 36318 44546 36370 44558
rect 36318 44482 36370 44494
rect 42702 44546 42754 44558
rect 42702 44482 42754 44494
rect 46174 44546 46226 44558
rect 46174 44482 46226 44494
rect 47406 44546 47458 44558
rect 54350 44546 54402 44558
rect 49634 44494 49646 44546
rect 49698 44543 49710 44546
rect 49970 44543 49982 44546
rect 49698 44497 49982 44543
rect 49698 44494 49710 44497
rect 49970 44494 49982 44497
rect 50034 44494 50046 44546
rect 51986 44543 51998 44546
rect 51553 44497 51998 44543
rect 47406 44482 47458 44494
rect 10446 44434 10498 44446
rect 23214 44434 23266 44446
rect 40238 44434 40290 44446
rect 20626 44382 20638 44434
rect 20690 44382 20702 44434
rect 25554 44382 25566 44434
rect 25618 44382 25630 44434
rect 10446 44370 10498 44382
rect 23214 44370 23266 44382
rect 40238 44370 40290 44382
rect 41134 44434 41186 44446
rect 41134 44370 41186 44382
rect 43934 44434 43986 44446
rect 43934 44370 43986 44382
rect 47854 44434 47906 44446
rect 47854 44370 47906 44382
rect 7870 44322 7922 44334
rect 14254 44322 14306 44334
rect 15038 44322 15090 44334
rect 16494 44322 16546 44334
rect 8530 44270 8542 44322
rect 8594 44270 8606 44322
rect 14802 44270 14814 44322
rect 14866 44270 14878 44322
rect 15810 44270 15822 44322
rect 15874 44319 15886 44322
rect 16034 44319 16046 44322
rect 15874 44273 16046 44319
rect 15874 44270 15886 44273
rect 16034 44270 16046 44273
rect 16098 44270 16110 44322
rect 7870 44258 7922 44270
rect 14254 44258 14306 44270
rect 15038 44258 15090 44270
rect 16494 44258 16546 44270
rect 16942 44322 16994 44334
rect 16942 44258 16994 44270
rect 17838 44322 17890 44334
rect 17838 44258 17890 44270
rect 18174 44322 18226 44334
rect 18174 44258 18226 44270
rect 19742 44322 19794 44334
rect 23102 44322 23154 44334
rect 20402 44270 20414 44322
rect 20466 44270 20478 44322
rect 22754 44270 22766 44322
rect 22818 44270 22830 44322
rect 19742 44258 19794 44270
rect 23102 44258 23154 44270
rect 23662 44322 23714 44334
rect 23662 44258 23714 44270
rect 24334 44322 24386 44334
rect 24334 44258 24386 44270
rect 24558 44322 24610 44334
rect 24558 44258 24610 44270
rect 24670 44322 24722 44334
rect 26462 44322 26514 44334
rect 26002 44270 26014 44322
rect 26066 44270 26078 44322
rect 24670 44258 24722 44270
rect 26462 44258 26514 44270
rect 29934 44322 29986 44334
rect 29934 44258 29986 44270
rect 30382 44322 30434 44334
rect 30382 44258 30434 44270
rect 35422 44322 35474 44334
rect 35422 44258 35474 44270
rect 36430 44322 36482 44334
rect 36430 44258 36482 44270
rect 42926 44322 42978 44334
rect 46398 44322 46450 44334
rect 46050 44270 46062 44322
rect 46114 44270 46126 44322
rect 42926 44258 42978 44270
rect 46398 44258 46450 44270
rect 47182 44322 47234 44334
rect 47182 44258 47234 44270
rect 47630 44322 47682 44334
rect 47630 44258 47682 44270
rect 48638 44322 48690 44334
rect 48638 44258 48690 44270
rect 48862 44322 48914 44334
rect 48862 44258 48914 44270
rect 49086 44322 49138 44334
rect 50194 44270 50206 44322
rect 50258 44270 50270 44322
rect 51314 44270 51326 44322
rect 51378 44270 51390 44322
rect 49086 44258 49138 44270
rect 6078 44210 6130 44222
rect 6078 44146 6130 44158
rect 6638 44210 6690 44222
rect 6638 44146 6690 44158
rect 7534 44210 7586 44222
rect 7534 44146 7586 44158
rect 8766 44210 8818 44222
rect 8766 44146 8818 44158
rect 9326 44210 9378 44222
rect 9326 44146 9378 44158
rect 9662 44210 9714 44222
rect 9662 44146 9714 44158
rect 10558 44210 10610 44222
rect 10558 44146 10610 44158
rect 11118 44210 11170 44222
rect 11118 44146 11170 44158
rect 15150 44210 15202 44222
rect 15150 44146 15202 44158
rect 18398 44210 18450 44222
rect 18398 44146 18450 44158
rect 29598 44210 29650 44222
rect 29598 44146 29650 44158
rect 30942 44210 30994 44222
rect 30942 44146 30994 44158
rect 31278 44210 31330 44222
rect 31278 44146 31330 44158
rect 31502 44210 31554 44222
rect 31502 44146 31554 44158
rect 32174 44210 32226 44222
rect 32174 44146 32226 44158
rect 35086 44210 35138 44222
rect 35086 44146 35138 44158
rect 36318 44210 36370 44222
rect 36318 44146 36370 44158
rect 38894 44210 38946 44222
rect 38894 44146 38946 44158
rect 39342 44210 39394 44222
rect 39342 44146 39394 44158
rect 45838 44210 45890 44222
rect 45838 44146 45890 44158
rect 48414 44210 48466 44222
rect 50866 44158 50878 44210
rect 50930 44158 50942 44210
rect 48414 44146 48466 44158
rect 5070 44098 5122 44110
rect 5070 44034 5122 44046
rect 5966 44098 6018 44110
rect 5966 44034 6018 44046
rect 6750 44098 6802 44110
rect 6750 44034 6802 44046
rect 6862 44098 6914 44110
rect 6862 44034 6914 44046
rect 10334 44098 10386 44110
rect 10334 44034 10386 44046
rect 11454 44098 11506 44110
rect 11454 44034 11506 44046
rect 12014 44098 12066 44110
rect 12014 44034 12066 44046
rect 12910 44098 12962 44110
rect 16270 44098 16322 44110
rect 15586 44046 15598 44098
rect 15650 44046 15662 44098
rect 12910 44034 12962 44046
rect 16270 44034 16322 44046
rect 16382 44098 16434 44110
rect 16382 44034 16434 44046
rect 17278 44098 17330 44110
rect 17278 44034 17330 44046
rect 18062 44098 18114 44110
rect 18062 44034 18114 44046
rect 31166 44098 31218 44110
rect 31166 44034 31218 44046
rect 32734 44098 32786 44110
rect 32734 44034 32786 44046
rect 32846 44098 32898 44110
rect 32846 44034 32898 44046
rect 32958 44098 33010 44110
rect 32958 44034 33010 44046
rect 33182 44098 33234 44110
rect 33182 44034 33234 44046
rect 37438 44098 37490 44110
rect 37438 44034 37490 44046
rect 37998 44098 38050 44110
rect 37998 44034 38050 44046
rect 38334 44098 38386 44110
rect 38334 44034 38386 44046
rect 38782 44098 38834 44110
rect 38782 44034 38834 44046
rect 39118 44098 39170 44110
rect 39118 44034 39170 44046
rect 39902 44098 39954 44110
rect 39902 44034 39954 44046
rect 40686 44098 40738 44110
rect 40686 44034 40738 44046
rect 41694 44098 41746 44110
rect 41694 44034 41746 44046
rect 42366 44098 42418 44110
rect 42366 44034 42418 44046
rect 42590 44098 42642 44110
rect 42590 44034 42642 44046
rect 43598 44098 43650 44110
rect 43598 44034 43650 44046
rect 44494 44098 44546 44110
rect 44494 44034 44546 44046
rect 46734 44098 46786 44110
rect 46734 44034 46786 44046
rect 49646 44098 49698 44110
rect 51553 44098 51599 44497
rect 51986 44494 51998 44497
rect 52050 44494 52062 44546
rect 54350 44482 54402 44494
rect 52222 44434 52274 44446
rect 55458 44382 55470 44434
rect 55522 44382 55534 44434
rect 52222 44370 52274 44382
rect 53454 44322 53506 44334
rect 53454 44258 53506 44270
rect 53678 44322 53730 44334
rect 53678 44258 53730 44270
rect 53902 44322 53954 44334
rect 57486 44322 57538 44334
rect 55570 44270 55582 44322
rect 55634 44270 55646 44322
rect 53902 44258 53954 44270
rect 57486 44258 57538 44270
rect 55134 44210 55186 44222
rect 55134 44146 55186 44158
rect 51886 44098 51938 44110
rect 50418 44046 50430 44098
rect 50482 44046 50494 44098
rect 51538 44046 51550 44098
rect 51602 44046 51614 44098
rect 49646 44034 49698 44046
rect 51886 44034 51938 44046
rect 52670 44098 52722 44110
rect 52670 44034 52722 44046
rect 56590 44098 56642 44110
rect 56590 44034 56642 44046
rect 57150 44098 57202 44110
rect 57150 44034 57202 44046
rect 57934 44098 57986 44110
rect 57934 44034 57986 44046
rect 1344 43930 58576 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 58576 43930
rect 1344 43844 58576 43878
rect 6302 43762 6354 43774
rect 8990 43762 9042 43774
rect 5730 43710 5742 43762
rect 5794 43710 5806 43762
rect 8194 43710 8206 43762
rect 8258 43710 8270 43762
rect 6302 43698 6354 43710
rect 8990 43698 9042 43710
rect 15934 43762 15986 43774
rect 15934 43698 15986 43710
rect 16942 43762 16994 43774
rect 16942 43698 16994 43710
rect 18062 43762 18114 43774
rect 18062 43698 18114 43710
rect 19406 43762 19458 43774
rect 19406 43698 19458 43710
rect 20974 43762 21026 43774
rect 20974 43698 21026 43710
rect 25902 43762 25954 43774
rect 25902 43698 25954 43710
rect 26126 43762 26178 43774
rect 26126 43698 26178 43710
rect 34526 43762 34578 43774
rect 39566 43762 39618 43774
rect 38770 43710 38782 43762
rect 38834 43710 38846 43762
rect 41906 43710 41918 43762
rect 41970 43710 41982 43762
rect 46274 43710 46286 43762
rect 46338 43710 46350 43762
rect 34526 43698 34578 43710
rect 39566 43698 39618 43710
rect 7086 43650 7138 43662
rect 7086 43586 7138 43598
rect 7310 43650 7362 43662
rect 7310 43586 7362 43598
rect 11790 43650 11842 43662
rect 11790 43586 11842 43598
rect 13134 43650 13186 43662
rect 13134 43586 13186 43598
rect 13582 43650 13634 43662
rect 13582 43586 13634 43598
rect 14254 43650 14306 43662
rect 14254 43586 14306 43598
rect 16830 43650 16882 43662
rect 16830 43586 16882 43598
rect 18398 43650 18450 43662
rect 18398 43586 18450 43598
rect 18510 43650 18562 43662
rect 18510 43586 18562 43598
rect 22990 43650 23042 43662
rect 22990 43586 23042 43598
rect 23214 43650 23266 43662
rect 23214 43586 23266 43598
rect 25790 43650 25842 43662
rect 32286 43650 32338 43662
rect 28466 43598 28478 43650
rect 28530 43598 28542 43650
rect 25790 43586 25842 43598
rect 32286 43586 32338 43598
rect 40238 43650 40290 43662
rect 40238 43586 40290 43598
rect 40350 43650 40402 43662
rect 45054 43650 45106 43662
rect 44706 43598 44718 43650
rect 44770 43598 44782 43650
rect 40350 43586 40402 43598
rect 45054 43586 45106 43598
rect 47294 43650 47346 43662
rect 47294 43586 47346 43598
rect 47518 43650 47570 43662
rect 47518 43586 47570 43598
rect 48078 43650 48130 43662
rect 54350 43650 54402 43662
rect 49746 43598 49758 43650
rect 49810 43598 49822 43650
rect 50306 43598 50318 43650
rect 50370 43598 50382 43650
rect 51650 43598 51662 43650
rect 51714 43598 51726 43650
rect 51986 43598 51998 43650
rect 52050 43598 52062 43650
rect 48078 43586 48130 43598
rect 54350 43586 54402 43598
rect 2830 43538 2882 43550
rect 6974 43538 7026 43550
rect 10222 43538 10274 43550
rect 11118 43538 11170 43550
rect 3154 43486 3166 43538
rect 3218 43486 3230 43538
rect 8418 43486 8430 43538
rect 8482 43486 8494 43538
rect 10882 43486 10894 43538
rect 10946 43486 10958 43538
rect 2830 43474 2882 43486
rect 6974 43474 7026 43486
rect 10222 43474 10274 43486
rect 11118 43474 11170 43486
rect 11902 43538 11954 43550
rect 15038 43538 15090 43550
rect 12562 43486 12574 43538
rect 12626 43486 12638 43538
rect 11902 43474 11954 43486
rect 15038 43474 15090 43486
rect 15486 43538 15538 43550
rect 15486 43474 15538 43486
rect 16270 43538 16322 43550
rect 18286 43538 18338 43550
rect 16594 43486 16606 43538
rect 16658 43486 16670 43538
rect 16270 43474 16322 43486
rect 18286 43474 18338 43486
rect 19070 43538 19122 43550
rect 19070 43474 19122 43486
rect 20302 43538 20354 43550
rect 20302 43474 20354 43486
rect 21422 43538 21474 43550
rect 21422 43474 21474 43486
rect 23102 43538 23154 43550
rect 23102 43474 23154 43486
rect 25678 43538 25730 43550
rect 35870 43538 35922 43550
rect 40014 43538 40066 43550
rect 42478 43538 42530 43550
rect 45278 43538 45330 43550
rect 29586 43486 29598 43538
rect 29650 43486 29662 43538
rect 31266 43486 31278 43538
rect 31330 43486 31342 43538
rect 31714 43486 31726 43538
rect 31778 43486 31790 43538
rect 36418 43486 36430 43538
rect 36482 43486 36494 43538
rect 40786 43486 40798 43538
rect 40850 43486 40862 43538
rect 41682 43486 41694 43538
rect 41746 43486 41758 43538
rect 42802 43486 42814 43538
rect 42866 43486 42878 43538
rect 44818 43486 44830 43538
rect 44882 43486 44894 43538
rect 25678 43474 25730 43486
rect 35870 43474 35922 43486
rect 40014 43474 40066 43486
rect 42478 43474 42530 43486
rect 45278 43474 45330 43486
rect 45838 43538 45890 43550
rect 45838 43474 45890 43486
rect 46174 43538 46226 43550
rect 48526 43538 48578 43550
rect 46610 43486 46622 43538
rect 46674 43486 46686 43538
rect 46174 43474 46226 43486
rect 48526 43474 48578 43486
rect 49646 43538 49698 43550
rect 49646 43474 49698 43486
rect 51326 43538 51378 43550
rect 57374 43538 57426 43550
rect 53890 43486 53902 43538
rect 53954 43486 53966 43538
rect 54114 43486 54126 43538
rect 54178 43486 54190 43538
rect 56130 43486 56142 43538
rect 56194 43486 56206 43538
rect 51326 43474 51378 43486
rect 57374 43474 57426 43486
rect 7646 43426 7698 43438
rect 7646 43362 7698 43374
rect 9662 43426 9714 43438
rect 9662 43362 9714 43374
rect 22318 43426 22370 43438
rect 32846 43426 32898 43438
rect 29026 43374 29038 43426
rect 29090 43374 29102 43426
rect 22318 43362 22370 43374
rect 32846 43362 32898 43374
rect 35086 43426 35138 43438
rect 35086 43362 35138 43374
rect 35422 43426 35474 43438
rect 43710 43426 43762 43438
rect 49422 43426 49474 43438
rect 40226 43374 40238 43426
rect 40290 43374 40302 43426
rect 44930 43374 44942 43426
rect 44994 43374 45006 43426
rect 47618 43374 47630 43426
rect 47682 43374 47694 43426
rect 35422 43362 35474 43374
rect 43710 43362 43762 43374
rect 49422 43362 49474 43374
rect 52110 43426 52162 43438
rect 52110 43362 52162 43374
rect 52782 43426 52834 43438
rect 52782 43362 52834 43374
rect 53230 43426 53282 43438
rect 56590 43426 56642 43438
rect 55346 43374 55358 43426
rect 55410 43374 55422 43426
rect 53230 43362 53282 43374
rect 56590 43362 56642 43374
rect 57934 43426 57986 43438
rect 57934 43362 57986 43374
rect 12126 43314 12178 43326
rect 12126 43250 12178 43262
rect 12350 43314 12402 43326
rect 12350 43250 12402 43262
rect 14142 43314 14194 43326
rect 14142 43250 14194 43262
rect 15262 43314 15314 43326
rect 15262 43250 15314 43262
rect 20078 43314 20130 43326
rect 20078 43250 20130 43262
rect 20638 43314 20690 43326
rect 20638 43250 20690 43262
rect 20862 43314 20914 43326
rect 46286 43314 46338 43326
rect 43138 43262 43150 43314
rect 43202 43262 43214 43314
rect 20862 43250 20914 43262
rect 46286 43250 46338 43262
rect 51102 43314 51154 43326
rect 54462 43314 54514 43326
rect 52434 43262 52446 43314
rect 52498 43311 52510 43314
rect 52658 43311 52670 43314
rect 52498 43265 52670 43311
rect 52498 43262 52510 43265
rect 52658 43262 52670 43265
rect 52722 43262 52734 43314
rect 51102 43250 51154 43262
rect 54462 43250 54514 43262
rect 1344 43146 58576 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 58576 43146
rect 1344 43060 58576 43094
rect 4958 42978 5010 42990
rect 4958 42914 5010 42926
rect 6414 42978 6466 42990
rect 6414 42914 6466 42926
rect 11342 42978 11394 42990
rect 20302 42978 20354 42990
rect 31054 42978 31106 42990
rect 11890 42926 11902 42978
rect 11954 42975 11966 42978
rect 12450 42975 12462 42978
rect 11954 42929 12462 42975
rect 11954 42926 11966 42929
rect 12450 42926 12462 42929
rect 12514 42926 12526 42978
rect 22978 42926 22990 42978
rect 23042 42926 23054 42978
rect 29810 42926 29822 42978
rect 29874 42926 29886 42978
rect 11342 42914 11394 42926
rect 20302 42914 20354 42926
rect 31054 42914 31106 42926
rect 38446 42978 38498 42990
rect 38446 42914 38498 42926
rect 39454 42978 39506 42990
rect 39454 42914 39506 42926
rect 40238 42978 40290 42990
rect 45726 42978 45778 42990
rect 43474 42926 43486 42978
rect 43538 42926 43550 42978
rect 40238 42914 40290 42926
rect 45726 42914 45778 42926
rect 46286 42978 46338 42990
rect 54014 42978 54066 42990
rect 47058 42926 47070 42978
rect 47122 42975 47134 42978
rect 47122 42929 47679 42975
rect 47122 42926 47134 42929
rect 46286 42914 46338 42926
rect 3054 42866 3106 42878
rect 3054 42802 3106 42814
rect 5742 42866 5794 42878
rect 12014 42866 12066 42878
rect 7186 42814 7198 42866
rect 7250 42814 7262 42866
rect 5742 42802 5794 42814
rect 12014 42802 12066 42814
rect 12462 42866 12514 42878
rect 12462 42802 12514 42814
rect 13806 42866 13858 42878
rect 13806 42802 13858 42814
rect 15374 42866 15426 42878
rect 15374 42802 15426 42814
rect 18846 42866 18898 42878
rect 26350 42866 26402 42878
rect 31950 42866 32002 42878
rect 23314 42814 23326 42866
rect 23378 42814 23390 42866
rect 24322 42814 24334 42866
rect 24386 42814 24398 42866
rect 28354 42814 28366 42866
rect 28418 42814 28430 42866
rect 18846 42802 18898 42814
rect 26350 42802 26402 42814
rect 31950 42802 32002 42814
rect 33966 42866 34018 42878
rect 33966 42802 34018 42814
rect 36094 42866 36146 42878
rect 36094 42802 36146 42814
rect 36654 42866 36706 42878
rect 41806 42866 41858 42878
rect 40002 42814 40014 42866
rect 40066 42814 40078 42866
rect 36654 42802 36706 42814
rect 41806 42802 41858 42814
rect 47070 42866 47122 42878
rect 47633 42863 47679 42929
rect 47730 42926 47742 42978
rect 47794 42975 47806 42978
rect 49298 42975 49310 42978
rect 47794 42929 49310 42975
rect 47794 42926 47806 42929
rect 49298 42926 49310 42929
rect 49362 42926 49374 42978
rect 57138 42926 57150 42978
rect 57202 42975 57214 42978
rect 57698 42975 57710 42978
rect 57202 42929 57710 42975
rect 57202 42926 57214 42929
rect 57698 42926 57710 42929
rect 57762 42926 57774 42978
rect 54014 42914 54066 42926
rect 48414 42866 48466 42878
rect 47842 42863 47854 42866
rect 47633 42817 47854 42863
rect 47842 42814 47854 42817
rect 47906 42814 47918 42866
rect 47070 42802 47122 42814
rect 48414 42802 48466 42814
rect 49310 42866 49362 42878
rect 49310 42802 49362 42814
rect 50094 42866 50146 42878
rect 50094 42802 50146 42814
rect 53342 42866 53394 42878
rect 53342 42802 53394 42814
rect 57710 42866 57762 42878
rect 57710 42802 57762 42814
rect 6302 42754 6354 42766
rect 11006 42754 11058 42766
rect 7298 42702 7310 42754
rect 7362 42702 7374 42754
rect 6302 42690 6354 42702
rect 11006 42690 11058 42702
rect 11118 42754 11170 42766
rect 11118 42690 11170 42702
rect 13582 42754 13634 42766
rect 13582 42690 13634 42702
rect 15822 42754 15874 42766
rect 26910 42754 26962 42766
rect 30382 42754 30434 42766
rect 31502 42754 31554 42766
rect 19506 42702 19518 42754
rect 19570 42702 19582 42754
rect 20514 42702 20526 42754
rect 20578 42751 20590 42754
rect 20738 42751 20750 42754
rect 20578 42705 20750 42751
rect 20578 42702 20590 42705
rect 20738 42702 20750 42705
rect 20802 42702 20814 42754
rect 22866 42702 22878 42754
rect 22930 42702 22942 42754
rect 28130 42702 28142 42754
rect 28194 42702 28206 42754
rect 30594 42702 30606 42754
rect 30658 42702 30670 42754
rect 15822 42690 15874 42702
rect 26910 42690 26962 42702
rect 30382 42690 30434 42702
rect 31502 42690 31554 42702
rect 31726 42754 31778 42766
rect 31726 42690 31778 42702
rect 32510 42754 32562 42766
rect 32510 42690 32562 42702
rect 32734 42754 32786 42766
rect 32734 42690 32786 42702
rect 37662 42754 37714 42766
rect 37662 42690 37714 42702
rect 37886 42754 37938 42766
rect 37886 42690 37938 42702
rect 39678 42754 39730 42766
rect 39678 42690 39730 42702
rect 40686 42754 40738 42766
rect 40686 42690 40738 42702
rect 42814 42754 42866 42766
rect 42814 42690 42866 42702
rect 43038 42754 43090 42766
rect 45950 42754 46002 42766
rect 44258 42702 44270 42754
rect 44322 42702 44334 42754
rect 43038 42690 43090 42702
rect 45950 42690 46002 42702
rect 46510 42754 46562 42766
rect 52558 42754 52610 42766
rect 50306 42702 50318 42754
rect 50370 42702 50382 42754
rect 50866 42702 50878 42754
rect 50930 42702 50942 42754
rect 51538 42702 51550 42754
rect 51602 42702 51614 42754
rect 46510 42690 46562 42702
rect 52558 42690 52610 42702
rect 54574 42754 54626 42766
rect 54574 42690 54626 42702
rect 55022 42754 55074 42766
rect 55022 42690 55074 42702
rect 55918 42754 55970 42766
rect 56242 42702 56254 42754
rect 56306 42702 56318 42754
rect 55918 42690 55970 42702
rect 2942 42642 2994 42654
rect 2942 42578 2994 42590
rect 3278 42642 3330 42654
rect 3278 42578 3330 42590
rect 3502 42642 3554 42654
rect 3502 42578 3554 42590
rect 4846 42642 4898 42654
rect 14142 42642 14194 42654
rect 6962 42590 6974 42642
rect 7026 42590 7038 42642
rect 4846 42578 4898 42590
rect 14142 42578 14194 42590
rect 15262 42642 15314 42654
rect 15262 42578 15314 42590
rect 15598 42642 15650 42654
rect 15598 42578 15650 42590
rect 20414 42642 20466 42654
rect 20414 42578 20466 42590
rect 20862 42642 20914 42654
rect 20862 42578 20914 42590
rect 24110 42642 24162 42654
rect 24110 42578 24162 42590
rect 28814 42642 28866 42654
rect 28814 42578 28866 42590
rect 30270 42642 30322 42654
rect 30270 42578 30322 42590
rect 32622 42642 32674 42654
rect 32622 42578 32674 42590
rect 35646 42642 35698 42654
rect 35646 42578 35698 42590
rect 38222 42642 38274 42654
rect 38222 42578 38274 42590
rect 40014 42642 40066 42654
rect 40014 42578 40066 42590
rect 42926 42642 42978 42654
rect 46062 42642 46114 42654
rect 54014 42642 54066 42654
rect 44034 42590 44046 42642
rect 44098 42590 44110 42642
rect 50418 42590 50430 42642
rect 50482 42590 50494 42642
rect 52210 42590 52222 42642
rect 52274 42590 52286 42642
rect 42926 42578 42978 42590
rect 46062 42578 46114 42590
rect 54014 42578 54066 42590
rect 54126 42642 54178 42654
rect 54126 42578 54178 42590
rect 55806 42642 55858 42654
rect 55806 42578 55858 42590
rect 6750 42530 6802 42542
rect 6750 42466 6802 42478
rect 7758 42530 7810 42542
rect 7758 42466 7810 42478
rect 11006 42530 11058 42542
rect 11006 42466 11058 42478
rect 13022 42530 13074 42542
rect 13022 42466 13074 42478
rect 13918 42530 13970 42542
rect 13918 42466 13970 42478
rect 14702 42530 14754 42542
rect 14702 42466 14754 42478
rect 16270 42530 16322 42542
rect 16270 42466 16322 42478
rect 17054 42530 17106 42542
rect 17054 42466 17106 42478
rect 17614 42530 17666 42542
rect 17614 42466 17666 42478
rect 18062 42530 18114 42542
rect 18062 42466 18114 42478
rect 19742 42530 19794 42542
rect 19742 42466 19794 42478
rect 24334 42530 24386 42542
rect 24334 42466 24386 42478
rect 27246 42530 27298 42542
rect 27246 42466 27298 42478
rect 32958 42530 33010 42542
rect 32958 42466 33010 42478
rect 33518 42530 33570 42542
rect 33518 42466 33570 42478
rect 34750 42530 34802 42542
rect 34750 42466 34802 42478
rect 35422 42530 35474 42542
rect 35422 42466 35474 42478
rect 35534 42530 35586 42542
rect 35534 42466 35586 42478
rect 37550 42530 37602 42542
rect 37550 42466 37602 42478
rect 41134 42530 41186 42542
rect 41134 42466 41186 42478
rect 41246 42530 41298 42542
rect 41246 42466 41298 42478
rect 41358 42530 41410 42542
rect 41358 42466 41410 42478
rect 47518 42530 47570 42542
rect 47518 42466 47570 42478
rect 48078 42530 48130 42542
rect 48078 42466 48130 42478
rect 48974 42530 49026 42542
rect 48974 42466 49026 42478
rect 55134 42530 55186 42542
rect 55134 42466 55186 42478
rect 55246 42530 55298 42542
rect 55246 42466 55298 42478
rect 57374 42530 57426 42542
rect 57374 42466 57426 42478
rect 1344 42362 58576 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 58576 42362
rect 1344 42276 58576 42310
rect 14030 42194 14082 42206
rect 14030 42130 14082 42142
rect 15710 42194 15762 42206
rect 15710 42130 15762 42142
rect 19966 42194 20018 42206
rect 19966 42130 20018 42142
rect 20190 42194 20242 42206
rect 20190 42130 20242 42142
rect 20750 42194 20802 42206
rect 20750 42130 20802 42142
rect 21310 42194 21362 42206
rect 21310 42130 21362 42142
rect 26014 42194 26066 42206
rect 26014 42130 26066 42142
rect 35870 42194 35922 42206
rect 35870 42130 35922 42142
rect 36094 42194 36146 42206
rect 36094 42130 36146 42142
rect 36990 42194 37042 42206
rect 36990 42130 37042 42142
rect 37998 42194 38050 42206
rect 37998 42130 38050 42142
rect 38894 42194 38946 42206
rect 38894 42130 38946 42142
rect 40238 42194 40290 42206
rect 40238 42130 40290 42142
rect 45278 42194 45330 42206
rect 52446 42194 52498 42206
rect 52098 42142 52110 42194
rect 52162 42142 52174 42194
rect 45278 42130 45330 42142
rect 52446 42130 52498 42142
rect 53118 42194 53170 42206
rect 53118 42130 53170 42142
rect 56366 42194 56418 42206
rect 56366 42130 56418 42142
rect 1822 42082 1874 42094
rect 5518 42082 5570 42094
rect 3714 42030 3726 42082
rect 3778 42030 3790 42082
rect 1822 42018 1874 42030
rect 5518 42018 5570 42030
rect 6750 42082 6802 42094
rect 6750 42018 6802 42030
rect 6974 42082 7026 42094
rect 6974 42018 7026 42030
rect 12350 42082 12402 42094
rect 12350 42018 12402 42030
rect 13918 42082 13970 42094
rect 32398 42082 32450 42094
rect 16594 42030 16606 42082
rect 16658 42030 16670 42082
rect 13918 42018 13970 42030
rect 32398 42018 32450 42030
rect 34078 42082 34130 42094
rect 34078 42018 34130 42030
rect 36766 42082 36818 42094
rect 36766 42018 36818 42030
rect 37326 42082 37378 42094
rect 37326 42018 37378 42030
rect 38110 42082 38162 42094
rect 38110 42018 38162 42030
rect 39342 42082 39394 42094
rect 39342 42018 39394 42030
rect 40462 42082 40514 42094
rect 55470 42082 55522 42094
rect 44818 42030 44830 42082
rect 44882 42030 44894 42082
rect 47618 42030 47630 42082
rect 47682 42030 47694 42082
rect 40462 42018 40514 42030
rect 55470 42018 55522 42030
rect 56142 42082 56194 42094
rect 56142 42018 56194 42030
rect 5406 41970 5458 41982
rect 2482 41918 2494 41970
rect 2546 41918 2558 41970
rect 5406 41906 5458 41918
rect 5742 41970 5794 41982
rect 5742 41906 5794 41918
rect 5966 41970 6018 41982
rect 5966 41906 6018 41918
rect 6414 41970 6466 41982
rect 9998 41970 10050 41982
rect 14254 41970 14306 41982
rect 9762 41918 9774 41970
rect 9826 41918 9838 41970
rect 12898 41918 12910 41970
rect 12962 41918 12974 41970
rect 6414 41906 6466 41918
rect 9998 41906 10050 41918
rect 14254 41906 14306 41918
rect 14478 41970 14530 41982
rect 18062 41970 18114 41982
rect 16706 41918 16718 41970
rect 16770 41918 16782 41970
rect 14478 41906 14530 41918
rect 18062 41906 18114 41918
rect 18958 41970 19010 41982
rect 18958 41906 19010 41918
rect 19854 41970 19906 41982
rect 19854 41906 19906 41918
rect 20638 41970 20690 41982
rect 20638 41906 20690 41918
rect 25790 41970 25842 41982
rect 25790 41906 25842 41918
rect 26014 41970 26066 41982
rect 26014 41906 26066 41918
rect 26350 41970 26402 41982
rect 26350 41906 26402 41918
rect 26686 41970 26738 41982
rect 33630 41970 33682 41982
rect 35646 41970 35698 41982
rect 31826 41918 31838 41970
rect 31890 41918 31902 41970
rect 34738 41918 34750 41970
rect 34802 41918 34814 41970
rect 26686 41906 26738 41918
rect 33630 41906 33682 41918
rect 35646 41906 35698 41918
rect 37102 41970 37154 41982
rect 37102 41906 37154 41918
rect 37774 41970 37826 41982
rect 37774 41906 37826 41918
rect 38670 41970 38722 41982
rect 38670 41906 38722 41918
rect 39118 41970 39170 41982
rect 39118 41906 39170 41918
rect 39902 41970 39954 41982
rect 39902 41906 39954 41918
rect 40126 41970 40178 41982
rect 45950 41970 46002 41982
rect 41794 41918 41806 41970
rect 41858 41918 41870 41970
rect 42018 41918 42030 41970
rect 42082 41918 42094 41970
rect 43810 41918 43822 41970
rect 43874 41918 43886 41970
rect 40126 41906 40178 41918
rect 45950 41906 46002 41918
rect 46622 41970 46674 41982
rect 46622 41906 46674 41918
rect 46846 41970 46898 41982
rect 50206 41970 50258 41982
rect 51102 41970 51154 41982
rect 48178 41918 48190 41970
rect 48242 41918 48254 41970
rect 48514 41918 48526 41970
rect 48578 41918 48590 41970
rect 50418 41918 50430 41970
rect 50482 41918 50494 41970
rect 46846 41906 46898 41918
rect 50206 41906 50258 41918
rect 51102 41906 51154 41918
rect 55246 41970 55298 41982
rect 56690 41918 56702 41970
rect 56754 41918 56766 41970
rect 55246 41906 55298 41918
rect 3838 41858 3890 41870
rect 8766 41858 8818 41870
rect 6850 41806 6862 41858
rect 6914 41806 6926 41858
rect 3838 41794 3890 41806
rect 8766 41794 8818 41806
rect 10782 41858 10834 41870
rect 10782 41794 10834 41806
rect 11342 41858 11394 41870
rect 14926 41858 14978 41870
rect 13122 41806 13134 41858
rect 13186 41806 13198 41858
rect 11342 41794 11394 41806
rect 14926 41794 14978 41806
rect 17726 41858 17778 41870
rect 17726 41794 17778 41806
rect 18622 41858 18674 41870
rect 35758 41858 35810 41870
rect 51550 41858 51602 41870
rect 31602 41806 31614 41858
rect 31666 41806 31678 41858
rect 34962 41806 34974 41858
rect 35026 41806 35038 41858
rect 47730 41806 47742 41858
rect 47794 41806 47806 41858
rect 49858 41806 49870 41858
rect 49922 41806 49934 41858
rect 18622 41794 18674 41806
rect 35758 41794 35810 41806
rect 51550 41794 51602 41806
rect 53678 41858 53730 41870
rect 53678 41794 53730 41806
rect 54126 41858 54178 41870
rect 54126 41794 54178 41806
rect 54574 41858 54626 41870
rect 56254 41858 56306 41870
rect 55570 41806 55582 41858
rect 55634 41806 55646 41858
rect 54574 41794 54626 41806
rect 56254 41794 56306 41806
rect 57374 41858 57426 41870
rect 57374 41794 57426 41806
rect 57822 41858 57874 41870
rect 57822 41794 57874 41806
rect 10110 41746 10162 41758
rect 10110 41682 10162 41694
rect 16046 41746 16098 41758
rect 20750 41746 20802 41758
rect 17714 41694 17726 41746
rect 17778 41743 17790 41746
rect 18610 41743 18622 41746
rect 17778 41697 18622 41743
rect 17778 41694 17790 41697
rect 18610 41694 18622 41697
rect 18674 41694 18686 41746
rect 16046 41682 16098 41694
rect 20750 41682 20802 41694
rect 39230 41746 39282 41758
rect 39230 41682 39282 41694
rect 46398 41746 46450 41758
rect 54114 41694 54126 41746
rect 54178 41743 54190 41746
rect 55010 41743 55022 41746
rect 54178 41697 55022 41743
rect 54178 41694 54190 41697
rect 55010 41694 55022 41697
rect 55074 41694 55086 41746
rect 46398 41682 46450 41694
rect 1344 41578 58576 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 58576 41578
rect 1344 41492 58576 41526
rect 3950 41410 4002 41422
rect 3950 41346 4002 41358
rect 7870 41410 7922 41422
rect 13918 41410 13970 41422
rect 23102 41410 23154 41422
rect 8978 41358 8990 41410
rect 9042 41358 9054 41410
rect 14242 41358 14254 41410
rect 14306 41358 14318 41410
rect 16146 41358 16158 41410
rect 16210 41358 16222 41410
rect 7870 41346 7922 41358
rect 13918 41346 13970 41358
rect 23102 41346 23154 41358
rect 27246 41410 27298 41422
rect 27246 41346 27298 41358
rect 49310 41410 49362 41422
rect 51314 41358 51326 41410
rect 51378 41407 51390 41410
rect 51538 41407 51550 41410
rect 51378 41361 51550 41407
rect 51378 41358 51390 41361
rect 51538 41358 51550 41361
rect 51602 41358 51614 41410
rect 49310 41346 49362 41358
rect 10446 41298 10498 41310
rect 3714 41246 3726 41298
rect 3778 41246 3790 41298
rect 10446 41234 10498 41246
rect 13694 41298 13746 41310
rect 18286 41298 18338 41310
rect 17826 41246 17838 41298
rect 17890 41246 17902 41298
rect 13694 41234 13746 41246
rect 18286 41234 18338 41246
rect 26350 41298 26402 41310
rect 26350 41234 26402 41246
rect 35646 41298 35698 41310
rect 35646 41234 35698 41246
rect 37886 41298 37938 41310
rect 40574 41298 40626 41310
rect 39106 41246 39118 41298
rect 39170 41246 39182 41298
rect 37886 41234 37938 41246
rect 40574 41234 40626 41246
rect 41022 41298 41074 41310
rect 41022 41234 41074 41246
rect 42142 41298 42194 41310
rect 42142 41234 42194 41246
rect 51326 41298 51378 41310
rect 51326 41234 51378 41246
rect 2942 41186 2994 41198
rect 8542 41186 8594 41198
rect 2594 41134 2606 41186
rect 2658 41134 2670 41186
rect 6514 41134 6526 41186
rect 6578 41134 6590 41186
rect 2942 41122 2994 41134
rect 8542 41122 8594 41134
rect 9438 41186 9490 41198
rect 9438 41122 9490 41134
rect 10222 41186 10274 41198
rect 10222 41122 10274 41134
rect 10782 41186 10834 41198
rect 10782 41122 10834 41134
rect 15822 41186 15874 41198
rect 19294 41186 19346 41198
rect 16482 41134 16494 41186
rect 16546 41134 16558 41186
rect 17602 41134 17614 41186
rect 17666 41134 17678 41186
rect 15822 41122 15874 41134
rect 19294 41122 19346 41134
rect 21870 41186 21922 41198
rect 27806 41186 27858 41198
rect 24994 41134 25006 41186
rect 25058 41134 25070 41186
rect 21870 41122 21922 41134
rect 27806 41122 27858 41134
rect 28590 41186 28642 41198
rect 28590 41122 28642 41134
rect 29598 41186 29650 41198
rect 29598 41122 29650 41134
rect 34190 41186 34242 41198
rect 34190 41122 34242 41134
rect 34302 41186 34354 41198
rect 46510 41186 46562 41198
rect 56590 41186 56642 41198
rect 35410 41134 35422 41186
rect 35474 41134 35486 41186
rect 36306 41134 36318 41186
rect 36370 41134 36382 41186
rect 38658 41134 38670 41186
rect 38722 41134 38734 41186
rect 38882 41134 38894 41186
rect 38946 41134 38958 41186
rect 42242 41134 42254 41186
rect 42306 41134 42318 41186
rect 42690 41134 42702 41186
rect 42754 41134 42766 41186
rect 43586 41134 43598 41186
rect 43650 41134 43662 41186
rect 54114 41134 54126 41186
rect 54178 41134 54190 41186
rect 55234 41134 55246 41186
rect 55298 41134 55310 41186
rect 34302 41122 34354 41134
rect 46510 41122 46562 41134
rect 56590 41122 56642 41134
rect 3054 41074 3106 41086
rect 3054 41010 3106 41022
rect 3726 41074 3778 41086
rect 6190 41074 6242 41086
rect 5730 41022 5742 41074
rect 5794 41022 5806 41074
rect 3726 41010 3778 41022
rect 6190 41010 6242 41022
rect 6302 41074 6354 41086
rect 6302 41010 6354 41022
rect 8206 41074 8258 41086
rect 8206 41010 8258 41022
rect 9550 41074 9602 41086
rect 9550 41010 9602 41022
rect 9662 41074 9714 41086
rect 9662 41010 9714 41022
rect 10670 41074 10722 41086
rect 10670 41010 10722 41022
rect 21646 41074 21698 41086
rect 21646 41010 21698 41022
rect 22766 41074 22818 41086
rect 27358 41074 27410 41086
rect 25890 41022 25902 41074
rect 25954 41022 25966 41074
rect 22766 41010 22818 41022
rect 27358 41010 27410 41022
rect 28702 41074 28754 41086
rect 28702 41010 28754 41022
rect 29934 41074 29986 41086
rect 29934 41010 29986 41022
rect 30158 41074 30210 41086
rect 30158 41010 30210 41022
rect 31502 41074 31554 41086
rect 31502 41010 31554 41022
rect 31726 41074 31778 41086
rect 31726 41010 31778 41022
rect 31838 41074 31890 41086
rect 31838 41010 31890 41022
rect 33854 41074 33906 41086
rect 39118 41074 39170 41086
rect 35634 41022 35646 41074
rect 35698 41022 35710 41074
rect 36082 41022 36094 41074
rect 36146 41022 36158 41074
rect 33854 41010 33906 41022
rect 39118 41010 39170 41022
rect 39678 41074 39730 41086
rect 39678 41010 39730 41022
rect 40014 41074 40066 41086
rect 45390 41074 45442 41086
rect 44370 41022 44382 41074
rect 44434 41022 44446 41074
rect 40014 41010 40066 41022
rect 45390 41010 45442 41022
rect 46286 41074 46338 41086
rect 46286 41010 46338 41022
rect 46846 41074 46898 41086
rect 46846 41010 46898 41022
rect 47742 41074 47794 41086
rect 47742 41010 47794 41022
rect 48974 41074 49026 41086
rect 48974 41010 49026 41022
rect 49198 41074 49250 41086
rect 56254 41074 56306 41086
rect 53778 41022 53790 41074
rect 53842 41022 53854 41074
rect 49198 41010 49250 41022
rect 56254 41010 56306 41022
rect 7310 40962 7362 40974
rect 7310 40898 7362 40910
rect 7982 40962 8034 40974
rect 7982 40898 8034 40910
rect 11678 40962 11730 40974
rect 11678 40898 11730 40910
rect 12574 40962 12626 40974
rect 12574 40898 12626 40910
rect 13022 40962 13074 40974
rect 13022 40898 13074 40910
rect 15150 40962 15202 40974
rect 15150 40898 15202 40910
rect 18846 40962 18898 40974
rect 18846 40898 18898 40910
rect 19630 40962 19682 40974
rect 19630 40898 19682 40910
rect 20190 40962 20242 40974
rect 20190 40898 20242 40910
rect 20862 40962 20914 40974
rect 22990 40962 23042 40974
rect 27246 40962 27298 40974
rect 22194 40910 22206 40962
rect 22258 40910 22270 40962
rect 24658 40910 24670 40962
rect 24722 40910 24734 40962
rect 20862 40898 20914 40910
rect 22990 40898 23042 40910
rect 27246 40898 27298 40910
rect 28926 40962 28978 40974
rect 28926 40898 28978 40910
rect 29822 40962 29874 40974
rect 29822 40898 29874 40910
rect 34078 40962 34130 40974
rect 34078 40898 34130 40910
rect 37550 40962 37602 40974
rect 37550 40898 37602 40910
rect 41582 40962 41634 40974
rect 41582 40898 41634 40910
rect 43822 40962 43874 40974
rect 43822 40898 43874 40910
rect 44718 40962 44770 40974
rect 44718 40898 44770 40910
rect 46398 40962 46450 40974
rect 49758 40962 49810 40974
rect 48066 40910 48078 40962
rect 48130 40910 48142 40962
rect 46398 40898 46450 40910
rect 49758 40898 49810 40910
rect 50206 40962 50258 40974
rect 50206 40898 50258 40910
rect 50654 40962 50706 40974
rect 50654 40898 50706 40910
rect 51774 40962 51826 40974
rect 51774 40898 51826 40910
rect 52222 40962 52274 40974
rect 52222 40898 52274 40910
rect 52782 40962 52834 40974
rect 56366 40962 56418 40974
rect 55346 40910 55358 40962
rect 55410 40910 55422 40962
rect 52782 40898 52834 40910
rect 56366 40898 56418 40910
rect 57038 40962 57090 40974
rect 57038 40898 57090 40910
rect 57374 40962 57426 40974
rect 57374 40898 57426 40910
rect 57822 40962 57874 40974
rect 57822 40898 57874 40910
rect 1344 40794 58576 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 58576 40794
rect 1344 40708 58576 40742
rect 4958 40626 5010 40638
rect 4958 40562 5010 40574
rect 6302 40626 6354 40638
rect 6302 40562 6354 40574
rect 6750 40626 6802 40638
rect 6750 40562 6802 40574
rect 9886 40626 9938 40638
rect 9886 40562 9938 40574
rect 9998 40626 10050 40638
rect 9998 40562 10050 40574
rect 13246 40626 13298 40638
rect 13246 40562 13298 40574
rect 19518 40626 19570 40638
rect 19518 40562 19570 40574
rect 20638 40626 20690 40638
rect 20638 40562 20690 40574
rect 25790 40626 25842 40638
rect 36206 40626 36258 40638
rect 34738 40574 34750 40626
rect 34802 40574 34814 40626
rect 25790 40562 25842 40574
rect 36206 40562 36258 40574
rect 36318 40626 36370 40638
rect 36318 40562 36370 40574
rect 36430 40626 36482 40638
rect 36430 40562 36482 40574
rect 36878 40626 36930 40638
rect 36878 40562 36930 40574
rect 39118 40626 39170 40638
rect 39118 40562 39170 40574
rect 39566 40626 39618 40638
rect 39566 40562 39618 40574
rect 40462 40626 40514 40638
rect 40462 40562 40514 40574
rect 41694 40626 41746 40638
rect 41694 40562 41746 40574
rect 43038 40626 43090 40638
rect 43038 40562 43090 40574
rect 43262 40626 43314 40638
rect 43262 40562 43314 40574
rect 44606 40626 44658 40638
rect 44606 40562 44658 40574
rect 44718 40626 44770 40638
rect 44718 40562 44770 40574
rect 45166 40626 45218 40638
rect 45166 40562 45218 40574
rect 45614 40626 45666 40638
rect 45614 40562 45666 40574
rect 48526 40626 48578 40638
rect 48526 40562 48578 40574
rect 48638 40626 48690 40638
rect 48638 40562 48690 40574
rect 48750 40626 48802 40638
rect 48750 40562 48802 40574
rect 51214 40626 51266 40638
rect 51874 40574 51886 40626
rect 51938 40574 51950 40626
rect 54338 40574 54350 40626
rect 54402 40574 54414 40626
rect 51214 40562 51266 40574
rect 7534 40514 7586 40526
rect 7534 40450 7586 40462
rect 7646 40514 7698 40526
rect 7646 40450 7698 40462
rect 10222 40514 10274 40526
rect 10222 40450 10274 40462
rect 14478 40514 14530 40526
rect 19406 40514 19458 40526
rect 16370 40462 16382 40514
rect 16434 40462 16446 40514
rect 14478 40450 14530 40462
rect 19406 40450 19458 40462
rect 20526 40514 20578 40526
rect 20526 40450 20578 40462
rect 21646 40514 21698 40526
rect 21646 40450 21698 40462
rect 23886 40514 23938 40526
rect 23886 40450 23938 40462
rect 26798 40514 26850 40526
rect 26798 40450 26850 40462
rect 33742 40514 33794 40526
rect 33742 40450 33794 40462
rect 33854 40514 33906 40526
rect 33854 40450 33906 40462
rect 38222 40514 38274 40526
rect 38222 40450 38274 40462
rect 41918 40514 41970 40526
rect 41918 40450 41970 40462
rect 42142 40514 42194 40526
rect 42142 40450 42194 40462
rect 44494 40514 44546 40526
rect 48302 40514 48354 40526
rect 46946 40462 46958 40514
rect 47010 40462 47022 40514
rect 44494 40450 44546 40462
rect 48302 40450 48354 40462
rect 49534 40514 49586 40526
rect 49534 40450 49586 40462
rect 49870 40514 49922 40526
rect 49870 40450 49922 40462
rect 52334 40514 52386 40526
rect 52334 40450 52386 40462
rect 52558 40514 52610 40526
rect 52558 40450 52610 40462
rect 55134 40514 55186 40526
rect 55134 40450 55186 40462
rect 8094 40402 8146 40414
rect 2818 40350 2830 40402
rect 2882 40350 2894 40402
rect 8094 40338 8146 40350
rect 9774 40402 9826 40414
rect 9774 40338 9826 40350
rect 11566 40402 11618 40414
rect 11566 40338 11618 40350
rect 12126 40402 12178 40414
rect 12126 40338 12178 40350
rect 15374 40402 15426 40414
rect 15374 40338 15426 40350
rect 16046 40402 16098 40414
rect 16046 40338 16098 40350
rect 16942 40402 16994 40414
rect 16942 40338 16994 40350
rect 17726 40402 17778 40414
rect 17726 40338 17778 40350
rect 18734 40402 18786 40414
rect 18734 40338 18786 40350
rect 19294 40402 19346 40414
rect 19294 40338 19346 40350
rect 19742 40402 19794 40414
rect 19742 40338 19794 40350
rect 20302 40402 20354 40414
rect 20302 40338 20354 40350
rect 20974 40402 21026 40414
rect 20974 40338 21026 40350
rect 21534 40402 21586 40414
rect 21534 40338 21586 40350
rect 23326 40402 23378 40414
rect 28366 40402 28418 40414
rect 30046 40402 30098 40414
rect 24322 40350 24334 40402
rect 24386 40350 24398 40402
rect 27458 40350 27470 40402
rect 27522 40350 27534 40402
rect 28914 40350 28926 40402
rect 28978 40350 28990 40402
rect 23326 40338 23378 40350
rect 28366 40338 28418 40350
rect 30046 40338 30098 40350
rect 30494 40402 30546 40414
rect 33518 40402 33570 40414
rect 31378 40350 31390 40402
rect 31442 40350 31454 40402
rect 30494 40338 30546 40350
rect 33518 40338 33570 40350
rect 35310 40402 35362 40414
rect 35310 40338 35362 40350
rect 35758 40402 35810 40414
rect 35758 40338 35810 40350
rect 37998 40402 38050 40414
rect 37998 40338 38050 40350
rect 38334 40402 38386 40414
rect 38334 40338 38386 40350
rect 38670 40402 38722 40414
rect 38670 40338 38722 40350
rect 41582 40402 41634 40414
rect 41582 40338 41634 40350
rect 42702 40402 42754 40414
rect 50766 40402 50818 40414
rect 44034 40350 44046 40402
rect 44098 40350 44110 40402
rect 44258 40350 44270 40402
rect 44322 40350 44334 40402
rect 46610 40350 46622 40402
rect 46674 40350 46686 40402
rect 47394 40350 47406 40402
rect 47458 40350 47470 40402
rect 53230 40402 53282 40414
rect 55022 40402 55074 40414
rect 42702 40338 42754 40350
rect 50766 40338 50818 40350
rect 52446 40346 52498 40358
rect 5406 40290 5458 40302
rect 1922 40238 1934 40290
rect 1986 40238 1998 40290
rect 5406 40226 5458 40238
rect 5854 40290 5906 40302
rect 5854 40226 5906 40238
rect 7870 40290 7922 40302
rect 7870 40226 7922 40238
rect 9102 40290 9154 40302
rect 9102 40226 9154 40238
rect 11118 40290 11170 40302
rect 11118 40226 11170 40238
rect 14142 40290 14194 40302
rect 14142 40226 14194 40238
rect 18286 40290 18338 40302
rect 18286 40226 18338 40238
rect 22206 40290 22258 40302
rect 22206 40226 22258 40238
rect 22654 40290 22706 40302
rect 37326 40290 37378 40302
rect 24658 40238 24670 40290
rect 24722 40238 24734 40290
rect 25666 40238 25678 40290
rect 25730 40238 25742 40290
rect 27682 40238 27694 40290
rect 27746 40238 27758 40290
rect 29138 40238 29150 40290
rect 29202 40238 29214 40290
rect 31154 40238 31166 40290
rect 31218 40238 31230 40290
rect 22654 40226 22706 40238
rect 37326 40226 37378 40238
rect 40014 40290 40066 40302
rect 40014 40226 40066 40238
rect 42926 40290 42978 40302
rect 50430 40290 50482 40302
rect 46834 40238 46846 40290
rect 46898 40238 46910 40290
rect 54114 40350 54126 40402
rect 54178 40350 54190 40402
rect 53230 40338 53282 40350
rect 55022 40338 55074 40350
rect 55806 40402 55858 40414
rect 56130 40350 56142 40402
rect 56194 40350 56206 40402
rect 55806 40338 55858 40350
rect 52446 40282 52498 40294
rect 56702 40290 56754 40302
rect 42926 40226 42978 40238
rect 50430 40226 50482 40238
rect 56702 40226 56754 40238
rect 57374 40290 57426 40302
rect 57374 40226 57426 40238
rect 57934 40290 57986 40302
rect 57934 40226 57986 40238
rect 7310 40178 7362 40190
rect 5506 40126 5518 40178
rect 5570 40175 5582 40178
rect 6178 40175 6190 40178
rect 5570 40129 6190 40175
rect 5570 40126 5582 40129
rect 6178 40126 6190 40129
rect 6242 40126 6254 40178
rect 7310 40114 7362 40126
rect 12350 40178 12402 40190
rect 12350 40114 12402 40126
rect 12574 40178 12626 40190
rect 12574 40114 12626 40126
rect 12798 40178 12850 40190
rect 12798 40114 12850 40126
rect 13806 40178 13858 40190
rect 13806 40114 13858 40126
rect 13918 40178 13970 40190
rect 13918 40114 13970 40126
rect 14366 40178 14418 40190
rect 21646 40178 21698 40190
rect 17602 40126 17614 40178
rect 17666 40175 17678 40178
rect 18274 40175 18286 40178
rect 17666 40129 18286 40175
rect 17666 40126 17678 40129
rect 18274 40126 18286 40129
rect 18338 40126 18350 40178
rect 14366 40114 14418 40126
rect 21646 40114 21698 40126
rect 26014 40178 26066 40190
rect 26014 40114 26066 40126
rect 35086 40178 35138 40190
rect 35086 40114 35138 40126
rect 1344 40010 58576 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 58576 40010
rect 1344 39924 58576 39958
rect 6862 39842 6914 39854
rect 6862 39778 6914 39790
rect 8430 39842 8482 39854
rect 8430 39778 8482 39790
rect 8654 39842 8706 39854
rect 8654 39778 8706 39790
rect 9102 39842 9154 39854
rect 9102 39778 9154 39790
rect 19630 39842 19682 39854
rect 19630 39778 19682 39790
rect 29598 39842 29650 39854
rect 29598 39778 29650 39790
rect 35646 39842 35698 39854
rect 52782 39842 52834 39854
rect 44034 39790 44046 39842
rect 44098 39839 44110 39842
rect 44594 39839 44606 39842
rect 44098 39793 44606 39839
rect 44098 39790 44110 39793
rect 44594 39790 44606 39793
rect 44658 39790 44670 39842
rect 35646 39778 35698 39790
rect 52782 39778 52834 39790
rect 56814 39842 56866 39854
rect 56814 39778 56866 39790
rect 3166 39730 3218 39742
rect 3166 39666 3218 39678
rect 5742 39730 5794 39742
rect 5742 39666 5794 39678
rect 7310 39730 7362 39742
rect 7310 39666 7362 39678
rect 7758 39730 7810 39742
rect 7758 39666 7810 39678
rect 8206 39730 8258 39742
rect 8206 39666 8258 39678
rect 13918 39730 13970 39742
rect 13918 39666 13970 39678
rect 22094 39730 22146 39742
rect 22094 39666 22146 39678
rect 22766 39730 22818 39742
rect 36206 39730 36258 39742
rect 39342 39730 39394 39742
rect 31714 39678 31726 39730
rect 31778 39678 31790 39730
rect 33506 39678 33518 39730
rect 33570 39678 33582 39730
rect 38658 39678 38670 39730
rect 38722 39678 38734 39730
rect 22766 39666 22818 39678
rect 36206 39666 36258 39678
rect 39342 39666 39394 39678
rect 41694 39730 41746 39742
rect 41694 39666 41746 39678
rect 43262 39730 43314 39742
rect 43262 39666 43314 39678
rect 46174 39730 46226 39742
rect 46174 39666 46226 39678
rect 54238 39730 54290 39742
rect 54238 39666 54290 39678
rect 2718 39618 2770 39630
rect 2718 39554 2770 39566
rect 4174 39618 4226 39630
rect 4174 39554 4226 39566
rect 4398 39618 4450 39630
rect 4398 39554 4450 39566
rect 4734 39618 4786 39630
rect 4734 39554 4786 39566
rect 5966 39618 6018 39630
rect 5966 39554 6018 39566
rect 6190 39618 6242 39630
rect 6190 39554 6242 39566
rect 6414 39618 6466 39630
rect 6414 39554 6466 39566
rect 13806 39618 13858 39630
rect 14478 39618 14530 39630
rect 19966 39618 20018 39630
rect 35758 39618 35810 39630
rect 14130 39566 14142 39618
rect 14194 39566 14206 39618
rect 17826 39566 17838 39618
rect 17890 39566 17902 39618
rect 21634 39566 21646 39618
rect 21698 39566 21710 39618
rect 31154 39566 31166 39618
rect 31218 39566 31230 39618
rect 32274 39566 32286 39618
rect 32338 39566 32350 39618
rect 33618 39566 33630 39618
rect 33682 39566 33694 39618
rect 13806 39554 13858 39566
rect 14478 39554 14530 39566
rect 19966 39554 20018 39566
rect 35758 39554 35810 39566
rect 38110 39618 38162 39630
rect 38110 39554 38162 39566
rect 39006 39618 39058 39630
rect 43374 39618 43426 39630
rect 42578 39566 42590 39618
rect 42642 39566 42654 39618
rect 39006 39554 39058 39566
rect 43374 39554 43426 39566
rect 46062 39618 46114 39630
rect 46062 39554 46114 39566
rect 46398 39618 46450 39630
rect 46398 39554 46450 39566
rect 46510 39618 46562 39630
rect 47742 39618 47794 39630
rect 46722 39566 46734 39618
rect 46786 39566 46798 39618
rect 46510 39554 46562 39566
rect 47742 39554 47794 39566
rect 49086 39618 49138 39630
rect 55246 39618 55298 39630
rect 49634 39566 49646 39618
rect 49698 39566 49710 39618
rect 49086 39554 49138 39566
rect 55246 39554 55298 39566
rect 55694 39618 55746 39630
rect 55694 39554 55746 39566
rect 55918 39618 55970 39630
rect 55918 39554 55970 39566
rect 56366 39618 56418 39630
rect 56366 39554 56418 39566
rect 57038 39618 57090 39630
rect 57038 39554 57090 39566
rect 57262 39618 57314 39630
rect 57262 39554 57314 39566
rect 57710 39618 57762 39630
rect 57710 39554 57762 39566
rect 2382 39506 2434 39518
rect 2382 39442 2434 39454
rect 4958 39506 5010 39518
rect 4958 39442 5010 39454
rect 10334 39506 10386 39518
rect 10334 39442 10386 39454
rect 10670 39506 10722 39518
rect 29822 39506 29874 39518
rect 32846 39506 32898 39518
rect 20178 39454 20190 39506
rect 20242 39454 20254 39506
rect 20514 39454 20526 39506
rect 20578 39454 20590 39506
rect 31602 39454 31614 39506
rect 31666 39454 31678 39506
rect 10670 39442 10722 39454
rect 29822 39442 29874 39454
rect 32846 39442 32898 39454
rect 36654 39506 36706 39518
rect 36654 39442 36706 39454
rect 37774 39506 37826 39518
rect 37774 39442 37826 39454
rect 43038 39506 43090 39518
rect 43038 39442 43090 39454
rect 43150 39506 43202 39518
rect 43150 39442 43202 39454
rect 44046 39506 44098 39518
rect 54910 39506 54962 39518
rect 48066 39454 48078 39506
rect 48130 39454 48142 39506
rect 44046 39442 44098 39454
rect 54910 39442 54962 39454
rect 55806 39506 55858 39518
rect 55806 39442 55858 39454
rect 4062 39394 4114 39406
rect 4062 39330 4114 39342
rect 9886 39394 9938 39406
rect 9886 39330 9938 39342
rect 11118 39394 11170 39406
rect 11118 39330 11170 39342
rect 11678 39394 11730 39406
rect 11678 39330 11730 39342
rect 12126 39394 12178 39406
rect 12126 39330 12178 39342
rect 12574 39394 12626 39406
rect 12574 39330 12626 39342
rect 13022 39394 13074 39406
rect 13022 39330 13074 39342
rect 14030 39394 14082 39406
rect 14030 39330 14082 39342
rect 15038 39394 15090 39406
rect 15038 39330 15090 39342
rect 15598 39394 15650 39406
rect 15598 39330 15650 39342
rect 16046 39394 16098 39406
rect 16046 39330 16098 39342
rect 16830 39394 16882 39406
rect 16830 39330 16882 39342
rect 17278 39394 17330 39406
rect 17278 39330 17330 39342
rect 18062 39394 18114 39406
rect 18062 39330 18114 39342
rect 18622 39394 18674 39406
rect 18622 39330 18674 39342
rect 19070 39394 19122 39406
rect 19070 39330 19122 39342
rect 21982 39394 22034 39406
rect 21982 39330 22034 39342
rect 22206 39394 22258 39406
rect 22206 39330 22258 39342
rect 23214 39394 23266 39406
rect 23214 39330 23266 39342
rect 24782 39394 24834 39406
rect 24782 39330 24834 39342
rect 25342 39394 25394 39406
rect 25342 39330 25394 39342
rect 25790 39394 25842 39406
rect 25790 39330 25842 39342
rect 29710 39394 29762 39406
rect 29710 39330 29762 39342
rect 30606 39394 30658 39406
rect 30606 39330 30658 39342
rect 35646 39394 35698 39406
rect 35646 39330 35698 39342
rect 37886 39394 37938 39406
rect 37886 39330 37938 39342
rect 39902 39394 39954 39406
rect 39902 39330 39954 39342
rect 40350 39394 40402 39406
rect 40350 39330 40402 39342
rect 40798 39394 40850 39406
rect 40798 39330 40850 39342
rect 41246 39394 41298 39406
rect 41246 39330 41298 39342
rect 42142 39394 42194 39406
rect 42142 39330 42194 39342
rect 44494 39394 44546 39406
rect 44494 39330 44546 39342
rect 45502 39394 45554 39406
rect 45502 39330 45554 39342
rect 48526 39394 48578 39406
rect 53454 39394 53506 39406
rect 52098 39342 52110 39394
rect 52162 39342 52174 39394
rect 48526 39330 48578 39342
rect 53454 39330 53506 39342
rect 53790 39394 53842 39406
rect 53790 39330 53842 39342
rect 55022 39394 55074 39406
rect 55022 39330 55074 39342
rect 57486 39394 57538 39406
rect 57486 39330 57538 39342
rect 57598 39394 57650 39406
rect 57598 39330 57650 39342
rect 1344 39226 58576 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 58576 39226
rect 1344 39140 58576 39174
rect 3726 39058 3778 39070
rect 3726 38994 3778 39006
rect 5518 39058 5570 39070
rect 5518 38994 5570 39006
rect 6190 39058 6242 39070
rect 6190 38994 6242 39006
rect 7646 39058 7698 39070
rect 7646 38994 7698 39006
rect 8206 39058 8258 39070
rect 8206 38994 8258 39006
rect 11566 39058 11618 39070
rect 11566 38994 11618 39006
rect 14478 39058 14530 39070
rect 14478 38994 14530 39006
rect 21086 39058 21138 39070
rect 21086 38994 21138 39006
rect 22542 39058 22594 39070
rect 37102 39058 37154 39070
rect 40574 39058 40626 39070
rect 33618 39006 33630 39058
rect 33682 39006 33694 39058
rect 39554 39006 39566 39058
rect 39618 39006 39630 39058
rect 22542 38994 22594 39006
rect 37102 38994 37154 39006
rect 40574 38994 40626 39006
rect 41806 39058 41858 39070
rect 47518 39058 47570 39070
rect 46050 39006 46062 39058
rect 46114 39006 46126 39058
rect 41806 38994 41858 39006
rect 47518 38994 47570 39006
rect 48302 39058 48354 39070
rect 48302 38994 48354 39006
rect 48526 39058 48578 39070
rect 48526 38994 48578 39006
rect 50990 39058 51042 39070
rect 50990 38994 51042 39006
rect 51438 39058 51490 39070
rect 51438 38994 51490 39006
rect 52334 39058 52386 39070
rect 57374 39058 57426 39070
rect 54562 39006 54574 39058
rect 54626 39006 54638 39058
rect 56578 39006 56590 39058
rect 56642 39006 56654 39058
rect 52334 38994 52386 39006
rect 8990 38946 9042 38958
rect 8990 38882 9042 38894
rect 12462 38946 12514 38958
rect 12462 38882 12514 38894
rect 15598 38946 15650 38958
rect 15598 38882 15650 38894
rect 16830 38946 16882 38958
rect 16830 38882 16882 38894
rect 16942 38946 16994 38958
rect 16942 38882 16994 38894
rect 18062 38946 18114 38958
rect 18062 38882 18114 38894
rect 20414 38946 20466 38958
rect 20414 38882 20466 38894
rect 20862 38946 20914 38958
rect 20862 38882 20914 38894
rect 21758 38946 21810 38958
rect 21758 38882 21810 38894
rect 22990 38946 23042 38958
rect 22990 38882 23042 38894
rect 24334 38946 24386 38958
rect 28814 38946 28866 38958
rect 25778 38894 25790 38946
rect 25842 38894 25854 38946
rect 24334 38882 24386 38894
rect 28814 38882 28866 38894
rect 30270 38946 30322 38958
rect 30270 38882 30322 38894
rect 34078 38946 34130 38958
rect 34078 38882 34130 38894
rect 34302 38946 34354 38958
rect 34302 38882 34354 38894
rect 38446 38946 38498 38958
rect 38446 38882 38498 38894
rect 42030 38946 42082 38958
rect 42030 38882 42082 38894
rect 43150 38946 43202 38958
rect 43150 38882 43202 38894
rect 44606 38946 44658 38958
rect 44606 38882 44658 38894
rect 46510 38946 46562 38958
rect 46510 38882 46562 38894
rect 47630 38946 47682 38958
rect 47630 38882 47682 38894
rect 51998 38946 52050 38958
rect 51998 38882 52050 38894
rect 54350 38946 54402 38958
rect 54350 38882 54402 38894
rect 4174 38834 4226 38846
rect 4174 38770 4226 38782
rect 4622 38834 4674 38846
rect 4622 38770 4674 38782
rect 4734 38834 4786 38846
rect 4734 38770 4786 38782
rect 5406 38834 5458 38846
rect 5406 38770 5458 38782
rect 7086 38834 7138 38846
rect 8654 38834 8706 38846
rect 7410 38782 7422 38834
rect 7474 38782 7486 38834
rect 7086 38770 7138 38782
rect 8654 38770 8706 38782
rect 10782 38834 10834 38846
rect 10782 38770 10834 38782
rect 10894 38834 10946 38846
rect 10894 38770 10946 38782
rect 11342 38834 11394 38846
rect 11342 38770 11394 38782
rect 13022 38834 13074 38846
rect 13022 38770 13074 38782
rect 14030 38834 14082 38846
rect 14926 38834 14978 38846
rect 14242 38782 14254 38834
rect 14306 38782 14318 38834
rect 14030 38770 14082 38782
rect 14926 38770 14978 38782
rect 15486 38834 15538 38846
rect 15486 38770 15538 38782
rect 15822 38834 15874 38846
rect 15822 38770 15874 38782
rect 16606 38834 16658 38846
rect 16606 38770 16658 38782
rect 17726 38834 17778 38846
rect 17726 38770 17778 38782
rect 17950 38834 18002 38846
rect 17950 38770 18002 38782
rect 19182 38834 19234 38846
rect 24446 38834 24498 38846
rect 30382 38834 30434 38846
rect 21970 38782 21982 38834
rect 22034 38782 22046 38834
rect 22530 38782 22542 38834
rect 22594 38782 22606 38834
rect 25890 38782 25902 38834
rect 25954 38782 25966 38834
rect 26898 38782 26910 38834
rect 26962 38782 26974 38834
rect 29810 38782 29822 38834
rect 29874 38782 29886 38834
rect 19182 38770 19234 38782
rect 24446 38770 24498 38782
rect 30382 38770 30434 38782
rect 34190 38834 34242 38846
rect 34190 38770 34242 38782
rect 35534 38834 35586 38846
rect 35534 38770 35586 38782
rect 36094 38834 36146 38846
rect 36094 38770 36146 38782
rect 36318 38834 36370 38846
rect 36318 38770 36370 38782
rect 36766 38834 36818 38846
rect 36766 38770 36818 38782
rect 37998 38834 38050 38846
rect 37998 38770 38050 38782
rect 38222 38834 38274 38846
rect 38222 38770 38274 38782
rect 39006 38834 39058 38846
rect 42478 38834 42530 38846
rect 48190 38834 48242 38846
rect 50542 38834 50594 38846
rect 54126 38834 54178 38846
rect 41570 38782 41582 38834
rect 41634 38782 41646 38834
rect 44146 38782 44158 38834
rect 44210 38782 44222 38834
rect 44930 38782 44942 38834
rect 44994 38782 45006 38834
rect 49858 38782 49870 38834
rect 49922 38782 49934 38834
rect 53666 38782 53678 38834
rect 53730 38782 53742 38834
rect 39006 38770 39058 38782
rect 42478 38770 42530 38782
rect 48190 38770 48242 38782
rect 50542 38770 50594 38782
rect 54126 38770 54178 38782
rect 6750 38722 6802 38734
rect 6750 38658 6802 38670
rect 9998 38722 10050 38734
rect 9998 38658 10050 38670
rect 10558 38722 10610 38734
rect 10558 38658 10610 38670
rect 12126 38722 12178 38734
rect 12126 38658 12178 38670
rect 13470 38722 13522 38734
rect 16158 38722 16210 38734
rect 13906 38670 13918 38722
rect 13970 38670 13982 38722
rect 13470 38658 13522 38670
rect 16158 38658 16210 38670
rect 19854 38722 19906 38734
rect 19854 38658 19906 38670
rect 22206 38722 22258 38734
rect 22206 38658 22258 38670
rect 23662 38722 23714 38734
rect 23662 38658 23714 38670
rect 25006 38722 25058 38734
rect 27806 38722 27858 38734
rect 26002 38670 26014 38722
rect 26066 38670 26078 38722
rect 27010 38670 27022 38722
rect 27074 38670 27086 38722
rect 25006 38658 25058 38670
rect 27806 38658 27858 38670
rect 28254 38722 28306 38734
rect 28254 38658 28306 38670
rect 36206 38722 36258 38734
rect 36206 38658 36258 38670
rect 38334 38722 38386 38734
rect 38334 38658 38386 38670
rect 39230 38722 39282 38734
rect 39230 38658 39282 38670
rect 40126 38722 40178 38734
rect 45502 38722 45554 38734
rect 41906 38670 41918 38722
rect 41970 38670 41982 38722
rect 40126 38658 40178 38670
rect 45502 38658 45554 38670
rect 47070 38722 47122 38734
rect 50082 38670 50094 38722
rect 50146 38670 50158 38722
rect 47070 38658 47122 38670
rect 5182 38610 5234 38622
rect 7758 38610 7810 38622
rect 14814 38610 14866 38622
rect 6178 38558 6190 38610
rect 6242 38607 6254 38610
rect 6626 38607 6638 38610
rect 6242 38561 6638 38607
rect 6242 38558 6254 38561
rect 6626 38558 6638 38561
rect 6690 38558 6702 38610
rect 12562 38558 12574 38610
rect 12626 38607 12638 38610
rect 12786 38607 12798 38610
rect 12626 38561 12798 38607
rect 12626 38558 12638 38561
rect 12786 38558 12798 38561
rect 12850 38558 12862 38610
rect 5182 38546 5234 38558
rect 7758 38546 7810 38558
rect 14814 38546 14866 38558
rect 18286 38610 18338 38622
rect 18286 38546 18338 38558
rect 18510 38610 18562 38622
rect 18510 38546 18562 38558
rect 21198 38610 21250 38622
rect 21198 38546 21250 38558
rect 24334 38610 24386 38622
rect 45726 38610 45778 38622
rect 29026 38558 29038 38610
rect 29090 38558 29102 38610
rect 43586 38558 43598 38610
rect 43650 38558 43662 38610
rect 54577 38607 54623 39006
rect 57374 38994 57426 39006
rect 57598 39058 57650 39070
rect 57598 38994 57650 39006
rect 55246 38946 55298 38958
rect 55246 38882 55298 38894
rect 57710 38946 57762 38958
rect 57710 38882 57762 38894
rect 56030 38834 56082 38846
rect 56030 38770 56082 38782
rect 54910 38722 54962 38734
rect 54910 38658 54962 38670
rect 56254 38610 56306 38622
rect 55010 38607 55022 38610
rect 54577 38561 55022 38607
rect 55010 38558 55022 38561
rect 55074 38558 55086 38610
rect 24334 38546 24386 38558
rect 45726 38546 45778 38558
rect 56254 38546 56306 38558
rect 1344 38442 58576 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 58576 38442
rect 1344 38356 58576 38390
rect 5070 38274 5122 38286
rect 5070 38210 5122 38222
rect 18510 38274 18562 38286
rect 18510 38210 18562 38222
rect 25230 38274 25282 38286
rect 25230 38210 25282 38222
rect 36766 38274 36818 38286
rect 42030 38274 42082 38286
rect 40786 38222 40798 38274
rect 40850 38222 40862 38274
rect 36766 38210 36818 38222
rect 42030 38210 42082 38222
rect 52782 38274 52834 38286
rect 56130 38222 56142 38274
rect 56194 38222 56206 38274
rect 57250 38222 57262 38274
rect 57314 38222 57326 38274
rect 52782 38210 52834 38222
rect 5630 38162 5682 38174
rect 8206 38162 8258 38174
rect 7410 38110 7422 38162
rect 7474 38110 7486 38162
rect 5630 38098 5682 38110
rect 8206 38098 8258 38110
rect 8766 38162 8818 38174
rect 8766 38098 8818 38110
rect 10222 38162 10274 38174
rect 14478 38162 14530 38174
rect 10994 38110 11006 38162
rect 11058 38110 11070 38162
rect 10222 38098 10274 38110
rect 14478 38098 14530 38110
rect 14590 38162 14642 38174
rect 14590 38098 14642 38110
rect 17390 38162 17442 38174
rect 17390 38098 17442 38110
rect 20862 38162 20914 38174
rect 20862 38098 20914 38110
rect 23214 38162 23266 38174
rect 23214 38098 23266 38110
rect 30046 38162 30098 38174
rect 33966 38162 34018 38174
rect 50206 38162 50258 38174
rect 30706 38110 30718 38162
rect 30770 38110 30782 38162
rect 34850 38110 34862 38162
rect 34914 38110 34926 38162
rect 36530 38110 36542 38162
rect 36594 38110 36606 38162
rect 40562 38110 40574 38162
rect 40626 38110 40638 38162
rect 43362 38110 43374 38162
rect 43426 38110 43438 38162
rect 30046 38098 30098 38110
rect 33966 38098 34018 38110
rect 50206 38098 50258 38110
rect 53342 38162 53394 38174
rect 57822 38162 57874 38174
rect 55794 38110 55806 38162
rect 55858 38110 55870 38162
rect 53342 38098 53394 38110
rect 57822 38098 57874 38110
rect 3614 38050 3666 38062
rect 3614 37986 3666 37998
rect 4174 38050 4226 38062
rect 5742 38050 5794 38062
rect 4610 37998 4622 38050
rect 4674 37998 4686 38050
rect 4174 37986 4226 37998
rect 5742 37986 5794 37998
rect 6302 38050 6354 38062
rect 9662 38050 9714 38062
rect 12238 38050 12290 38062
rect 7746 37998 7758 38050
rect 7810 37998 7822 38050
rect 11442 37998 11454 38050
rect 11506 37998 11518 38050
rect 6302 37986 6354 37998
rect 9662 37986 9714 37998
rect 12238 37986 12290 37998
rect 12686 38050 12738 38062
rect 12686 37986 12738 37998
rect 12910 38050 12962 38062
rect 17614 38050 17666 38062
rect 14018 37998 14030 38050
rect 14082 37998 14094 38050
rect 14802 37998 14814 38050
rect 14866 37998 14878 38050
rect 12910 37986 12962 37998
rect 17614 37986 17666 37998
rect 19518 38050 19570 38062
rect 19518 37986 19570 37998
rect 19742 38050 19794 38062
rect 25454 38050 25506 38062
rect 27806 38050 27858 38062
rect 30158 38050 30210 38062
rect 34078 38050 34130 38062
rect 22194 37998 22206 38050
rect 22258 37998 22270 38050
rect 23986 37998 23998 38050
rect 24050 37998 24062 38050
rect 25890 37998 25902 38050
rect 25954 37998 25966 38050
rect 28354 37998 28366 38050
rect 28418 37998 28430 38050
rect 33506 37998 33518 38050
rect 33570 37998 33582 38050
rect 19742 37986 19794 37998
rect 25454 37986 25506 37998
rect 27806 37986 27858 37998
rect 30158 37986 30210 37998
rect 34078 37986 34130 37998
rect 35982 38050 36034 38062
rect 35982 37986 36034 37998
rect 36206 38050 36258 38062
rect 36206 37986 36258 37998
rect 37438 38050 37490 38062
rect 37438 37986 37490 37998
rect 37774 38050 37826 38062
rect 37774 37986 37826 37998
rect 39342 38050 39394 38062
rect 41694 38050 41746 38062
rect 40450 37998 40462 38050
rect 40514 37998 40526 38050
rect 39342 37986 39394 37998
rect 41694 37986 41746 37998
rect 45838 38050 45890 38062
rect 45838 37986 45890 37998
rect 51886 38050 51938 38062
rect 51886 37986 51938 37998
rect 52110 38050 52162 38062
rect 52110 37986 52162 37998
rect 52334 38050 52386 38062
rect 52334 37986 52386 37998
rect 54910 38050 54962 38062
rect 57598 38050 57650 38062
rect 56018 37998 56030 38050
rect 56082 37998 56094 38050
rect 54910 37986 54962 37998
rect 57598 37986 57650 37998
rect 4286 37938 4338 37950
rect 4286 37874 4338 37886
rect 4398 37938 4450 37950
rect 4398 37874 4450 37886
rect 5966 37938 6018 37950
rect 5966 37874 6018 37886
rect 11006 37938 11058 37950
rect 11006 37874 11058 37886
rect 11230 37938 11282 37950
rect 16046 37938 16098 37950
rect 15026 37886 15038 37938
rect 15090 37886 15102 37938
rect 11230 37874 11282 37886
rect 16046 37874 16098 37886
rect 16158 37938 16210 37950
rect 18846 37938 18898 37950
rect 16258 37886 16270 37938
rect 16322 37886 16334 37938
rect 16158 37874 16210 37886
rect 18846 37874 18898 37886
rect 20078 37938 20130 37950
rect 20078 37874 20130 37886
rect 22430 37938 22482 37950
rect 27694 37938 27746 37950
rect 24322 37886 24334 37938
rect 24386 37886 24398 37938
rect 22430 37874 22482 37886
rect 27694 37874 27746 37886
rect 31054 37938 31106 37950
rect 31054 37874 31106 37886
rect 31838 37938 31890 37950
rect 31838 37874 31890 37886
rect 34862 37938 34914 37950
rect 34862 37874 34914 37886
rect 35310 37938 35362 37950
rect 35310 37874 35362 37886
rect 36542 37938 36594 37950
rect 36542 37874 36594 37886
rect 37662 37938 37714 37950
rect 37662 37874 37714 37886
rect 39006 37938 39058 37950
rect 39006 37874 39058 37886
rect 41470 37938 41522 37950
rect 43262 37938 43314 37950
rect 43138 37886 43150 37938
rect 43202 37886 43214 37938
rect 41470 37874 41522 37886
rect 43262 37874 43314 37886
rect 44046 37938 44098 37950
rect 44046 37874 44098 37886
rect 45502 37938 45554 37950
rect 45502 37874 45554 37886
rect 48750 37938 48802 37950
rect 48750 37874 48802 37886
rect 55022 37938 55074 37950
rect 55022 37874 55074 37886
rect 6190 37826 6242 37838
rect 6190 37762 6242 37774
rect 9102 37826 9154 37838
rect 9102 37762 9154 37774
rect 10894 37826 10946 37838
rect 10894 37762 10946 37774
rect 12350 37826 12402 37838
rect 12350 37762 12402 37774
rect 12462 37826 12514 37838
rect 12462 37762 12514 37774
rect 15822 37826 15874 37838
rect 15822 37762 15874 37774
rect 15934 37826 15986 37838
rect 18622 37826 18674 37838
rect 17938 37774 17950 37826
rect 18002 37774 18014 37826
rect 15934 37762 15986 37774
rect 18622 37762 18674 37774
rect 19630 37826 19682 37838
rect 19630 37762 19682 37774
rect 21534 37826 21586 37838
rect 21534 37762 21586 37774
rect 29710 37826 29762 37838
rect 29710 37762 29762 37774
rect 29934 37826 29986 37838
rect 29934 37762 29986 37774
rect 30830 37826 30882 37838
rect 30830 37762 30882 37774
rect 31502 37826 31554 37838
rect 31502 37762 31554 37774
rect 31726 37826 31778 37838
rect 31726 37762 31778 37774
rect 32398 37826 32450 37838
rect 32398 37762 32450 37774
rect 32734 37826 32786 37838
rect 32734 37762 32786 37774
rect 33854 37826 33906 37838
rect 33854 37762 33906 37774
rect 35086 37826 35138 37838
rect 35086 37762 35138 37774
rect 38446 37826 38498 37838
rect 38446 37762 38498 37774
rect 43374 37826 43426 37838
rect 43374 37762 43426 37774
rect 43598 37826 43650 37838
rect 43598 37762 43650 37774
rect 44494 37826 44546 37838
rect 44494 37762 44546 37774
rect 45614 37826 45666 37838
rect 45614 37762 45666 37774
rect 46174 37826 46226 37838
rect 46174 37762 46226 37774
rect 46622 37826 46674 37838
rect 46622 37762 46674 37774
rect 47182 37826 47234 37838
rect 47182 37762 47234 37774
rect 47966 37826 48018 37838
rect 47966 37762 48018 37774
rect 48302 37826 48354 37838
rect 48302 37762 48354 37774
rect 49422 37826 49474 37838
rect 49422 37762 49474 37774
rect 49758 37826 49810 37838
rect 49758 37762 49810 37774
rect 50654 37826 50706 37838
rect 50654 37762 50706 37774
rect 51214 37826 51266 37838
rect 51214 37762 51266 37774
rect 53790 37826 53842 37838
rect 53790 37762 53842 37774
rect 54798 37826 54850 37838
rect 54798 37762 54850 37774
rect 1344 37658 58576 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 58576 37658
rect 1344 37572 58576 37606
rect 4062 37490 4114 37502
rect 4062 37426 4114 37438
rect 4734 37490 4786 37502
rect 4734 37426 4786 37438
rect 4846 37490 4898 37502
rect 4846 37426 4898 37438
rect 4958 37490 5010 37502
rect 7086 37490 7138 37502
rect 6850 37438 6862 37490
rect 6914 37438 6926 37490
rect 4958 37426 5010 37438
rect 7086 37426 7138 37438
rect 8094 37490 8146 37502
rect 8094 37426 8146 37438
rect 10558 37490 10610 37502
rect 10558 37426 10610 37438
rect 12238 37490 12290 37502
rect 12238 37426 12290 37438
rect 13918 37490 13970 37502
rect 25566 37490 25618 37502
rect 20626 37438 20638 37490
rect 20690 37438 20702 37490
rect 13918 37426 13970 37438
rect 25566 37426 25618 37438
rect 26350 37490 26402 37502
rect 26350 37426 26402 37438
rect 27358 37490 27410 37502
rect 27358 37426 27410 37438
rect 27470 37490 27522 37502
rect 27470 37426 27522 37438
rect 32958 37490 33010 37502
rect 32958 37426 33010 37438
rect 35310 37490 35362 37502
rect 35310 37426 35362 37438
rect 36878 37490 36930 37502
rect 36878 37426 36930 37438
rect 36990 37490 37042 37502
rect 36990 37426 37042 37438
rect 38334 37490 38386 37502
rect 38334 37426 38386 37438
rect 39566 37490 39618 37502
rect 39566 37426 39618 37438
rect 44158 37490 44210 37502
rect 44158 37426 44210 37438
rect 47406 37490 47458 37502
rect 52658 37438 52670 37490
rect 52722 37438 52734 37490
rect 47406 37426 47458 37438
rect 11454 37378 11506 37390
rect 11454 37314 11506 37326
rect 13806 37378 13858 37390
rect 16718 37378 16770 37390
rect 22654 37378 22706 37390
rect 25790 37378 25842 37390
rect 14578 37326 14590 37378
rect 14642 37326 14654 37378
rect 19842 37326 19854 37378
rect 19906 37326 19918 37378
rect 20850 37326 20862 37378
rect 20914 37326 20926 37378
rect 24098 37326 24110 37378
rect 24162 37326 24174 37378
rect 13806 37314 13858 37326
rect 16718 37314 16770 37326
rect 22654 37314 22706 37326
rect 25790 37314 25842 37326
rect 25902 37378 25954 37390
rect 25902 37314 25954 37326
rect 27582 37378 27634 37390
rect 27582 37314 27634 37326
rect 28030 37378 28082 37390
rect 28030 37314 28082 37326
rect 28814 37378 28866 37390
rect 28814 37314 28866 37326
rect 32622 37378 32674 37390
rect 32622 37314 32674 37326
rect 32734 37378 32786 37390
rect 41694 37378 41746 37390
rect 39890 37326 39902 37378
rect 39954 37326 39966 37378
rect 32734 37314 32786 37326
rect 41694 37314 41746 37326
rect 46398 37378 46450 37390
rect 50206 37378 50258 37390
rect 48290 37326 48302 37378
rect 48354 37326 48366 37378
rect 46398 37314 46450 37326
rect 50206 37314 50258 37326
rect 53566 37378 53618 37390
rect 53566 37314 53618 37326
rect 57374 37378 57426 37390
rect 57374 37314 57426 37326
rect 6862 37266 6914 37278
rect 4498 37214 4510 37266
rect 4562 37214 4574 37266
rect 5170 37214 5182 37266
rect 5234 37214 5246 37266
rect 6862 37202 6914 37214
rect 7310 37266 7362 37278
rect 7310 37202 7362 37214
rect 7422 37266 7474 37278
rect 7422 37202 7474 37214
rect 11902 37266 11954 37278
rect 14366 37266 14418 37278
rect 18398 37266 18450 37278
rect 13346 37214 13358 37266
rect 13410 37214 13422 37266
rect 13570 37214 13582 37266
rect 13634 37214 13646 37266
rect 14914 37214 14926 37266
rect 14978 37214 14990 37266
rect 15586 37214 15598 37266
rect 15650 37214 15662 37266
rect 11902 37202 11954 37214
rect 14366 37202 14418 37214
rect 18398 37202 18450 37214
rect 19070 37266 19122 37278
rect 23886 37266 23938 37278
rect 33630 37266 33682 37278
rect 19954 37214 19966 37266
rect 20018 37214 20030 37266
rect 20626 37214 20638 37266
rect 20690 37214 20702 37266
rect 21522 37214 21534 37266
rect 21586 37214 21598 37266
rect 23426 37214 23438 37266
rect 23490 37214 23502 37266
rect 24658 37214 24670 37266
rect 24722 37214 24734 37266
rect 29698 37214 29710 37266
rect 29762 37214 29774 37266
rect 31826 37214 31838 37266
rect 31890 37214 31902 37266
rect 19070 37202 19122 37214
rect 23886 37202 23938 37214
rect 33630 37202 33682 37214
rect 33742 37266 33794 37278
rect 36206 37266 36258 37278
rect 34066 37214 34078 37266
rect 34130 37214 34142 37266
rect 33742 37202 33794 37214
rect 36206 37202 36258 37214
rect 36766 37266 36818 37278
rect 36766 37202 36818 37214
rect 37438 37266 37490 37278
rect 37438 37202 37490 37214
rect 41806 37266 41858 37278
rect 41806 37202 41858 37214
rect 41918 37266 41970 37278
rect 41918 37202 41970 37214
rect 42814 37266 42866 37278
rect 42814 37202 42866 37214
rect 43934 37266 43986 37278
rect 43934 37202 43986 37214
rect 44158 37266 44210 37278
rect 44158 37202 44210 37214
rect 44494 37266 44546 37278
rect 44494 37202 44546 37214
rect 46734 37266 46786 37278
rect 50766 37266 50818 37278
rect 48402 37214 48414 37266
rect 48466 37214 48478 37266
rect 50418 37214 50430 37266
rect 50482 37214 50494 37266
rect 46734 37202 46786 37214
rect 50766 37202 50818 37214
rect 52782 37266 52834 37278
rect 52994 37214 53006 37266
rect 53058 37214 53070 37266
rect 56354 37214 56366 37266
rect 56418 37214 56430 37266
rect 52782 37202 52834 37214
rect 5630 37154 5682 37166
rect 5630 37090 5682 37102
rect 6302 37154 6354 37166
rect 6302 37090 6354 37102
rect 11006 37154 11058 37166
rect 11006 37090 11058 37102
rect 12910 37154 12962 37166
rect 12910 37090 12962 37102
rect 14254 37154 14306 37166
rect 17726 37154 17778 37166
rect 16594 37102 16606 37154
rect 16658 37102 16670 37154
rect 14254 37090 14306 37102
rect 17726 37090 17778 37102
rect 18174 37154 18226 37166
rect 31054 37154 31106 37166
rect 37998 37154 38050 37166
rect 24546 37102 24558 37154
rect 24610 37102 24622 37154
rect 29474 37102 29486 37154
rect 29538 37102 29550 37154
rect 31154 37102 31166 37154
rect 31218 37102 31230 37154
rect 18174 37090 18226 37102
rect 31054 37090 31106 37102
rect 37998 37090 38050 37102
rect 38782 37154 38834 37166
rect 38782 37090 38834 37102
rect 40350 37154 40402 37166
rect 40350 37090 40402 37102
rect 40798 37154 40850 37166
rect 40798 37090 40850 37102
rect 43262 37154 43314 37166
rect 43262 37090 43314 37102
rect 44942 37154 44994 37166
rect 44942 37090 44994 37102
rect 45502 37154 45554 37166
rect 45502 37090 45554 37102
rect 45950 37154 46002 37166
rect 45950 37090 46002 37102
rect 49534 37154 49586 37166
rect 51214 37154 51266 37166
rect 57822 37154 57874 37166
rect 50306 37102 50318 37154
rect 50370 37102 50382 37154
rect 55682 37102 55694 37154
rect 55746 37102 55758 37154
rect 49534 37090 49586 37102
rect 51214 37090 51266 37102
rect 57822 37090 57874 37102
rect 16942 37042 16994 37054
rect 16942 36978 16994 36990
rect 18622 37042 18674 37054
rect 18622 36978 18674 36990
rect 35758 37042 35810 37054
rect 35758 36978 35810 36990
rect 35982 37042 36034 37054
rect 47742 37042 47794 37054
rect 37650 36990 37662 37042
rect 37714 37039 37726 37042
rect 38434 37039 38446 37042
rect 37714 36993 38446 37039
rect 37714 36990 37726 36993
rect 38434 36990 38446 36993
rect 38498 36990 38510 37042
rect 42354 36990 42366 37042
rect 42418 36990 42430 37042
rect 42578 36990 42590 37042
rect 42642 37039 42654 37042
rect 43586 37039 43598 37042
rect 42642 36993 43598 37039
rect 42642 36990 42654 36993
rect 43586 36990 43598 36993
rect 43650 36990 43662 37042
rect 35982 36978 36034 36990
rect 47742 36978 47794 36990
rect 1344 36874 58576 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 58576 36874
rect 1344 36788 58576 36822
rect 38670 36706 38722 36718
rect 7410 36654 7422 36706
rect 7474 36703 7486 36706
rect 7634 36703 7646 36706
rect 7474 36657 7646 36703
rect 7474 36654 7486 36657
rect 7634 36654 7646 36657
rect 7698 36654 7710 36706
rect 38670 36642 38722 36654
rect 45502 36706 45554 36718
rect 54338 36654 54350 36706
rect 54402 36703 54414 36706
rect 55234 36703 55246 36706
rect 54402 36657 55246 36703
rect 54402 36654 54414 36657
rect 55234 36654 55246 36657
rect 55298 36654 55310 36706
rect 45502 36642 45554 36654
rect 7870 36594 7922 36606
rect 9550 36594 9602 36606
rect 8754 36542 8766 36594
rect 8818 36542 8830 36594
rect 7870 36530 7922 36542
rect 9550 36530 9602 36542
rect 13918 36594 13970 36606
rect 13918 36530 13970 36542
rect 15598 36594 15650 36606
rect 15598 36530 15650 36542
rect 16270 36594 16322 36606
rect 16270 36530 16322 36542
rect 18734 36594 18786 36606
rect 33182 36594 33234 36606
rect 24322 36542 24334 36594
rect 24386 36542 24398 36594
rect 18734 36530 18786 36542
rect 33182 36530 33234 36542
rect 37438 36594 37490 36606
rect 52222 36594 52274 36606
rect 47954 36542 47966 36594
rect 48018 36542 48030 36594
rect 37438 36530 37490 36542
rect 52222 36530 52274 36542
rect 56142 36594 56194 36606
rect 56142 36530 56194 36542
rect 14814 36482 14866 36494
rect 16718 36482 16770 36494
rect 8306 36430 8318 36482
rect 8370 36430 8382 36482
rect 9762 36430 9774 36482
rect 9826 36430 9838 36482
rect 15138 36430 15150 36482
rect 15202 36430 15214 36482
rect 14814 36418 14866 36430
rect 16718 36418 16770 36430
rect 19854 36482 19906 36494
rect 19854 36418 19906 36430
rect 20190 36482 20242 36494
rect 20190 36418 20242 36430
rect 27134 36482 27186 36494
rect 27134 36418 27186 36430
rect 32286 36482 32338 36494
rect 33630 36482 33682 36494
rect 32722 36430 32734 36482
rect 32786 36430 32798 36482
rect 32286 36418 32338 36430
rect 33630 36418 33682 36430
rect 39678 36482 39730 36494
rect 39678 36418 39730 36430
rect 45838 36482 45890 36494
rect 52110 36482 52162 36494
rect 48066 36430 48078 36482
rect 48130 36430 48142 36482
rect 49634 36430 49646 36482
rect 49698 36430 49710 36482
rect 51202 36430 51214 36482
rect 51266 36430 51278 36482
rect 45838 36418 45890 36430
rect 52110 36418 52162 36430
rect 52670 36482 52722 36494
rect 52670 36418 52722 36430
rect 53902 36482 53954 36494
rect 57710 36482 57762 36494
rect 54226 36430 54238 36482
rect 54290 36430 54302 36482
rect 57250 36430 57262 36482
rect 57314 36430 57326 36482
rect 53902 36418 53954 36430
rect 57710 36418 57762 36430
rect 9438 36370 9490 36382
rect 9438 36306 9490 36318
rect 14366 36370 14418 36382
rect 17278 36370 17330 36382
rect 14578 36318 14590 36370
rect 14642 36318 14654 36370
rect 14366 36306 14418 36318
rect 17278 36306 17330 36318
rect 20414 36370 20466 36382
rect 20414 36306 20466 36318
rect 21646 36370 21698 36382
rect 21646 36306 21698 36318
rect 21982 36370 22034 36382
rect 24782 36370 24834 36382
rect 24546 36318 24558 36370
rect 24610 36318 24622 36370
rect 21982 36306 22034 36318
rect 24782 36306 24834 36318
rect 24894 36370 24946 36382
rect 24894 36306 24946 36318
rect 37998 36370 38050 36382
rect 37998 36306 38050 36318
rect 38782 36370 38834 36382
rect 38782 36306 38834 36318
rect 40574 36370 40626 36382
rect 40574 36306 40626 36318
rect 43038 36370 43090 36382
rect 43038 36306 43090 36318
rect 43262 36370 43314 36382
rect 43262 36306 43314 36318
rect 43822 36370 43874 36382
rect 43822 36306 43874 36318
rect 44158 36370 44210 36382
rect 44158 36306 44210 36318
rect 46062 36370 46114 36382
rect 46062 36306 46114 36318
rect 47294 36370 47346 36382
rect 52446 36370 52498 36382
rect 48178 36318 48190 36370
rect 48242 36318 48254 36370
rect 47294 36306 47346 36318
rect 52446 36306 52498 36318
rect 53454 36370 53506 36382
rect 56814 36370 56866 36382
rect 53666 36318 53678 36370
rect 53730 36318 53742 36370
rect 53454 36306 53506 36318
rect 56814 36306 56866 36318
rect 5070 36258 5122 36270
rect 5070 36194 5122 36206
rect 6078 36258 6130 36270
rect 6078 36194 6130 36206
rect 6526 36258 6578 36270
rect 6526 36194 6578 36206
rect 6974 36258 7026 36270
rect 6974 36194 7026 36206
rect 7310 36258 7362 36270
rect 7310 36194 7362 36206
rect 10222 36258 10274 36270
rect 10222 36194 10274 36206
rect 11006 36258 11058 36270
rect 11006 36194 11058 36206
rect 12014 36258 12066 36270
rect 12014 36194 12066 36206
rect 12462 36258 12514 36270
rect 12462 36194 12514 36206
rect 12910 36258 12962 36270
rect 17166 36258 17218 36270
rect 14690 36206 14702 36258
rect 14754 36206 14766 36258
rect 12910 36194 12962 36206
rect 17166 36194 17218 36206
rect 17726 36258 17778 36270
rect 17726 36194 17778 36206
rect 18174 36258 18226 36270
rect 18174 36194 18226 36206
rect 19182 36258 19234 36270
rect 19182 36194 19234 36206
rect 20078 36258 20130 36270
rect 20078 36194 20130 36206
rect 23774 36258 23826 36270
rect 23774 36194 23826 36206
rect 25118 36258 25170 36270
rect 25118 36194 25170 36206
rect 25678 36258 25730 36270
rect 25678 36194 25730 36206
rect 26014 36258 26066 36270
rect 26014 36194 26066 36206
rect 26798 36258 26850 36270
rect 26798 36194 26850 36206
rect 31278 36258 31330 36270
rect 31278 36194 31330 36206
rect 36430 36258 36482 36270
rect 36430 36194 36482 36206
rect 38670 36258 38722 36270
rect 38670 36194 38722 36206
rect 39342 36258 39394 36270
rect 39342 36194 39394 36206
rect 40238 36258 40290 36270
rect 40238 36194 40290 36206
rect 41022 36258 41074 36270
rect 41022 36194 41074 36206
rect 41582 36258 41634 36270
rect 41582 36194 41634 36206
rect 41918 36258 41970 36270
rect 41918 36194 41970 36206
rect 42478 36258 42530 36270
rect 42478 36194 42530 36206
rect 43150 36258 43202 36270
rect 43150 36194 43202 36206
rect 44606 36258 44658 36270
rect 44606 36194 44658 36206
rect 46734 36258 46786 36270
rect 54798 36258 54850 36270
rect 53778 36206 53790 36258
rect 53842 36206 53854 36258
rect 46734 36194 46786 36206
rect 54798 36194 54850 36206
rect 55134 36258 55186 36270
rect 55134 36194 55186 36206
rect 55582 36258 55634 36270
rect 55582 36194 55634 36206
rect 56254 36258 56306 36270
rect 56254 36194 56306 36206
rect 1344 36090 58576 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 58576 36090
rect 1344 36004 58576 36038
rect 7086 35922 7138 35934
rect 7086 35858 7138 35870
rect 7198 35922 7250 35934
rect 7198 35858 7250 35870
rect 8318 35922 8370 35934
rect 8318 35858 8370 35870
rect 8654 35922 8706 35934
rect 8654 35858 8706 35870
rect 9998 35922 10050 35934
rect 9998 35858 10050 35870
rect 13134 35922 13186 35934
rect 16942 35922 16994 35934
rect 14130 35870 14142 35922
rect 14194 35870 14206 35922
rect 16594 35870 16606 35922
rect 16658 35870 16670 35922
rect 13134 35858 13186 35870
rect 16942 35858 16994 35870
rect 17726 35922 17778 35934
rect 17726 35858 17778 35870
rect 30494 35922 30546 35934
rect 32398 35922 32450 35934
rect 31826 35870 31838 35922
rect 31890 35870 31902 35922
rect 30494 35858 30546 35870
rect 32398 35858 32450 35870
rect 35646 35922 35698 35934
rect 35646 35858 35698 35870
rect 36990 35922 37042 35934
rect 36990 35858 37042 35870
rect 38558 35922 38610 35934
rect 48302 35922 48354 35934
rect 51662 35922 51714 35934
rect 57822 35922 57874 35934
rect 45714 35870 45726 35922
rect 45778 35870 45790 35922
rect 46274 35870 46286 35922
rect 46338 35870 46350 35922
rect 51090 35870 51102 35922
rect 51154 35870 51166 35922
rect 52658 35870 52670 35922
rect 52722 35870 52734 35922
rect 38558 35858 38610 35870
rect 48302 35858 48354 35870
rect 51662 35858 51714 35870
rect 57822 35858 57874 35870
rect 4398 35810 4450 35822
rect 4398 35746 4450 35758
rect 8878 35810 8930 35822
rect 8878 35746 8930 35758
rect 11230 35810 11282 35822
rect 11230 35746 11282 35758
rect 11790 35810 11842 35822
rect 11790 35746 11842 35758
rect 12462 35810 12514 35822
rect 12462 35746 12514 35758
rect 12910 35810 12962 35822
rect 20414 35810 20466 35822
rect 14018 35758 14030 35810
rect 14082 35758 14094 35810
rect 18050 35758 18062 35810
rect 18114 35758 18126 35810
rect 12910 35746 12962 35758
rect 20414 35746 20466 35758
rect 36318 35810 36370 35822
rect 36318 35746 36370 35758
rect 36430 35810 36482 35822
rect 36430 35746 36482 35758
rect 37438 35810 37490 35822
rect 37438 35746 37490 35758
rect 38222 35810 38274 35822
rect 38222 35746 38274 35758
rect 42926 35810 42978 35822
rect 44606 35810 44658 35822
rect 43698 35758 43710 35810
rect 43762 35758 43774 35810
rect 42926 35746 42978 35758
rect 44606 35746 44658 35758
rect 50542 35810 50594 35822
rect 50542 35746 50594 35758
rect 51550 35810 51602 35822
rect 51550 35746 51602 35758
rect 51886 35810 51938 35822
rect 56590 35810 56642 35822
rect 54002 35758 54014 35810
rect 54066 35758 54078 35810
rect 51886 35746 51938 35758
rect 56590 35746 56642 35758
rect 57486 35810 57538 35822
rect 57486 35746 57538 35758
rect 58046 35810 58098 35822
rect 58046 35746 58098 35758
rect 6526 35698 6578 35710
rect 4946 35646 4958 35698
rect 5010 35646 5022 35698
rect 6526 35634 6578 35646
rect 6974 35698 7026 35710
rect 6974 35634 7026 35646
rect 8990 35698 9042 35710
rect 8990 35634 9042 35646
rect 10222 35698 10274 35710
rect 10670 35698 10722 35710
rect 20078 35698 20130 35710
rect 10322 35646 10334 35698
rect 10386 35646 10398 35698
rect 14242 35646 14254 35698
rect 14306 35646 14318 35698
rect 14802 35646 14814 35698
rect 14866 35646 14878 35698
rect 15362 35646 15374 35698
rect 15426 35646 15438 35698
rect 19842 35646 19854 35698
rect 19906 35646 19918 35698
rect 10222 35634 10274 35646
rect 10670 35634 10722 35646
rect 20078 35634 20130 35646
rect 24110 35698 24162 35710
rect 24110 35634 24162 35646
rect 24670 35698 24722 35710
rect 24670 35634 24722 35646
rect 30046 35698 30098 35710
rect 30046 35634 30098 35646
rect 30718 35698 30770 35710
rect 30718 35634 30770 35646
rect 31502 35698 31554 35710
rect 31502 35634 31554 35646
rect 35310 35698 35362 35710
rect 35310 35634 35362 35646
rect 38446 35698 38498 35710
rect 38446 35634 38498 35646
rect 38670 35698 38722 35710
rect 45166 35698 45218 35710
rect 38882 35646 38894 35698
rect 38946 35646 38958 35698
rect 39554 35646 39566 35698
rect 39618 35646 39630 35698
rect 39890 35646 39902 35698
rect 39954 35646 39966 35698
rect 40898 35646 40910 35698
rect 40962 35646 40974 35698
rect 43138 35646 43150 35698
rect 43202 35646 43214 35698
rect 43586 35646 43598 35698
rect 43650 35646 43662 35698
rect 38670 35634 38722 35646
rect 45166 35634 45218 35646
rect 46846 35698 46898 35710
rect 46846 35634 46898 35646
rect 48190 35698 48242 35710
rect 48190 35634 48242 35646
rect 48526 35698 48578 35710
rect 48526 35634 48578 35646
rect 48750 35698 48802 35710
rect 48750 35634 48802 35646
rect 50430 35698 50482 35710
rect 50430 35634 50482 35646
rect 50654 35698 50706 35710
rect 50654 35634 50706 35646
rect 52222 35698 52274 35710
rect 57710 35698 57762 35710
rect 52882 35646 52894 35698
rect 52946 35646 52958 35698
rect 52222 35634 52274 35646
rect 57710 35634 57762 35646
rect 6078 35586 6130 35598
rect 7758 35586 7810 35598
rect 5282 35534 5294 35586
rect 5346 35534 5358 35586
rect 6402 35534 6414 35586
rect 6466 35534 6478 35586
rect 6078 35522 6130 35534
rect 6066 35422 6078 35474
rect 6130 35471 6142 35474
rect 6417 35471 6463 35534
rect 7758 35522 7810 35534
rect 10110 35586 10162 35598
rect 16046 35586 16098 35598
rect 13234 35534 13246 35586
rect 13298 35534 13310 35586
rect 10110 35522 10162 35534
rect 16046 35522 16098 35534
rect 18846 35586 18898 35598
rect 18846 35522 18898 35534
rect 19294 35586 19346 35598
rect 19294 35522 19346 35534
rect 20862 35586 20914 35598
rect 20862 35522 20914 35534
rect 21422 35586 21474 35598
rect 21422 35522 21474 35534
rect 21870 35586 21922 35598
rect 21870 35522 21922 35534
rect 25566 35586 25618 35598
rect 25566 35522 25618 35534
rect 26126 35586 26178 35598
rect 26126 35522 26178 35534
rect 30606 35586 30658 35598
rect 30606 35522 30658 35534
rect 32734 35586 32786 35598
rect 32734 35522 32786 35534
rect 34750 35586 34802 35598
rect 34750 35522 34802 35534
rect 41470 35586 41522 35598
rect 41470 35522 41522 35534
rect 41918 35586 41970 35598
rect 47742 35586 47794 35598
rect 43474 35534 43486 35586
rect 43538 35534 43550 35586
rect 41918 35522 41970 35534
rect 47742 35522 47794 35534
rect 49534 35586 49586 35598
rect 49534 35522 49586 35534
rect 6130 35425 6463 35471
rect 11342 35474 11394 35486
rect 6130 35422 6142 35425
rect 11342 35410 11394 35422
rect 20302 35474 20354 35486
rect 20302 35410 20354 35422
rect 36430 35474 36482 35486
rect 36430 35410 36482 35422
rect 40686 35474 40738 35486
rect 40686 35410 40738 35422
rect 45390 35474 45442 35486
rect 45390 35410 45442 35422
rect 46622 35474 46674 35486
rect 46622 35410 46674 35422
rect 56254 35474 56306 35486
rect 56254 35410 56306 35422
rect 1344 35306 58576 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 58576 35306
rect 1344 35220 58576 35254
rect 4846 35138 4898 35150
rect 4050 35086 4062 35138
rect 4114 35135 4126 35138
rect 4274 35135 4286 35138
rect 4114 35089 4286 35135
rect 4114 35086 4126 35089
rect 4274 35086 4286 35089
rect 4338 35086 4350 35138
rect 4846 35074 4898 35086
rect 8654 35138 8706 35150
rect 8654 35074 8706 35086
rect 10334 35138 10386 35150
rect 32398 35138 32450 35150
rect 15362 35086 15374 35138
rect 15426 35086 15438 35138
rect 18274 35086 18286 35138
rect 18338 35086 18350 35138
rect 10334 35074 10386 35086
rect 32398 35074 32450 35086
rect 36094 35138 36146 35150
rect 36094 35074 36146 35086
rect 36430 35138 36482 35150
rect 41010 35086 41022 35138
rect 41074 35086 41086 35138
rect 36430 35074 36482 35086
rect 6190 35026 6242 35038
rect 6190 34962 6242 34974
rect 7198 35026 7250 35038
rect 7198 34962 7250 34974
rect 9102 35026 9154 35038
rect 9102 34962 9154 34974
rect 9550 35026 9602 35038
rect 9550 34962 9602 34974
rect 12238 35026 12290 35038
rect 17390 35026 17442 35038
rect 19854 35026 19906 35038
rect 24334 35026 24386 35038
rect 14354 34974 14366 35026
rect 14418 34974 14430 35026
rect 18386 34974 18398 35026
rect 18450 34974 18462 35026
rect 20290 34974 20302 35026
rect 20354 34974 20366 35026
rect 12238 34962 12290 34974
rect 17390 34962 17442 34974
rect 19854 34962 19906 34974
rect 24334 34962 24386 34974
rect 28366 35026 28418 35038
rect 28366 34962 28418 34974
rect 32958 35026 33010 35038
rect 38994 34974 39006 35026
rect 39058 34974 39070 35026
rect 42130 34974 42142 35026
rect 42194 34974 42206 35026
rect 49634 34974 49646 35026
rect 49698 34974 49710 35026
rect 56914 34974 56926 35026
rect 56978 34974 56990 35026
rect 32958 34962 33010 34974
rect 3502 34914 3554 34926
rect 2818 34862 2830 34914
rect 2882 34862 2894 34914
rect 3502 34850 3554 34862
rect 5070 34914 5122 34926
rect 5070 34850 5122 34862
rect 6302 34914 6354 34926
rect 6302 34850 6354 34862
rect 7870 34914 7922 34926
rect 7870 34850 7922 34862
rect 8094 34914 8146 34926
rect 8094 34850 8146 34862
rect 10110 34914 10162 34926
rect 11342 34914 11394 34926
rect 16942 34914 16994 34926
rect 23214 34914 23266 34926
rect 10658 34862 10670 34914
rect 10722 34862 10734 34914
rect 11778 34862 11790 34914
rect 11842 34862 11854 34914
rect 13682 34862 13694 34914
rect 13746 34862 13758 34914
rect 14802 34862 14814 34914
rect 14866 34862 14878 34914
rect 20514 34862 20526 34914
rect 20578 34862 20590 34914
rect 10110 34850 10162 34862
rect 11342 34850 11394 34862
rect 16942 34850 16994 34862
rect 23214 34850 23266 34862
rect 23774 34914 23826 34926
rect 27806 34914 27858 34926
rect 27346 34862 27358 34914
rect 27410 34862 27422 34914
rect 23774 34850 23826 34862
rect 27806 34850 27858 34862
rect 32510 34914 32562 34926
rect 55358 34914 55410 34926
rect 36082 34862 36094 34914
rect 36146 34862 36158 34914
rect 37762 34862 37774 34914
rect 37826 34862 37838 34914
rect 38546 34862 38558 34914
rect 38610 34862 38622 34914
rect 39218 34862 39230 34914
rect 39282 34862 39294 34914
rect 40562 34862 40574 34914
rect 40626 34862 40638 34914
rect 42018 34862 42030 34914
rect 42082 34862 42094 34914
rect 48514 34862 48526 34914
rect 48578 34862 48590 34914
rect 51650 34862 51662 34914
rect 51714 34862 51726 34914
rect 51986 34862 51998 34914
rect 52050 34862 52062 34914
rect 53778 34862 53790 34914
rect 53842 34862 53854 34914
rect 54450 34862 54462 34914
rect 54514 34862 54526 34914
rect 57026 34862 57038 34914
rect 57090 34862 57102 34914
rect 32510 34850 32562 34862
rect 55358 34850 55410 34862
rect 4510 34802 4562 34814
rect 1922 34750 1934 34802
rect 1986 34750 1998 34802
rect 4510 34738 4562 34750
rect 6078 34802 6130 34814
rect 6078 34738 6130 34750
rect 6638 34802 6690 34814
rect 6638 34738 6690 34750
rect 8430 34802 8482 34814
rect 15822 34802 15874 34814
rect 13794 34750 13806 34802
rect 13858 34750 13870 34802
rect 8430 34738 8482 34750
rect 15822 34738 15874 34750
rect 15934 34802 15986 34814
rect 15934 34738 15986 34750
rect 16046 34802 16098 34814
rect 16046 34738 16098 34750
rect 18846 34802 18898 34814
rect 22430 34802 22482 34814
rect 21970 34750 21982 34802
rect 22034 34750 22046 34802
rect 18846 34738 18898 34750
rect 22430 34738 22482 34750
rect 23886 34802 23938 34814
rect 33630 34802 33682 34814
rect 44382 34802 44434 34814
rect 30034 34750 30046 34802
rect 30098 34750 30110 34802
rect 40674 34750 40686 34802
rect 40738 34750 40750 34802
rect 23886 34738 23938 34750
rect 33630 34738 33682 34750
rect 44382 34738 44434 34750
rect 46062 34802 46114 34814
rect 46062 34738 46114 34750
rect 46398 34802 46450 34814
rect 53454 34802 53506 34814
rect 48626 34750 48638 34802
rect 48690 34750 48702 34802
rect 46398 34738 46450 34750
rect 53454 34738 53506 34750
rect 53566 34802 53618 34814
rect 53566 34738 53618 34750
rect 56590 34802 56642 34814
rect 56590 34738 56642 34750
rect 4062 34690 4114 34702
rect 4062 34626 4114 34638
rect 4734 34690 4786 34702
rect 4734 34626 4786 34638
rect 7758 34690 7810 34702
rect 7758 34626 7810 34638
rect 12910 34690 12962 34702
rect 12910 34626 12962 34638
rect 19294 34690 19346 34702
rect 19294 34626 19346 34638
rect 21646 34690 21698 34702
rect 31838 34690 31890 34702
rect 25106 34638 25118 34690
rect 25170 34638 25182 34690
rect 21646 34626 21698 34638
rect 31838 34626 31890 34638
rect 32398 34690 32450 34702
rect 32398 34626 32450 34638
rect 33742 34690 33794 34702
rect 33742 34626 33794 34638
rect 33966 34690 34018 34702
rect 33966 34626 34018 34638
rect 34414 34690 34466 34702
rect 34414 34626 34466 34638
rect 35646 34690 35698 34702
rect 38782 34690 38834 34702
rect 37538 34638 37550 34690
rect 37602 34638 37614 34690
rect 35646 34626 35698 34638
rect 38782 34626 38834 34638
rect 39006 34690 39058 34702
rect 39006 34626 39058 34638
rect 43934 34690 43986 34702
rect 43934 34626 43986 34638
rect 44830 34690 44882 34702
rect 44830 34626 44882 34638
rect 45502 34690 45554 34702
rect 45502 34626 45554 34638
rect 46846 34690 46898 34702
rect 46846 34626 46898 34638
rect 47294 34690 47346 34702
rect 47294 34626 47346 34638
rect 47742 34690 47794 34702
rect 47742 34626 47794 34638
rect 52446 34690 52498 34702
rect 55694 34690 55746 34702
rect 54674 34638 54686 34690
rect 54738 34638 54750 34690
rect 52446 34626 52498 34638
rect 55694 34626 55746 34638
rect 58046 34690 58098 34702
rect 58046 34626 58098 34638
rect 1344 34522 58576 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 58576 34522
rect 1344 34436 58576 34470
rect 4622 34354 4674 34366
rect 4622 34290 4674 34302
rect 6526 34354 6578 34366
rect 6526 34290 6578 34302
rect 6974 34354 7026 34366
rect 11006 34354 11058 34366
rect 10546 34302 10558 34354
rect 10610 34302 10622 34354
rect 6974 34290 7026 34302
rect 11006 34290 11058 34302
rect 14590 34354 14642 34366
rect 16606 34354 16658 34366
rect 24894 34354 24946 34366
rect 16258 34302 16270 34354
rect 16322 34302 16334 34354
rect 24322 34302 24334 34354
rect 24386 34302 24398 34354
rect 14590 34290 14642 34302
rect 16606 34290 16658 34302
rect 24894 34290 24946 34302
rect 29822 34354 29874 34366
rect 29822 34290 29874 34302
rect 30942 34354 30994 34366
rect 30942 34290 30994 34302
rect 31166 34354 31218 34366
rect 31166 34290 31218 34302
rect 31726 34354 31778 34366
rect 47630 34354 47682 34366
rect 37986 34302 37998 34354
rect 38050 34302 38062 34354
rect 40562 34302 40574 34354
rect 40626 34302 40638 34354
rect 46386 34302 46398 34354
rect 46450 34302 46462 34354
rect 31726 34290 31778 34302
rect 47630 34290 47682 34302
rect 49758 34354 49810 34366
rect 49758 34290 49810 34302
rect 51326 34354 51378 34366
rect 55582 34354 55634 34366
rect 52434 34302 52446 34354
rect 52498 34302 52510 34354
rect 51326 34290 51378 34302
rect 55582 34290 55634 34302
rect 55806 34354 55858 34366
rect 55806 34290 55858 34302
rect 6414 34242 6466 34254
rect 6414 34178 6466 34190
rect 7982 34242 8034 34254
rect 7982 34178 8034 34190
rect 9102 34242 9154 34254
rect 9102 34178 9154 34190
rect 11230 34242 11282 34254
rect 11230 34178 11282 34190
rect 11342 34242 11394 34254
rect 11342 34178 11394 34190
rect 13806 34242 13858 34254
rect 13806 34178 13858 34190
rect 14142 34242 14194 34254
rect 14142 34178 14194 34190
rect 17950 34242 18002 34254
rect 17950 34178 18002 34190
rect 20638 34242 20690 34254
rect 20638 34178 20690 34190
rect 26350 34242 26402 34254
rect 26350 34178 26402 34190
rect 27022 34242 27074 34254
rect 27022 34178 27074 34190
rect 30046 34242 30098 34254
rect 30046 34178 30098 34190
rect 34638 34242 34690 34254
rect 49646 34242 49698 34254
rect 38098 34190 38110 34242
rect 38162 34190 38174 34242
rect 40002 34190 40014 34242
rect 40066 34190 40078 34242
rect 40450 34190 40462 34242
rect 40514 34190 40526 34242
rect 42130 34190 42142 34242
rect 42194 34190 42206 34242
rect 47282 34190 47294 34242
rect 47346 34190 47358 34242
rect 34638 34178 34690 34190
rect 49646 34178 49698 34190
rect 50654 34242 50706 34254
rect 50654 34178 50706 34190
rect 52782 34242 52834 34254
rect 52782 34178 52834 34190
rect 53678 34242 53730 34254
rect 53678 34178 53730 34190
rect 55470 34242 55522 34254
rect 57486 34242 57538 34254
rect 56354 34190 56366 34242
rect 56418 34190 56430 34242
rect 55470 34178 55522 34190
rect 57486 34178 57538 34190
rect 9998 34130 10050 34142
rect 5954 34078 5966 34130
rect 6018 34078 6030 34130
rect 6178 34078 6190 34130
rect 6242 34078 6254 34130
rect 7186 34078 7198 34130
rect 7250 34078 7262 34130
rect 9762 34078 9774 34130
rect 9826 34078 9838 34130
rect 9998 34066 10050 34078
rect 10110 34130 10162 34142
rect 10110 34066 10162 34078
rect 18062 34130 18114 34142
rect 21198 34130 21250 34142
rect 25902 34130 25954 34142
rect 18610 34078 18622 34130
rect 18674 34078 18686 34130
rect 19730 34078 19742 34130
rect 19794 34078 19806 34130
rect 21746 34078 21758 34130
rect 21810 34078 21822 34130
rect 18062 34066 18114 34078
rect 21198 34066 21250 34078
rect 25902 34066 25954 34078
rect 26574 34130 26626 34142
rect 26574 34066 26626 34078
rect 27918 34130 27970 34142
rect 27918 34066 27970 34078
rect 30158 34130 30210 34142
rect 30158 34066 30210 34078
rect 30718 34130 30770 34142
rect 30718 34066 30770 34078
rect 30830 34130 30882 34142
rect 36318 34130 36370 34142
rect 40798 34130 40850 34142
rect 46734 34130 46786 34142
rect 33954 34078 33966 34130
rect 34018 34078 34030 34130
rect 37202 34078 37214 34130
rect 37266 34078 37278 34130
rect 38434 34078 38446 34130
rect 38498 34078 38510 34130
rect 41682 34078 41694 34130
rect 41746 34078 41758 34130
rect 41906 34078 41918 34130
rect 41970 34078 41982 34130
rect 43026 34078 43038 34130
rect 43090 34078 43102 34130
rect 44258 34078 44270 34130
rect 44322 34078 44334 34130
rect 44930 34078 44942 34130
rect 44994 34078 45006 34130
rect 45154 34078 45166 34130
rect 45218 34078 45230 34130
rect 30830 34066 30882 34078
rect 36318 34066 36370 34078
rect 40798 34066 40850 34078
rect 46734 34066 46786 34078
rect 49870 34130 49922 34142
rect 51886 34130 51938 34142
rect 50194 34078 50206 34130
rect 50258 34078 50270 34130
rect 49870 34066 49922 34078
rect 51886 34066 51938 34078
rect 53790 34130 53842 34142
rect 53790 34066 53842 34078
rect 54686 34130 54738 34142
rect 56578 34078 56590 34130
rect 56642 34078 56654 34130
rect 54686 34066 54738 34078
rect 5070 34018 5122 34030
rect 5070 33954 5122 33966
rect 5406 34018 5458 34030
rect 5406 33954 5458 33966
rect 8542 34018 8594 34030
rect 8542 33954 8594 33966
rect 12798 34018 12850 34030
rect 12798 33954 12850 33966
rect 13246 34018 13298 34030
rect 13246 33954 13298 33966
rect 15038 34018 15090 34030
rect 15038 33954 15090 33966
rect 15822 34018 15874 34030
rect 26462 34018 26514 34030
rect 20402 33966 20414 34018
rect 20466 33966 20478 34018
rect 15822 33954 15874 33966
rect 26462 33954 26514 33966
rect 29486 34018 29538 34030
rect 35198 34018 35250 34030
rect 38894 34018 38946 34030
rect 48190 34018 48242 34030
rect 33730 33966 33742 34018
rect 33794 33966 33806 34018
rect 35858 33966 35870 34018
rect 35922 33966 35934 34018
rect 37538 33966 37550 34018
rect 37602 33966 37614 34018
rect 43922 33966 43934 34018
rect 43986 33966 43998 34018
rect 45042 33966 45054 34018
rect 45106 33966 45118 34018
rect 29486 33954 29538 33966
rect 35198 33954 35250 33966
rect 38894 33954 38946 33966
rect 48190 33954 48242 33966
rect 48526 34018 48578 34030
rect 48526 33954 48578 33966
rect 54910 34018 54962 34030
rect 54910 33954 54962 33966
rect 58046 34018 58098 34030
rect 58046 33954 58098 33966
rect 7870 33906 7922 33918
rect 53678 33906 53730 33918
rect 57598 33906 57650 33918
rect 34962 33854 34974 33906
rect 35026 33903 35038 33906
rect 35186 33903 35198 33906
rect 35026 33857 35198 33903
rect 35026 33854 35038 33857
rect 35186 33854 35198 33857
rect 35250 33854 35262 33906
rect 44034 33854 44046 33906
rect 44098 33854 44110 33906
rect 54338 33854 54350 33906
rect 54402 33854 54414 33906
rect 7870 33842 7922 33854
rect 53678 33842 53730 33854
rect 57598 33842 57650 33854
rect 1344 33738 58576 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 58576 33738
rect 1344 33652 58576 33686
rect 26910 33570 26962 33582
rect 51438 33570 51490 33582
rect 4386 33518 4398 33570
rect 4450 33518 4462 33570
rect 27906 33518 27918 33570
rect 27970 33518 27982 33570
rect 37426 33518 37438 33570
rect 37490 33567 37502 33570
rect 37874 33567 37886 33570
rect 37490 33521 37886 33567
rect 37490 33518 37502 33521
rect 37874 33518 37886 33521
rect 37938 33518 37950 33570
rect 26910 33506 26962 33518
rect 51438 33506 51490 33518
rect 15150 33458 15202 33470
rect 8306 33406 8318 33458
rect 8370 33406 8382 33458
rect 15150 33394 15202 33406
rect 17614 33458 17666 33470
rect 17614 33394 17666 33406
rect 22094 33458 22146 33470
rect 22094 33394 22146 33406
rect 22542 33458 22594 33470
rect 22542 33394 22594 33406
rect 27358 33458 27410 33470
rect 27358 33394 27410 33406
rect 29710 33458 29762 33470
rect 29710 33394 29762 33406
rect 34190 33458 34242 33470
rect 34190 33394 34242 33406
rect 36766 33458 36818 33470
rect 36766 33394 36818 33406
rect 37438 33458 37490 33470
rect 37438 33394 37490 33406
rect 40574 33458 40626 33470
rect 50430 33458 50482 33470
rect 48402 33406 48414 33458
rect 48466 33406 48478 33458
rect 40574 33394 40626 33406
rect 50430 33394 50482 33406
rect 51550 33458 51602 33470
rect 56254 33458 56306 33470
rect 54338 33406 54350 33458
rect 54402 33406 54414 33458
rect 51550 33394 51602 33406
rect 56254 33394 56306 33406
rect 4734 33346 4786 33358
rect 7982 33346 8034 33358
rect 4498 33294 4510 33346
rect 4562 33294 4574 33346
rect 5730 33294 5742 33346
rect 5794 33294 5806 33346
rect 6738 33294 6750 33346
rect 6802 33294 6814 33346
rect 4734 33282 4786 33294
rect 7982 33282 8034 33294
rect 9214 33346 9266 33358
rect 27582 33346 27634 33358
rect 23650 33294 23662 33346
rect 23714 33294 23726 33346
rect 9214 33282 9266 33294
rect 27582 33282 27634 33294
rect 28478 33346 28530 33358
rect 28478 33282 28530 33294
rect 29934 33346 29986 33358
rect 29934 33282 29986 33294
rect 31950 33346 32002 33358
rect 31950 33282 32002 33294
rect 32510 33346 32562 33358
rect 32510 33282 32562 33294
rect 33294 33346 33346 33358
rect 36318 33346 36370 33358
rect 33506 33294 33518 33346
rect 33570 33294 33582 33346
rect 33294 33282 33346 33294
rect 36318 33282 36370 33294
rect 39790 33346 39842 33358
rect 41582 33346 41634 33358
rect 40002 33294 40014 33346
rect 40066 33294 40078 33346
rect 39790 33282 39842 33294
rect 41582 33282 41634 33294
rect 44158 33346 44210 33358
rect 50990 33346 51042 33358
rect 47954 33294 47966 33346
rect 48018 33294 48030 33346
rect 48514 33294 48526 33346
rect 48578 33294 48590 33346
rect 44158 33282 44210 33294
rect 50990 33282 51042 33294
rect 53902 33346 53954 33358
rect 53902 33282 53954 33294
rect 54238 33346 54290 33358
rect 54562 33294 54574 33346
rect 54626 33294 54638 33346
rect 54238 33282 54290 33294
rect 8318 33234 8370 33246
rect 12462 33234 12514 33246
rect 28814 33234 28866 33246
rect 5842 33182 5854 33234
rect 5906 33182 5918 33234
rect 7298 33182 7310 33234
rect 7362 33182 7374 33234
rect 8530 33182 8542 33234
rect 8594 33182 8606 33234
rect 23090 33182 23102 33234
rect 23154 33182 23166 33234
rect 23426 33182 23438 33234
rect 23490 33182 23502 33234
rect 24434 33182 24446 33234
rect 24498 33182 24510 33234
rect 8318 33170 8370 33182
rect 12462 33170 12514 33182
rect 28814 33170 28866 33182
rect 39678 33234 39730 33246
rect 39678 33170 39730 33182
rect 41806 33234 41858 33246
rect 41806 33170 41858 33182
rect 41918 33234 41970 33246
rect 45502 33234 45554 33246
rect 42018 33182 42030 33234
rect 42082 33182 42094 33234
rect 41918 33170 41970 33182
rect 45502 33170 45554 33182
rect 47182 33234 47234 33246
rect 55918 33234 55970 33246
rect 49074 33182 49086 33234
rect 49138 33182 49150 33234
rect 47182 33170 47234 33182
rect 55918 33170 55970 33182
rect 57150 33234 57202 33246
rect 57150 33170 57202 33182
rect 8206 33122 8258 33134
rect 7186 33070 7198 33122
rect 7250 33070 7262 33122
rect 8206 33058 8258 33070
rect 9662 33122 9714 33134
rect 9662 33058 9714 33070
rect 12126 33122 12178 33134
rect 12126 33058 12178 33070
rect 12350 33122 12402 33134
rect 12350 33058 12402 33070
rect 12910 33122 12962 33134
rect 14030 33122 14082 33134
rect 13682 33070 13694 33122
rect 13746 33070 13758 33122
rect 12910 33058 12962 33070
rect 14030 33058 14082 33070
rect 16158 33122 16210 33134
rect 16158 33058 16210 33070
rect 16270 33122 16322 33134
rect 16270 33058 16322 33070
rect 16382 33122 16434 33134
rect 16382 33058 16434 33070
rect 16606 33122 16658 33134
rect 16606 33058 16658 33070
rect 17278 33122 17330 33134
rect 17278 33058 17330 33070
rect 19182 33122 19234 33134
rect 19182 33058 19234 33070
rect 19854 33122 19906 33134
rect 19854 33058 19906 33070
rect 20862 33122 20914 33134
rect 30830 33122 30882 33134
rect 30258 33070 30270 33122
rect 30322 33070 30334 33122
rect 20862 33058 20914 33070
rect 30830 33058 30882 33070
rect 32398 33122 32450 33134
rect 32398 33058 32450 33070
rect 32622 33122 32674 33134
rect 32622 33058 32674 33070
rect 34750 33122 34802 33134
rect 34750 33058 34802 33070
rect 35422 33122 35474 33134
rect 35422 33058 35474 33070
rect 35982 33122 36034 33134
rect 35982 33058 36034 33070
rect 37886 33122 37938 33134
rect 37886 33058 37938 33070
rect 38446 33122 38498 33134
rect 40910 33122 40962 33134
rect 39218 33070 39230 33122
rect 39282 33070 39294 33122
rect 38446 33058 38498 33070
rect 40910 33058 40962 33070
rect 41694 33122 41746 33134
rect 41694 33058 41746 33070
rect 42926 33122 42978 33134
rect 42926 33058 42978 33070
rect 43262 33122 43314 33134
rect 43262 33058 43314 33070
rect 43710 33122 43762 33134
rect 43710 33058 43762 33070
rect 44606 33122 44658 33134
rect 44606 33058 44658 33070
rect 45614 33122 45666 33134
rect 45614 33058 45666 33070
rect 45726 33122 45778 33134
rect 45726 33058 45778 33070
rect 46398 33122 46450 33134
rect 46398 33058 46450 33070
rect 46734 33122 46786 33134
rect 46734 33058 46786 33070
rect 49534 33122 49586 33134
rect 49534 33058 49586 33070
rect 50318 33122 50370 33134
rect 50318 33058 50370 33070
rect 50542 33122 50594 33134
rect 50542 33058 50594 33070
rect 51662 33122 51714 33134
rect 52670 33122 52722 33134
rect 52322 33070 52334 33122
rect 52386 33070 52398 33122
rect 51662 33058 51714 33070
rect 52670 33058 52722 33070
rect 53342 33122 53394 33134
rect 53342 33058 53394 33070
rect 56142 33122 56194 33134
rect 56142 33058 56194 33070
rect 56366 33122 56418 33134
rect 56366 33058 56418 33070
rect 57486 33122 57538 33134
rect 57486 33058 57538 33070
rect 57934 33122 57986 33134
rect 57934 33058 57986 33070
rect 1344 32954 58576 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 58576 32954
rect 1344 32868 58576 32902
rect 4734 32786 4786 32798
rect 4734 32722 4786 32734
rect 6526 32786 6578 32798
rect 6526 32722 6578 32734
rect 7646 32786 7698 32798
rect 7646 32722 7698 32734
rect 8654 32786 8706 32798
rect 8654 32722 8706 32734
rect 13582 32786 13634 32798
rect 13582 32722 13634 32734
rect 17726 32786 17778 32798
rect 17726 32722 17778 32734
rect 21870 32786 21922 32798
rect 21870 32722 21922 32734
rect 22878 32786 22930 32798
rect 22878 32722 22930 32734
rect 25790 32786 25842 32798
rect 25790 32722 25842 32734
rect 26014 32786 26066 32798
rect 26014 32722 26066 32734
rect 26910 32786 26962 32798
rect 26910 32722 26962 32734
rect 35310 32786 35362 32798
rect 35310 32722 35362 32734
rect 38558 32786 38610 32798
rect 38558 32722 38610 32734
rect 39454 32786 39506 32798
rect 39454 32722 39506 32734
rect 39790 32786 39842 32798
rect 39790 32722 39842 32734
rect 40350 32786 40402 32798
rect 40350 32722 40402 32734
rect 41806 32786 41858 32798
rect 41806 32722 41858 32734
rect 45278 32786 45330 32798
rect 45278 32722 45330 32734
rect 46398 32786 46450 32798
rect 46398 32722 46450 32734
rect 47182 32786 47234 32798
rect 47182 32722 47234 32734
rect 50094 32786 50146 32798
rect 52894 32786 52946 32798
rect 50754 32734 50766 32786
rect 50818 32734 50830 32786
rect 50094 32722 50146 32734
rect 52894 32722 52946 32734
rect 7758 32674 7810 32686
rect 7758 32610 7810 32622
rect 8766 32674 8818 32686
rect 8766 32610 8818 32622
rect 11790 32674 11842 32686
rect 11790 32610 11842 32622
rect 14926 32674 14978 32686
rect 14926 32610 14978 32622
rect 15038 32674 15090 32686
rect 15038 32610 15090 32622
rect 18622 32674 18674 32686
rect 18622 32610 18674 32622
rect 20638 32674 20690 32686
rect 20638 32610 20690 32622
rect 22654 32674 22706 32686
rect 22654 32610 22706 32622
rect 23326 32674 23378 32686
rect 40910 32674 40962 32686
rect 31826 32622 31838 32674
rect 31890 32622 31902 32674
rect 36866 32622 36878 32674
rect 36930 32622 36942 32674
rect 37538 32622 37550 32674
rect 37602 32622 37614 32674
rect 23326 32610 23378 32622
rect 40910 32610 40962 32622
rect 42142 32674 42194 32686
rect 42142 32610 42194 32622
rect 53454 32674 53506 32686
rect 53454 32610 53506 32622
rect 57486 32674 57538 32686
rect 57486 32610 57538 32622
rect 3838 32562 3890 32574
rect 3838 32498 3890 32510
rect 5406 32562 5458 32574
rect 8430 32562 8482 32574
rect 6290 32510 6302 32562
rect 6354 32510 6366 32562
rect 5406 32498 5458 32510
rect 8430 32498 8482 32510
rect 8878 32562 8930 32574
rect 13358 32562 13410 32574
rect 12450 32510 12462 32562
rect 12514 32510 12526 32562
rect 8878 32498 8930 32510
rect 13358 32498 13410 32510
rect 13470 32562 13522 32574
rect 13470 32498 13522 32510
rect 14030 32562 14082 32574
rect 14030 32498 14082 32510
rect 15262 32562 15314 32574
rect 18062 32562 18114 32574
rect 20526 32562 20578 32574
rect 16594 32510 16606 32562
rect 16658 32510 16670 32562
rect 19506 32510 19518 32562
rect 19570 32510 19582 32562
rect 15262 32498 15314 32510
rect 18062 32498 18114 32510
rect 20526 32498 20578 32510
rect 21646 32562 21698 32574
rect 21646 32498 21698 32510
rect 21982 32562 22034 32574
rect 21982 32498 22034 32510
rect 22542 32562 22594 32574
rect 24222 32562 24274 32574
rect 23762 32510 23774 32562
rect 23826 32510 23838 32562
rect 22542 32498 22594 32510
rect 24222 32498 24274 32510
rect 26126 32562 26178 32574
rect 26126 32498 26178 32510
rect 26686 32562 26738 32574
rect 26686 32498 26738 32510
rect 26798 32562 26850 32574
rect 26798 32498 26850 32510
rect 27358 32562 27410 32574
rect 27358 32498 27410 32510
rect 31502 32562 31554 32574
rect 39678 32562 39730 32574
rect 35522 32510 35534 32562
rect 35586 32510 35598 32562
rect 36418 32510 36430 32562
rect 36482 32510 36494 32562
rect 37426 32510 37438 32562
rect 37490 32510 37502 32562
rect 31502 32498 31554 32510
rect 39678 32498 39730 32510
rect 39902 32562 39954 32574
rect 39902 32498 39954 32510
rect 41470 32562 41522 32574
rect 41470 32498 41522 32510
rect 41918 32562 41970 32574
rect 41918 32498 41970 32510
rect 43038 32562 43090 32574
rect 43822 32562 43874 32574
rect 43586 32510 43598 32562
rect 43650 32510 43662 32562
rect 43038 32498 43090 32510
rect 43822 32498 43874 32510
rect 44046 32562 44098 32574
rect 44718 32562 44770 32574
rect 44258 32510 44270 32562
rect 44322 32510 44334 32562
rect 44046 32498 44098 32510
rect 44718 32498 44770 32510
rect 45166 32562 45218 32574
rect 45166 32498 45218 32510
rect 45390 32562 45442 32574
rect 46286 32562 46338 32574
rect 45938 32510 45950 32562
rect 46002 32510 46014 32562
rect 45390 32498 45442 32510
rect 46286 32498 46338 32510
rect 46510 32562 46562 32574
rect 46510 32498 46562 32510
rect 47294 32562 47346 32574
rect 49982 32562 50034 32574
rect 47954 32510 47966 32562
rect 48018 32510 48030 32562
rect 49634 32510 49646 32562
rect 49698 32510 49710 32562
rect 47294 32498 47346 32510
rect 49982 32498 50034 32510
rect 50206 32562 50258 32574
rect 50206 32498 50258 32510
rect 51102 32562 51154 32574
rect 51102 32498 51154 32510
rect 53678 32562 53730 32574
rect 53678 32498 53730 32510
rect 54014 32562 54066 32574
rect 56590 32562 56642 32574
rect 55010 32510 55022 32562
rect 55074 32510 55086 32562
rect 54014 32498 54066 32510
rect 56590 32498 56642 32510
rect 57822 32562 57874 32574
rect 57822 32498 57874 32510
rect 3390 32450 3442 32462
rect 3390 32386 3442 32398
rect 4286 32450 4338 32462
rect 4286 32386 4338 32398
rect 7086 32450 7138 32462
rect 7086 32386 7138 32398
rect 9662 32450 9714 32462
rect 9662 32386 9714 32398
rect 10222 32450 10274 32462
rect 10222 32386 10274 32398
rect 10894 32450 10946 32462
rect 14478 32450 14530 32462
rect 12674 32398 12686 32450
rect 12738 32398 12750 32450
rect 10894 32386 10946 32398
rect 14478 32386 14530 32398
rect 15822 32450 15874 32462
rect 21310 32450 21362 32462
rect 16258 32398 16270 32450
rect 16322 32398 16334 32450
rect 19394 32398 19406 32450
rect 19458 32398 19470 32450
rect 15822 32386 15874 32398
rect 21310 32386 21362 32398
rect 24782 32450 24834 32462
rect 24782 32386 24834 32398
rect 27694 32450 27746 32462
rect 27694 32386 27746 32398
rect 28142 32450 28194 32462
rect 28142 32386 28194 32398
rect 30494 32450 30546 32462
rect 30494 32386 30546 32398
rect 32846 32450 32898 32462
rect 32846 32386 32898 32398
rect 34974 32450 35026 32462
rect 34974 32386 35026 32398
rect 38110 32450 38162 32462
rect 38110 32386 38162 32398
rect 42590 32450 42642 32462
rect 48414 32450 48466 32462
rect 44146 32398 44158 32450
rect 44210 32398 44222 32450
rect 42590 32386 42642 32398
rect 48414 32386 48466 32398
rect 51550 32450 51602 32462
rect 52434 32398 52446 32450
rect 52498 32398 52510 32450
rect 53778 32398 53790 32450
rect 53842 32398 53854 32450
rect 56018 32398 56030 32450
rect 56082 32398 56094 32450
rect 51550 32386 51602 32398
rect 4846 32338 4898 32350
rect 4846 32274 4898 32286
rect 5070 32338 5122 32350
rect 5070 32274 5122 32286
rect 5630 32338 5682 32350
rect 7534 32338 7586 32350
rect 7074 32286 7086 32338
rect 7138 32335 7150 32338
rect 7298 32335 7310 32338
rect 7138 32289 7310 32335
rect 7138 32286 7150 32289
rect 7298 32286 7310 32289
rect 7362 32286 7374 32338
rect 5630 32274 5682 32286
rect 7534 32274 7586 32286
rect 47182 32338 47234 32350
rect 47182 32274 47234 32286
rect 54238 32338 54290 32350
rect 54238 32274 54290 32286
rect 1344 32170 58576 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 58576 32170
rect 1344 32084 58576 32118
rect 14142 32002 14194 32014
rect 14142 31938 14194 31950
rect 14590 32002 14642 32014
rect 44606 32002 44658 32014
rect 22194 31950 22206 32002
rect 22258 31950 22270 32002
rect 23090 31950 23102 32002
rect 23154 31950 23166 32002
rect 48066 31950 48078 32002
rect 48130 31950 48142 32002
rect 14590 31938 14642 31950
rect 44606 31938 44658 31950
rect 6078 31890 6130 31902
rect 6078 31826 6130 31838
rect 8990 31890 9042 31902
rect 8990 31826 9042 31838
rect 10334 31890 10386 31902
rect 10334 31826 10386 31838
rect 11454 31890 11506 31902
rect 13918 31890 13970 31902
rect 12338 31838 12350 31890
rect 12402 31838 12414 31890
rect 11454 31826 11506 31838
rect 13918 31826 13970 31838
rect 15262 31890 15314 31902
rect 17726 31890 17778 31902
rect 16034 31838 16046 31890
rect 16098 31838 16110 31890
rect 15262 31826 15314 31838
rect 17726 31826 17778 31838
rect 20190 31890 20242 31902
rect 20190 31826 20242 31838
rect 20862 31890 20914 31902
rect 20862 31826 20914 31838
rect 21646 31890 21698 31902
rect 34302 31890 34354 31902
rect 33954 31838 33966 31890
rect 34018 31838 34030 31890
rect 21646 31826 21698 31838
rect 34302 31826 34354 31838
rect 36654 31890 36706 31902
rect 40450 31838 40462 31890
rect 40514 31838 40526 31890
rect 46274 31838 46286 31890
rect 46338 31838 46350 31890
rect 46722 31838 46734 31890
rect 46786 31838 46798 31890
rect 48178 31838 48190 31890
rect 48242 31838 48254 31890
rect 53666 31838 53678 31890
rect 53730 31838 53742 31890
rect 55346 31838 55358 31890
rect 55410 31838 55422 31890
rect 56690 31838 56702 31890
rect 56754 31838 56766 31890
rect 36654 31826 36706 31838
rect 8654 31778 8706 31790
rect 8654 31714 8706 31726
rect 8878 31778 8930 31790
rect 8878 31714 8930 31726
rect 9102 31778 9154 31790
rect 9102 31714 9154 31726
rect 9774 31778 9826 31790
rect 13694 31778 13746 31790
rect 18062 31778 18114 31790
rect 12114 31726 12126 31778
rect 12178 31726 12190 31778
rect 15698 31726 15710 31778
rect 15762 31726 15774 31778
rect 9774 31714 9826 31726
rect 13694 31714 13746 31726
rect 18062 31714 18114 31726
rect 21870 31778 21922 31790
rect 21870 31714 21922 31726
rect 23550 31778 23602 31790
rect 23550 31714 23602 31726
rect 23662 31778 23714 31790
rect 34862 31778 34914 31790
rect 24658 31726 24670 31778
rect 24722 31726 24734 31778
rect 33730 31726 33742 31778
rect 33794 31726 33806 31778
rect 23662 31714 23714 31726
rect 34862 31714 34914 31726
rect 35758 31778 35810 31790
rect 35758 31714 35810 31726
rect 37438 31778 37490 31790
rect 37438 31714 37490 31726
rect 39230 31778 39282 31790
rect 41470 31778 41522 31790
rect 43150 31778 43202 31790
rect 39666 31726 39678 31778
rect 39730 31726 39742 31778
rect 42690 31726 42702 31778
rect 42754 31726 42766 31778
rect 39230 31714 39282 31726
rect 41470 31714 41522 31726
rect 43150 31714 43202 31726
rect 44158 31778 44210 31790
rect 44158 31714 44210 31726
rect 44494 31778 44546 31790
rect 51326 31778 51378 31790
rect 46162 31726 46174 31778
rect 46226 31726 46238 31778
rect 46498 31726 46510 31778
rect 46562 31726 46574 31778
rect 47730 31726 47742 31778
rect 47794 31726 47806 31778
rect 48402 31726 48414 31778
rect 48466 31726 48478 31778
rect 49298 31726 49310 31778
rect 49362 31726 49374 31778
rect 44494 31714 44546 31726
rect 51326 31714 51378 31726
rect 51998 31778 52050 31790
rect 51998 31714 52050 31726
rect 52446 31778 52498 31790
rect 52446 31714 52498 31726
rect 52670 31778 52722 31790
rect 52670 31714 52722 31726
rect 54238 31778 54290 31790
rect 57934 31778 57986 31790
rect 54898 31726 54910 31778
rect 54962 31726 54974 31778
rect 55234 31726 55246 31778
rect 55298 31726 55310 31778
rect 56466 31726 56478 31778
rect 56530 31726 56542 31778
rect 57474 31726 57486 31778
rect 57538 31726 57550 31778
rect 54238 31714 54290 31726
rect 57934 31714 57986 31726
rect 4174 31666 4226 31678
rect 4174 31602 4226 31614
rect 7534 31666 7586 31678
rect 7534 31602 7586 31614
rect 18510 31666 18562 31678
rect 18510 31602 18562 31614
rect 20078 31666 20130 31678
rect 20078 31602 20130 31614
rect 23774 31666 23826 31678
rect 23774 31602 23826 31614
rect 24446 31666 24498 31678
rect 31278 31666 31330 31678
rect 26450 31614 26462 31666
rect 26514 31614 26526 31666
rect 24446 31602 24498 31614
rect 31278 31602 31330 31614
rect 35422 31666 35474 31678
rect 35422 31602 35474 31614
rect 37886 31666 37938 31678
rect 37886 31602 37938 31614
rect 38110 31666 38162 31678
rect 38110 31602 38162 31614
rect 44718 31666 44770 31678
rect 50990 31666 51042 31678
rect 49634 31614 49646 31666
rect 49698 31614 49710 31666
rect 50194 31614 50206 31666
rect 50258 31614 50270 31666
rect 44718 31602 44770 31614
rect 50990 31602 51042 31614
rect 53454 31666 53506 31678
rect 53454 31602 53506 31614
rect 53678 31666 53730 31678
rect 56802 31614 56814 31666
rect 56866 31614 56878 31666
rect 53678 31602 53730 31614
rect 2382 31554 2434 31566
rect 2382 31490 2434 31502
rect 2830 31554 2882 31566
rect 2830 31490 2882 31502
rect 3278 31554 3330 31566
rect 3278 31490 3330 31502
rect 3726 31554 3778 31566
rect 3726 31490 3778 31502
rect 4622 31554 4674 31566
rect 4622 31490 4674 31502
rect 5070 31554 5122 31566
rect 5070 31490 5122 31502
rect 5742 31554 5794 31566
rect 5742 31490 5794 31502
rect 6526 31554 6578 31566
rect 6526 31490 6578 31502
rect 6974 31554 7026 31566
rect 6974 31490 7026 31502
rect 10222 31554 10274 31566
rect 10222 31490 10274 31502
rect 10446 31554 10498 31566
rect 10446 31490 10498 31502
rect 10894 31554 10946 31566
rect 10894 31490 10946 31502
rect 13022 31554 13074 31566
rect 13022 31490 13074 31502
rect 19406 31554 19458 31566
rect 19406 31490 19458 31502
rect 20302 31554 20354 31566
rect 20302 31490 20354 31502
rect 28142 31554 28194 31566
rect 28142 31490 28194 31502
rect 30718 31554 30770 31566
rect 30718 31490 30770 31502
rect 31390 31554 31442 31566
rect 31390 31490 31442 31502
rect 35534 31554 35586 31566
rect 35534 31490 35586 31502
rect 36318 31554 36370 31566
rect 36318 31490 36370 31502
rect 36542 31554 36594 31566
rect 36542 31490 36594 31502
rect 36766 31554 36818 31566
rect 36766 31490 36818 31502
rect 37662 31554 37714 31566
rect 37662 31490 37714 31502
rect 38558 31554 38610 31566
rect 38558 31490 38610 31502
rect 40910 31554 40962 31566
rect 40910 31490 40962 31502
rect 42030 31554 42082 31566
rect 42030 31490 42082 31502
rect 44270 31554 44322 31566
rect 52222 31554 52274 31566
rect 49858 31502 49870 31554
rect 49922 31502 49934 31554
rect 44270 31490 44322 31502
rect 52222 31490 52274 31502
rect 1344 31386 58576 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 58576 31386
rect 1344 31300 58576 31334
rect 3726 31218 3778 31230
rect 3726 31154 3778 31166
rect 4622 31218 4674 31230
rect 10894 31218 10946 31230
rect 13134 31218 13186 31230
rect 5058 31166 5070 31218
rect 5122 31166 5134 31218
rect 11890 31166 11902 31218
rect 11954 31166 11966 31218
rect 4622 31154 4674 31166
rect 10894 31154 10946 31166
rect 13134 31154 13186 31166
rect 14702 31218 14754 31230
rect 14702 31154 14754 31166
rect 16494 31218 16546 31230
rect 16494 31154 16546 31166
rect 21646 31218 21698 31230
rect 21646 31154 21698 31166
rect 22430 31218 22482 31230
rect 22430 31154 22482 31166
rect 23662 31218 23714 31230
rect 23662 31154 23714 31166
rect 24782 31218 24834 31230
rect 24782 31154 24834 31166
rect 26014 31218 26066 31230
rect 26014 31154 26066 31166
rect 26126 31218 26178 31230
rect 26126 31154 26178 31166
rect 27358 31218 27410 31230
rect 27358 31154 27410 31166
rect 27582 31218 27634 31230
rect 27582 31154 27634 31166
rect 28254 31218 28306 31230
rect 28254 31154 28306 31166
rect 31950 31218 32002 31230
rect 40910 31218 40962 31230
rect 35746 31166 35758 31218
rect 35810 31166 35822 31218
rect 31950 31154 32002 31166
rect 40910 31154 40962 31166
rect 42926 31218 42978 31230
rect 42926 31154 42978 31166
rect 43038 31218 43090 31230
rect 43038 31154 43090 31166
rect 43822 31218 43874 31230
rect 43822 31154 43874 31166
rect 44830 31218 44882 31230
rect 44830 31154 44882 31166
rect 44942 31218 44994 31230
rect 44942 31154 44994 31166
rect 45054 31218 45106 31230
rect 45054 31154 45106 31166
rect 45838 31218 45890 31230
rect 45838 31154 45890 31166
rect 49422 31218 49474 31230
rect 49422 31154 49474 31166
rect 49758 31218 49810 31230
rect 49758 31154 49810 31166
rect 53118 31218 53170 31230
rect 53118 31154 53170 31166
rect 8318 31106 8370 31118
rect 8318 31042 8370 31054
rect 12686 31106 12738 31118
rect 22766 31106 22818 31118
rect 19394 31054 19406 31106
rect 19458 31054 19470 31106
rect 12686 31042 12738 31054
rect 22766 31042 22818 31054
rect 24894 31106 24946 31118
rect 24894 31042 24946 31054
rect 26238 31106 26290 31118
rect 26238 31042 26290 31054
rect 27694 31106 27746 31118
rect 27694 31042 27746 31054
rect 30382 31106 30434 31118
rect 30382 31042 30434 31054
rect 31166 31106 31218 31118
rect 31166 31042 31218 31054
rect 31502 31106 31554 31118
rect 31502 31042 31554 31054
rect 33630 31106 33682 31118
rect 33630 31042 33682 31054
rect 33966 31106 34018 31118
rect 40798 31106 40850 31118
rect 36530 31054 36542 31106
rect 36594 31054 36606 31106
rect 39778 31054 39790 31106
rect 39842 31054 39854 31106
rect 33966 31042 34018 31054
rect 40798 31042 40850 31054
rect 42814 31106 42866 31118
rect 42814 31042 42866 31054
rect 47070 31106 47122 31118
rect 49534 31106 49586 31118
rect 48626 31054 48638 31106
rect 48690 31054 48702 31106
rect 47070 31042 47122 31054
rect 49534 31042 49586 31054
rect 50878 31106 50930 31118
rect 50878 31042 50930 31054
rect 50990 31106 51042 31118
rect 56366 31106 56418 31118
rect 52322 31054 52334 31106
rect 52386 31054 52398 31106
rect 54786 31054 54798 31106
rect 54850 31054 54862 31106
rect 57474 31054 57486 31106
rect 57538 31054 57550 31106
rect 50990 31042 51042 31054
rect 56366 31042 56418 31054
rect 8094 30994 8146 31006
rect 12238 30994 12290 31006
rect 22318 30994 22370 31006
rect 5282 30942 5294 30994
rect 5346 30942 5358 30994
rect 8530 30942 8542 30994
rect 8594 30942 8606 30994
rect 8754 30942 8766 30994
rect 8818 30942 8830 30994
rect 19842 30942 19854 30994
rect 19906 30942 19918 30994
rect 21522 30942 21534 30994
rect 21586 30942 21598 30994
rect 8094 30930 8146 30942
rect 12238 30930 12290 30942
rect 22318 30930 22370 30942
rect 22542 30994 22594 31006
rect 22542 30930 22594 30942
rect 24558 30994 24610 31006
rect 24558 30930 24610 30942
rect 25566 30994 25618 31006
rect 33854 30994 33906 31006
rect 43934 30994 43986 31006
rect 29922 30942 29934 30994
rect 29986 30942 29998 30994
rect 35634 30942 35646 30994
rect 35698 30942 35710 30994
rect 37874 30942 37886 30994
rect 37938 30942 37950 30994
rect 39666 30942 39678 30994
rect 39730 30942 39742 30994
rect 40338 30942 40350 30994
rect 40402 30942 40414 30994
rect 40562 30942 40574 30994
rect 40626 30942 40638 30994
rect 25566 30930 25618 30942
rect 33854 30930 33906 30942
rect 43934 30930 43986 30942
rect 44158 30994 44210 31006
rect 44158 30930 44210 30942
rect 45502 30994 45554 31006
rect 56702 30994 56754 31006
rect 47506 30942 47518 30994
rect 47570 30942 47582 30994
rect 48290 30942 48302 30994
rect 48354 30942 48366 30994
rect 49970 30942 49982 30994
rect 50034 30942 50046 30994
rect 51650 30942 51662 30994
rect 51714 30942 51726 30994
rect 53666 30942 53678 30994
rect 53730 30942 53742 30994
rect 55346 30942 55358 30994
rect 55410 30942 55422 30994
rect 57698 30942 57710 30994
rect 57762 30942 57774 30994
rect 45502 30930 45554 30942
rect 56702 30930 56754 30942
rect 1934 30882 1986 30894
rect 1934 30818 1986 30830
rect 2270 30882 2322 30894
rect 2270 30818 2322 30830
rect 2830 30882 2882 30894
rect 2830 30818 2882 30830
rect 3166 30882 3218 30894
rect 3166 30818 3218 30830
rect 4174 30882 4226 30894
rect 4174 30818 4226 30830
rect 6190 30882 6242 30894
rect 6190 30818 6242 30830
rect 6638 30882 6690 30894
rect 6638 30818 6690 30830
rect 7086 30882 7138 30894
rect 7086 30818 7138 30830
rect 7534 30882 7586 30894
rect 9662 30882 9714 30894
rect 8418 30830 8430 30882
rect 8482 30830 8494 30882
rect 7534 30818 7586 30830
rect 9662 30818 9714 30830
rect 10558 30882 10610 30894
rect 10558 30818 10610 30830
rect 11454 30882 11506 30894
rect 11454 30818 11506 30830
rect 13918 30882 13970 30894
rect 13918 30818 13970 30830
rect 14366 30882 14418 30894
rect 14366 30818 14418 30830
rect 15262 30882 15314 30894
rect 15262 30818 15314 30830
rect 16046 30882 16098 30894
rect 16046 30818 16098 30830
rect 16942 30882 16994 30894
rect 16942 30818 16994 30830
rect 17726 30882 17778 30894
rect 17726 30818 17778 30830
rect 18398 30882 18450 30894
rect 18398 30818 18450 30830
rect 18846 30882 18898 30894
rect 18846 30818 18898 30830
rect 24110 30882 24162 30894
rect 34190 30882 34242 30894
rect 30146 30830 30158 30882
rect 30210 30830 30222 30882
rect 24110 30818 24162 30830
rect 34190 30818 34242 30830
rect 34974 30882 35026 30894
rect 34974 30818 35026 30830
rect 41470 30882 41522 30894
rect 41470 30818 41522 30830
rect 42590 30882 42642 30894
rect 42590 30818 42642 30830
rect 46286 30882 46338 30894
rect 46286 30818 46338 30830
rect 34414 30770 34466 30782
rect 1922 30718 1934 30770
rect 1986 30767 1998 30770
rect 2818 30767 2830 30770
rect 1986 30721 2830 30767
rect 1986 30718 1998 30721
rect 2818 30718 2830 30721
rect 2882 30718 2894 30770
rect 13906 30718 13918 30770
rect 13970 30767 13982 30770
rect 14690 30767 14702 30770
rect 13970 30721 14702 30767
rect 13970 30718 13982 30721
rect 14690 30718 14702 30721
rect 14754 30718 14766 30770
rect 18498 30718 18510 30770
rect 18562 30767 18574 30770
rect 18834 30767 18846 30770
rect 18562 30721 18846 30767
rect 18562 30718 18574 30721
rect 18834 30718 18846 30721
rect 18898 30718 18910 30770
rect 23538 30718 23550 30770
rect 23602 30767 23614 30770
rect 23762 30767 23774 30770
rect 23602 30721 23774 30767
rect 23602 30718 23614 30721
rect 23762 30718 23774 30721
rect 23826 30767 23838 30770
rect 24098 30767 24110 30770
rect 23826 30721 24110 30767
rect 23826 30718 23838 30721
rect 24098 30718 24110 30721
rect 24162 30718 24174 30770
rect 34414 30706 34466 30718
rect 42142 30770 42194 30782
rect 42142 30706 42194 30718
rect 42366 30770 42418 30782
rect 42366 30706 42418 30718
rect 43822 30770 43874 30782
rect 50878 30770 50930 30782
rect 47394 30718 47406 30770
rect 47458 30718 47470 30770
rect 43822 30706 43874 30718
rect 50878 30706 50930 30718
rect 1344 30602 58576 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 58576 30602
rect 1344 30516 58576 30550
rect 6190 30434 6242 30446
rect 3154 30382 3166 30434
rect 3218 30431 3230 30434
rect 3602 30431 3614 30434
rect 3218 30385 3614 30431
rect 3218 30382 3230 30385
rect 3602 30382 3614 30385
rect 3666 30431 3678 30434
rect 4274 30431 4286 30434
rect 3666 30385 4286 30431
rect 3666 30382 3678 30385
rect 4274 30382 4286 30385
rect 4338 30382 4350 30434
rect 6190 30370 6242 30382
rect 6862 30434 6914 30446
rect 6862 30370 6914 30382
rect 8654 30434 8706 30446
rect 15374 30434 15426 30446
rect 8866 30382 8878 30434
rect 8930 30431 8942 30434
rect 9762 30431 9774 30434
rect 8930 30385 9774 30431
rect 8930 30382 8942 30385
rect 9762 30382 9774 30385
rect 9826 30382 9838 30434
rect 8654 30370 8706 30382
rect 15374 30370 15426 30382
rect 15710 30434 15762 30446
rect 15710 30370 15762 30382
rect 21758 30434 21810 30446
rect 21758 30370 21810 30382
rect 22094 30434 22146 30446
rect 29710 30434 29762 30446
rect 24322 30382 24334 30434
rect 24386 30382 24398 30434
rect 22094 30370 22146 30382
rect 29710 30370 29762 30382
rect 31502 30434 31554 30446
rect 52558 30434 52610 30446
rect 44594 30382 44606 30434
rect 44658 30382 44670 30434
rect 47282 30382 47294 30434
rect 47346 30382 47358 30434
rect 51314 30382 51326 30434
rect 51378 30382 51390 30434
rect 31502 30370 31554 30382
rect 52558 30370 52610 30382
rect 5742 30322 5794 30334
rect 5742 30258 5794 30270
rect 5966 30322 6018 30334
rect 5966 30258 6018 30270
rect 8318 30322 8370 30334
rect 25342 30322 25394 30334
rect 44270 30322 44322 30334
rect 17714 30270 17726 30322
rect 17778 30270 17790 30322
rect 23650 30270 23662 30322
rect 23714 30270 23726 30322
rect 24210 30270 24222 30322
rect 24274 30270 24286 30322
rect 40226 30270 40238 30322
rect 40290 30270 40302 30322
rect 51202 30270 51214 30322
rect 51266 30270 51278 30322
rect 56914 30270 56926 30322
rect 56978 30270 56990 30322
rect 8318 30258 8370 30270
rect 25342 30258 25394 30270
rect 44270 30258 44322 30270
rect 2382 30210 2434 30222
rect 2382 30146 2434 30158
rect 6414 30210 6466 30222
rect 6414 30146 6466 30158
rect 9102 30210 9154 30222
rect 9102 30146 9154 30158
rect 11678 30210 11730 30222
rect 11678 30146 11730 30158
rect 13918 30210 13970 30222
rect 13918 30146 13970 30158
rect 19742 30210 19794 30222
rect 19742 30146 19794 30158
rect 20078 30210 20130 30222
rect 28142 30210 28194 30222
rect 20626 30158 20638 30210
rect 20690 30158 20702 30210
rect 23202 30158 23214 30210
rect 23266 30158 23278 30210
rect 24434 30158 24446 30210
rect 24498 30158 24510 30210
rect 20078 30146 20130 30158
rect 28142 30146 28194 30158
rect 30942 30210 30994 30222
rect 32286 30210 32338 30222
rect 35086 30210 35138 30222
rect 42030 30210 42082 30222
rect 31490 30158 31502 30210
rect 31554 30158 31566 30210
rect 34738 30158 34750 30210
rect 34802 30158 34814 30210
rect 38994 30158 39006 30210
rect 39058 30158 39070 30210
rect 40450 30158 40462 30210
rect 40514 30158 40526 30210
rect 30942 30146 30994 30158
rect 32286 30146 32338 30158
rect 35086 30146 35138 30158
rect 42030 30146 42082 30158
rect 44046 30210 44098 30222
rect 44046 30146 44098 30158
rect 45726 30210 45778 30222
rect 45726 30146 45778 30158
rect 46174 30210 46226 30222
rect 46174 30146 46226 30158
rect 47406 30210 47458 30222
rect 52446 30210 52498 30222
rect 49410 30158 49422 30210
rect 49474 30158 49486 30210
rect 47406 30146 47458 30158
rect 52446 30146 52498 30158
rect 53790 30210 53842 30222
rect 53790 30146 53842 30158
rect 54238 30210 54290 30222
rect 54238 30146 54290 30158
rect 54686 30210 54738 30222
rect 56690 30158 56702 30210
rect 56754 30158 56766 30210
rect 57362 30158 57374 30210
rect 57426 30158 57438 30210
rect 54686 30146 54738 30158
rect 3726 30098 3778 30110
rect 3726 30034 3778 30046
rect 8094 30098 8146 30110
rect 8094 30034 8146 30046
rect 11006 30098 11058 30110
rect 11006 30034 11058 30046
rect 11118 30098 11170 30110
rect 11118 30034 11170 30046
rect 14142 30098 14194 30110
rect 14142 30034 14194 30046
rect 14366 30098 14418 30110
rect 14366 30034 14418 30046
rect 14590 30098 14642 30110
rect 14590 30034 14642 30046
rect 15150 30098 15202 30110
rect 15150 30034 15202 30046
rect 18734 30098 18786 30110
rect 18734 30034 18786 30046
rect 19294 30098 19346 30110
rect 21982 30098 22034 30110
rect 20850 30046 20862 30098
rect 20914 30046 20926 30098
rect 19294 30034 19346 30046
rect 21982 30034 22034 30046
rect 28702 30098 28754 30110
rect 28702 30034 28754 30046
rect 28814 30098 28866 30110
rect 28814 30034 28866 30046
rect 29598 30098 29650 30110
rect 29598 30034 29650 30046
rect 30830 30098 30882 30110
rect 31838 30098 31890 30110
rect 31154 30046 31166 30098
rect 31218 30095 31230 30098
rect 31378 30095 31390 30098
rect 31218 30049 31390 30095
rect 31218 30046 31230 30049
rect 31378 30046 31390 30049
rect 31442 30046 31454 30098
rect 30830 30034 30882 30046
rect 31838 30034 31890 30046
rect 34190 30098 34242 30110
rect 34190 30034 34242 30046
rect 35646 30098 35698 30110
rect 35646 30034 35698 30046
rect 37886 30098 37938 30110
rect 41246 30098 41298 30110
rect 40786 30046 40798 30098
rect 40850 30046 40862 30098
rect 37886 30034 37938 30046
rect 41246 30034 41298 30046
rect 42142 30098 42194 30110
rect 42142 30034 42194 30046
rect 42366 30098 42418 30110
rect 42366 30034 42418 30046
rect 42590 30098 42642 30110
rect 55582 30098 55634 30110
rect 48850 30046 48862 30098
rect 48914 30046 48926 30098
rect 50978 30046 50990 30098
rect 51042 30046 51054 30098
rect 56242 30046 56254 30098
rect 56306 30046 56318 30098
rect 42590 30034 42642 30046
rect 55582 30034 55634 30046
rect 1934 29986 1986 29998
rect 1934 29922 1986 29934
rect 2830 29986 2882 29998
rect 2830 29922 2882 29934
rect 3278 29986 3330 29998
rect 3278 29922 3330 29934
rect 4174 29986 4226 29998
rect 4174 29922 4226 29934
rect 4622 29986 4674 29998
rect 4622 29922 4674 29934
rect 5070 29986 5122 29998
rect 5070 29922 5122 29934
rect 7646 29986 7698 29998
rect 7646 29922 7698 29934
rect 9550 29986 9602 29998
rect 9550 29922 9602 29934
rect 10110 29986 10162 29998
rect 10110 29922 10162 29934
rect 10446 29986 10498 29998
rect 10446 29922 10498 29934
rect 11342 29986 11394 29998
rect 11342 29922 11394 29934
rect 12462 29986 12514 29998
rect 12462 29922 12514 29934
rect 12686 29986 12738 29998
rect 12686 29922 12738 29934
rect 12798 29986 12850 29998
rect 12798 29922 12850 29934
rect 12910 29986 12962 29998
rect 12910 29922 12962 29934
rect 16270 29986 16322 29998
rect 16270 29922 16322 29934
rect 16830 29986 16882 29998
rect 16830 29922 16882 29934
rect 17278 29986 17330 29998
rect 17278 29922 17330 29934
rect 18398 29986 18450 29998
rect 18398 29922 18450 29934
rect 19854 29986 19906 29998
rect 19854 29922 19906 29934
rect 25902 29986 25954 29998
rect 25902 29922 25954 29934
rect 26238 29986 26290 29998
rect 26238 29922 26290 29934
rect 28478 29986 28530 29998
rect 28478 29922 28530 29934
rect 29710 29986 29762 29998
rect 29710 29922 29762 29934
rect 30494 29986 30546 29998
rect 30494 29922 30546 29934
rect 30718 29986 30770 29998
rect 37550 29986 37602 29998
rect 33170 29934 33182 29986
rect 33234 29934 33246 29986
rect 30718 29922 30770 29934
rect 37550 29922 37602 29934
rect 43038 29986 43090 29998
rect 43038 29922 43090 29934
rect 43486 29986 43538 29998
rect 43486 29922 43538 29934
rect 45390 29986 45442 29998
rect 45390 29922 45442 29934
rect 45614 29986 45666 29998
rect 45614 29922 45666 29934
rect 46622 29986 46674 29998
rect 46622 29922 46674 29934
rect 50206 29986 50258 29998
rect 50206 29922 50258 29934
rect 53342 29986 53394 29998
rect 53342 29922 53394 29934
rect 55134 29986 55186 29998
rect 55134 29922 55186 29934
rect 57822 29986 57874 29998
rect 57822 29922 57874 29934
rect 1344 29818 58576 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 58576 29818
rect 1344 29732 58576 29766
rect 2158 29650 2210 29662
rect 2158 29586 2210 29598
rect 2494 29650 2546 29662
rect 2494 29586 2546 29598
rect 2942 29650 2994 29662
rect 7646 29650 7698 29662
rect 5282 29598 5294 29650
rect 5346 29598 5358 29650
rect 2942 29586 2994 29598
rect 7646 29586 7698 29598
rect 8430 29650 8482 29662
rect 8430 29586 8482 29598
rect 8542 29650 8594 29662
rect 8542 29586 8594 29598
rect 8654 29650 8706 29662
rect 8654 29586 8706 29598
rect 18062 29650 18114 29662
rect 18062 29586 18114 29598
rect 20974 29650 21026 29662
rect 20974 29586 21026 29598
rect 21870 29650 21922 29662
rect 21870 29586 21922 29598
rect 26126 29650 26178 29662
rect 26126 29586 26178 29598
rect 26238 29650 26290 29662
rect 26238 29586 26290 29598
rect 29486 29650 29538 29662
rect 29486 29586 29538 29598
rect 32846 29650 32898 29662
rect 32846 29586 32898 29598
rect 33518 29650 33570 29662
rect 33518 29586 33570 29598
rect 35198 29650 35250 29662
rect 35198 29586 35250 29598
rect 38334 29650 38386 29662
rect 38334 29586 38386 29598
rect 38446 29650 38498 29662
rect 38446 29586 38498 29598
rect 39342 29650 39394 29662
rect 39342 29586 39394 29598
rect 44718 29650 44770 29662
rect 44718 29586 44770 29598
rect 47966 29650 48018 29662
rect 47966 29586 48018 29598
rect 54238 29650 54290 29662
rect 54238 29586 54290 29598
rect 55022 29650 55074 29662
rect 55022 29586 55074 29598
rect 56366 29650 56418 29662
rect 57474 29598 57486 29650
rect 57538 29598 57550 29650
rect 56366 29586 56418 29598
rect 4846 29538 4898 29550
rect 4846 29474 4898 29486
rect 7534 29538 7586 29550
rect 16830 29538 16882 29550
rect 22654 29538 22706 29550
rect 27582 29538 27634 29550
rect 11666 29486 11678 29538
rect 11730 29486 11742 29538
rect 13570 29486 13582 29538
rect 13634 29486 13646 29538
rect 20178 29486 20190 29538
rect 20242 29486 20254 29538
rect 23762 29486 23774 29538
rect 23826 29486 23838 29538
rect 7534 29474 7586 29486
rect 16830 29474 16882 29486
rect 22654 29474 22706 29486
rect 27582 29474 27634 29486
rect 29374 29538 29426 29550
rect 37998 29538 38050 29550
rect 30258 29486 30270 29538
rect 30322 29486 30334 29538
rect 32498 29486 32510 29538
rect 32562 29486 32574 29538
rect 29374 29474 29426 29486
rect 37998 29474 38050 29486
rect 38222 29538 38274 29550
rect 38222 29474 38274 29486
rect 39006 29538 39058 29550
rect 39006 29474 39058 29486
rect 41582 29538 41634 29550
rect 48078 29538 48130 29550
rect 44034 29486 44046 29538
rect 44098 29486 44110 29538
rect 46386 29486 46398 29538
rect 46450 29486 46462 29538
rect 41582 29474 41634 29486
rect 48078 29474 48130 29486
rect 50878 29538 50930 29550
rect 53554 29486 53566 29538
rect 53618 29486 53630 29538
rect 50878 29474 50930 29486
rect 5630 29426 5682 29438
rect 5630 29362 5682 29374
rect 6974 29426 7026 29438
rect 9102 29426 9154 29438
rect 14254 29426 14306 29438
rect 16270 29426 16322 29438
rect 7298 29374 7310 29426
rect 7362 29374 7374 29426
rect 10434 29374 10446 29426
rect 10498 29374 10510 29426
rect 11554 29374 11566 29426
rect 11618 29374 11630 29426
rect 13458 29374 13470 29426
rect 13522 29374 13534 29426
rect 15698 29374 15710 29426
rect 15762 29374 15774 29426
rect 6974 29362 7026 29374
rect 9102 29362 9154 29374
rect 14254 29362 14306 29374
rect 16270 29362 16322 29374
rect 18622 29426 18674 29438
rect 18622 29362 18674 29374
rect 19630 29426 19682 29438
rect 25566 29426 25618 29438
rect 20402 29374 20414 29426
rect 20466 29374 20478 29426
rect 23538 29374 23550 29426
rect 23602 29374 23614 29426
rect 24322 29374 24334 29426
rect 24386 29374 24398 29426
rect 19630 29362 19682 29374
rect 25566 29362 25618 29374
rect 26014 29426 26066 29438
rect 26014 29362 26066 29374
rect 26686 29426 26738 29438
rect 39342 29426 39394 29438
rect 27346 29374 27358 29426
rect 27410 29374 27422 29426
rect 30706 29374 30718 29426
rect 30770 29374 30782 29426
rect 31042 29374 31054 29426
rect 31106 29374 31118 29426
rect 34626 29374 34638 29426
rect 34690 29374 34702 29426
rect 36306 29374 36318 29426
rect 36370 29374 36382 29426
rect 36866 29374 36878 29426
rect 36930 29374 36942 29426
rect 26686 29362 26738 29374
rect 39342 29362 39394 29374
rect 39678 29426 39730 29438
rect 39678 29362 39730 29374
rect 40126 29426 40178 29438
rect 40126 29362 40178 29374
rect 40350 29426 40402 29438
rect 40350 29362 40402 29374
rect 40798 29426 40850 29438
rect 40798 29362 40850 29374
rect 41918 29426 41970 29438
rect 48750 29426 48802 29438
rect 54910 29426 54962 29438
rect 43362 29374 43374 29426
rect 43426 29374 43438 29426
rect 44930 29374 44942 29426
rect 44994 29374 45006 29426
rect 46946 29374 46958 29426
rect 47010 29374 47022 29426
rect 49746 29374 49758 29426
rect 49810 29374 49822 29426
rect 53218 29374 53230 29426
rect 53282 29374 53294 29426
rect 41918 29362 41970 29374
rect 48750 29362 48802 29374
rect 54910 29362 54962 29374
rect 55134 29426 55186 29438
rect 55134 29362 55186 29374
rect 56030 29426 56082 29438
rect 56030 29362 56082 29374
rect 56478 29426 56530 29438
rect 56478 29362 56530 29374
rect 56702 29426 56754 29438
rect 57698 29374 57710 29426
rect 57762 29374 57774 29426
rect 56702 29362 56754 29374
rect 3502 29314 3554 29326
rect 3502 29250 3554 29262
rect 3950 29314 4002 29326
rect 3950 29250 4002 29262
rect 4398 29314 4450 29326
rect 4398 29250 4450 29262
rect 5854 29314 5906 29326
rect 5854 29250 5906 29262
rect 6526 29314 6578 29326
rect 6526 29250 6578 29262
rect 9998 29314 10050 29326
rect 9998 29250 10050 29262
rect 11006 29314 11058 29326
rect 11006 29250 11058 29262
rect 19182 29314 19234 29326
rect 19182 29250 19234 29262
rect 21534 29314 21586 29326
rect 21534 29250 21586 29262
rect 22430 29314 22482 29326
rect 23998 29314 24050 29326
rect 22754 29262 22766 29314
rect 22818 29262 22830 29314
rect 22430 29250 22482 29262
rect 23998 29250 24050 29262
rect 24110 29314 24162 29326
rect 24110 29250 24162 29262
rect 28030 29314 28082 29326
rect 31726 29314 31778 29326
rect 40238 29314 40290 29326
rect 30818 29262 30830 29314
rect 30882 29262 30894 29314
rect 34290 29262 34302 29314
rect 34354 29262 34366 29314
rect 36978 29262 36990 29314
rect 37042 29262 37054 29314
rect 28030 29250 28082 29262
rect 31726 29250 31778 29262
rect 40238 29250 40290 29262
rect 42366 29314 42418 29326
rect 42366 29250 42418 29262
rect 48638 29314 48690 29326
rect 48638 29250 48690 29262
rect 49982 29314 50034 29326
rect 55358 29314 55410 29326
rect 52322 29262 52334 29314
rect 52386 29262 52398 29314
rect 49982 29250 50034 29262
rect 55358 29250 55410 29262
rect 10782 29202 10834 29214
rect 10782 29138 10834 29150
rect 29598 29202 29650 29214
rect 29598 29138 29650 29150
rect 36094 29202 36146 29214
rect 36094 29138 36146 29150
rect 47966 29202 48018 29214
rect 47966 29138 48018 29150
rect 50094 29202 50146 29214
rect 50094 29138 50146 29150
rect 50990 29202 51042 29214
rect 50990 29138 51042 29150
rect 51214 29202 51266 29214
rect 51214 29138 51266 29150
rect 51326 29202 51378 29214
rect 51326 29138 51378 29150
rect 55582 29202 55634 29214
rect 55582 29138 55634 29150
rect 1344 29034 58576 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 58576 29034
rect 1344 28948 58576 28982
rect 5854 28866 5906 28878
rect 17950 28866 18002 28878
rect 24670 28866 24722 28878
rect 7746 28814 7758 28866
rect 7810 28814 7822 28866
rect 11218 28814 11230 28866
rect 11282 28814 11294 28866
rect 22194 28814 22206 28866
rect 22258 28863 22270 28866
rect 22754 28863 22766 28866
rect 22258 28817 22766 28863
rect 22258 28814 22270 28817
rect 22754 28814 22766 28817
rect 22818 28814 22830 28866
rect 24098 28814 24110 28866
rect 24162 28814 24174 28866
rect 5854 28802 5906 28814
rect 17950 28802 18002 28814
rect 24670 28802 24722 28814
rect 31278 28866 31330 28878
rect 47394 28814 47406 28866
rect 47458 28814 47470 28866
rect 49410 28814 49422 28866
rect 49474 28814 49486 28866
rect 31278 28802 31330 28814
rect 3726 28754 3778 28766
rect 3726 28690 3778 28702
rect 4174 28754 4226 28766
rect 4174 28690 4226 28702
rect 4622 28754 4674 28766
rect 4622 28690 4674 28702
rect 5070 28754 5122 28766
rect 5070 28690 5122 28702
rect 5966 28754 6018 28766
rect 12910 28754 12962 28766
rect 10882 28702 10894 28754
rect 10946 28702 10958 28754
rect 5966 28690 6018 28702
rect 12910 28690 12962 28702
rect 13806 28754 13858 28766
rect 21758 28754 21810 28766
rect 19394 28702 19406 28754
rect 19458 28702 19470 28754
rect 13806 28690 13858 28702
rect 21758 28690 21810 28702
rect 23774 28754 23826 28766
rect 23774 28690 23826 28702
rect 24782 28754 24834 28766
rect 24782 28690 24834 28702
rect 28702 28754 28754 28766
rect 28702 28690 28754 28702
rect 32286 28754 32338 28766
rect 33966 28754 34018 28766
rect 38894 28754 38946 28766
rect 33058 28702 33070 28754
rect 33122 28702 33134 28754
rect 34962 28702 34974 28754
rect 35026 28702 35038 28754
rect 37538 28702 37550 28754
rect 37602 28702 37614 28754
rect 32286 28690 32338 28702
rect 33966 28690 34018 28702
rect 38894 28690 38946 28702
rect 39230 28754 39282 28766
rect 39230 28690 39282 28702
rect 45390 28754 45442 28766
rect 53678 28754 53730 28766
rect 47058 28702 47070 28754
rect 47122 28702 47134 28754
rect 48962 28702 48974 28754
rect 49026 28702 49038 28754
rect 45390 28690 45442 28702
rect 53678 28690 53730 28702
rect 56142 28754 56194 28766
rect 56142 28690 56194 28702
rect 7086 28642 7138 28654
rect 2930 28590 2942 28642
rect 2994 28590 3006 28642
rect 7086 28578 7138 28590
rect 7310 28642 7362 28654
rect 7310 28578 7362 28590
rect 8654 28642 8706 28654
rect 16270 28642 16322 28654
rect 20974 28642 21026 28654
rect 9314 28590 9326 28642
rect 9378 28590 9390 28642
rect 11218 28590 11230 28642
rect 11282 28590 11294 28642
rect 14018 28590 14030 28642
rect 14082 28590 14094 28642
rect 14242 28590 14254 28642
rect 14306 28590 14318 28642
rect 16818 28590 16830 28642
rect 16882 28590 16894 28642
rect 17266 28590 17278 28642
rect 17330 28590 17342 28642
rect 18162 28590 18174 28642
rect 18226 28590 18238 28642
rect 18498 28590 18510 28642
rect 18562 28590 18574 28642
rect 19282 28590 19294 28642
rect 19346 28590 19358 28642
rect 8654 28578 8706 28590
rect 16270 28578 16322 28590
rect 20974 28578 21026 28590
rect 22206 28642 22258 28654
rect 22206 28578 22258 28590
rect 22654 28642 22706 28654
rect 22654 28578 22706 28590
rect 23102 28642 23154 28654
rect 23102 28578 23154 28590
rect 23550 28642 23602 28654
rect 23550 28578 23602 28590
rect 26686 28642 26738 28654
rect 26686 28578 26738 28590
rect 27918 28642 27970 28654
rect 27918 28578 27970 28590
rect 30606 28642 30658 28654
rect 35534 28642 35586 28654
rect 33506 28590 33518 28642
rect 33570 28590 33582 28642
rect 30606 28578 30658 28590
rect 35534 28578 35586 28590
rect 35870 28642 35922 28654
rect 35870 28578 35922 28590
rect 36430 28642 36482 28654
rect 36430 28578 36482 28590
rect 39678 28642 39730 28654
rect 52334 28642 52386 28654
rect 40674 28590 40686 28642
rect 40738 28590 40750 28642
rect 42802 28590 42814 28642
rect 42866 28590 42878 28642
rect 44370 28590 44382 28642
rect 44434 28590 44446 28642
rect 46498 28590 46510 28642
rect 46562 28590 46574 28642
rect 47506 28590 47518 28642
rect 47570 28590 47582 28642
rect 48626 28590 48638 28642
rect 48690 28590 48702 28642
rect 49522 28590 49534 28642
rect 49586 28590 49598 28642
rect 39678 28578 39730 28590
rect 52334 28578 52386 28590
rect 52558 28642 52610 28654
rect 52558 28578 52610 28590
rect 54014 28642 54066 28654
rect 54014 28578 54066 28590
rect 54238 28642 54290 28654
rect 54238 28578 54290 28590
rect 56030 28642 56082 28654
rect 56030 28578 56082 28590
rect 56702 28642 56754 28654
rect 56702 28578 56754 28590
rect 57710 28642 57762 28654
rect 57710 28578 57762 28590
rect 7198 28530 7250 28542
rect 15598 28530 15650 28542
rect 1922 28478 1934 28530
rect 1986 28478 1998 28530
rect 9986 28478 9998 28530
rect 10050 28478 10062 28530
rect 7198 28466 7250 28478
rect 15598 28466 15650 28478
rect 15822 28530 15874 28542
rect 24894 28530 24946 28542
rect 19730 28478 19742 28530
rect 19794 28478 19806 28530
rect 15822 28466 15874 28478
rect 24894 28466 24946 28478
rect 26350 28530 26402 28542
rect 26350 28466 26402 28478
rect 27358 28530 27410 28542
rect 27358 28466 27410 28478
rect 30270 28530 30322 28542
rect 30270 28466 30322 28478
rect 31278 28530 31330 28542
rect 31278 28466 31330 28478
rect 31390 28530 31442 28542
rect 31390 28466 31442 28478
rect 32174 28530 32226 28542
rect 32174 28466 32226 28478
rect 32398 28530 32450 28542
rect 32398 28466 32450 28478
rect 34526 28530 34578 28542
rect 34526 28466 34578 28478
rect 34750 28530 34802 28542
rect 34750 28466 34802 28478
rect 36766 28530 36818 28542
rect 37998 28530 38050 28542
rect 37762 28478 37774 28530
rect 37826 28478 37838 28530
rect 36766 28466 36818 28478
rect 37998 28466 38050 28478
rect 38334 28530 38386 28542
rect 46062 28530 46114 28542
rect 50654 28530 50706 28542
rect 40562 28478 40574 28530
rect 40626 28478 40638 28530
rect 44706 28478 44718 28530
rect 44770 28478 44782 28530
rect 49858 28478 49870 28530
rect 49922 28478 49934 28530
rect 38334 28466 38386 28478
rect 46062 28466 46114 28478
rect 50654 28466 50706 28478
rect 50990 28530 51042 28542
rect 50990 28466 51042 28478
rect 51214 28530 51266 28542
rect 51214 28466 51266 28478
rect 51774 28530 51826 28542
rect 51774 28466 51826 28478
rect 51998 28530 52050 28542
rect 51998 28466 52050 28478
rect 52110 28530 52162 28542
rect 52110 28466 52162 28478
rect 56254 28530 56306 28542
rect 56254 28466 56306 28478
rect 57150 28530 57202 28542
rect 57150 28466 57202 28478
rect 57374 28530 57426 28542
rect 57374 28466 57426 28478
rect 6078 28418 6130 28430
rect 6078 28354 6130 28366
rect 15710 28418 15762 28430
rect 15710 28354 15762 28366
rect 20526 28418 20578 28430
rect 20526 28354 20578 28366
rect 25902 28418 25954 28430
rect 25902 28354 25954 28366
rect 27134 28418 27186 28430
rect 27134 28354 27186 28366
rect 27246 28418 27298 28430
rect 27246 28354 27298 28366
rect 28254 28418 28306 28430
rect 28254 28354 28306 28366
rect 34974 28418 35026 28430
rect 34974 28354 35026 28366
rect 36654 28418 36706 28430
rect 36654 28354 36706 28366
rect 38110 28418 38162 28430
rect 50878 28418 50930 28430
rect 40786 28366 40798 28418
rect 40850 28366 40862 28418
rect 38110 28354 38162 28366
rect 50878 28354 50930 28366
rect 53566 28418 53618 28430
rect 53566 28354 53618 28366
rect 53790 28418 53842 28430
rect 55470 28418 55522 28430
rect 55122 28366 55134 28418
rect 55186 28366 55198 28418
rect 53790 28354 53842 28366
rect 55470 28354 55522 28366
rect 57598 28418 57650 28430
rect 57598 28354 57650 28366
rect 1344 28250 58576 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 58576 28250
rect 1344 28164 58576 28198
rect 5294 28082 5346 28094
rect 5294 28018 5346 28030
rect 6526 28082 6578 28094
rect 9774 28082 9826 28094
rect 8418 28030 8430 28082
rect 8482 28030 8494 28082
rect 6526 28018 6578 28030
rect 9774 28018 9826 28030
rect 10222 28082 10274 28094
rect 10222 28018 10274 28030
rect 10670 28082 10722 28094
rect 16046 28082 16098 28094
rect 12002 28030 12014 28082
rect 12066 28030 12078 28082
rect 13010 28030 13022 28082
rect 13074 28030 13086 28082
rect 10670 28018 10722 28030
rect 16046 28018 16098 28030
rect 16942 28082 16994 28094
rect 16942 28018 16994 28030
rect 18734 28082 18786 28094
rect 18734 28018 18786 28030
rect 18846 28082 18898 28094
rect 18846 28018 18898 28030
rect 20750 28082 20802 28094
rect 20750 28018 20802 28030
rect 23662 28082 23714 28094
rect 24670 28082 24722 28094
rect 23986 28030 23998 28082
rect 24050 28030 24062 28082
rect 23662 28018 23714 28030
rect 24670 28018 24722 28030
rect 24894 28082 24946 28094
rect 24894 28018 24946 28030
rect 31054 28082 31106 28094
rect 31054 28018 31106 28030
rect 31166 28082 31218 28094
rect 31166 28018 31218 28030
rect 31726 28082 31778 28094
rect 31726 28018 31778 28030
rect 32622 28082 32674 28094
rect 32622 28018 32674 28030
rect 39342 28082 39394 28094
rect 39342 28018 39394 28030
rect 40014 28082 40066 28094
rect 42814 28082 42866 28094
rect 41570 28030 41582 28082
rect 41634 28030 41646 28082
rect 40014 28018 40066 28030
rect 42814 28018 42866 28030
rect 47854 28082 47906 28094
rect 47854 28018 47906 28030
rect 49870 28082 49922 28094
rect 52994 28030 53006 28082
rect 53058 28030 53070 28082
rect 49870 28018 49922 28030
rect 3166 27970 3218 27982
rect 14030 27970 14082 27982
rect 11442 27918 11454 27970
rect 11506 27918 11518 27970
rect 3166 27906 3218 27918
rect 14030 27906 14082 27918
rect 14254 27970 14306 27982
rect 14254 27906 14306 27918
rect 14366 27970 14418 27982
rect 14366 27906 14418 27918
rect 16718 27970 16770 27982
rect 16718 27906 16770 27918
rect 18174 27970 18226 27982
rect 28142 27970 28194 27982
rect 21970 27918 21982 27970
rect 22034 27918 22046 27970
rect 22642 27918 22654 27970
rect 22706 27918 22718 27970
rect 26114 27918 26126 27970
rect 26178 27918 26190 27970
rect 18174 27906 18226 27918
rect 28142 27906 28194 27918
rect 28254 27970 28306 27982
rect 35534 27970 35586 27982
rect 39230 27970 39282 27982
rect 34178 27918 34190 27970
rect 34242 27918 34254 27970
rect 36642 27918 36654 27970
rect 36706 27918 36718 27970
rect 37538 27918 37550 27970
rect 37602 27918 37614 27970
rect 28254 27906 28306 27918
rect 35534 27906 35586 27918
rect 39230 27906 39282 27918
rect 40574 27970 40626 27982
rect 40574 27906 40626 27918
rect 50430 27970 50482 27982
rect 50430 27906 50482 27918
rect 50654 27970 50706 27982
rect 50654 27906 50706 27918
rect 51886 27970 51938 27982
rect 51886 27906 51938 27918
rect 52110 27970 52162 27982
rect 57486 27970 57538 27982
rect 53106 27918 53118 27970
rect 53170 27918 53182 27970
rect 52110 27906 52162 27918
rect 57486 27906 57538 27918
rect 57822 27970 57874 27982
rect 57822 27906 57874 27918
rect 3950 27858 4002 27870
rect 7422 27858 7474 27870
rect 7186 27806 7198 27858
rect 7250 27806 7262 27858
rect 3950 27794 4002 27806
rect 7422 27794 7474 27806
rect 7646 27858 7698 27870
rect 8766 27858 8818 27870
rect 12798 27858 12850 27870
rect 13246 27858 13298 27870
rect 15262 27858 15314 27870
rect 7858 27806 7870 27858
rect 7922 27806 7934 27858
rect 11666 27806 11678 27858
rect 11730 27806 11742 27858
rect 12226 27806 12238 27858
rect 12290 27806 12302 27858
rect 13010 27806 13022 27858
rect 13074 27806 13086 27858
rect 13346 27806 13358 27858
rect 13410 27806 13422 27858
rect 7646 27794 7698 27806
rect 8766 27794 8818 27806
rect 12798 27794 12850 27806
rect 13246 27794 13298 27806
rect 15262 27794 15314 27806
rect 16606 27858 16658 27870
rect 16606 27794 16658 27806
rect 18622 27858 18674 27870
rect 19742 27858 19794 27870
rect 19170 27806 19182 27858
rect 19234 27806 19246 27858
rect 18622 27794 18674 27806
rect 19742 27794 19794 27806
rect 20302 27858 20354 27870
rect 24558 27858 24610 27870
rect 30606 27858 30658 27870
rect 20850 27806 20862 27858
rect 20914 27806 20926 27858
rect 22194 27806 22206 27858
rect 22258 27806 22270 27858
rect 22754 27806 22766 27858
rect 22818 27806 22830 27858
rect 26450 27806 26462 27858
rect 26514 27806 26526 27858
rect 27122 27806 27134 27858
rect 27186 27806 27198 27858
rect 20302 27794 20354 27806
rect 24558 27794 24610 27806
rect 30606 27794 30658 27806
rect 31278 27858 31330 27870
rect 42702 27858 42754 27870
rect 34402 27806 34414 27858
rect 34466 27806 34478 27858
rect 35186 27806 35198 27858
rect 35250 27806 35262 27858
rect 36754 27806 36766 27858
rect 36818 27806 36830 27858
rect 37314 27806 37326 27858
rect 37378 27806 37390 27858
rect 38546 27806 38558 27858
rect 38610 27806 38622 27858
rect 31278 27794 31330 27806
rect 42702 27794 42754 27806
rect 42926 27858 42978 27870
rect 47742 27858 47794 27870
rect 43250 27806 43262 27858
rect 43314 27806 43326 27858
rect 43922 27806 43934 27858
rect 43986 27806 43998 27858
rect 44930 27806 44942 27858
rect 44994 27806 45006 27858
rect 45714 27806 45726 27858
rect 45778 27806 45790 27858
rect 46834 27806 46846 27858
rect 46898 27806 46910 27858
rect 47954 27806 47966 27858
rect 48018 27806 48030 27858
rect 49634 27806 49646 27858
rect 49698 27806 49710 27858
rect 52994 27806 53006 27858
rect 53058 27806 53070 27858
rect 54562 27806 54574 27858
rect 54626 27806 54638 27858
rect 56018 27806 56030 27858
rect 56082 27806 56094 27858
rect 42926 27794 42978 27806
rect 47742 27794 47794 27806
rect 1822 27746 1874 27758
rect 1822 27682 1874 27694
rect 2270 27746 2322 27758
rect 2270 27682 2322 27694
rect 2718 27746 2770 27758
rect 2718 27682 2770 27694
rect 3614 27746 3666 27758
rect 3614 27682 3666 27694
rect 4398 27746 4450 27758
rect 4398 27682 4450 27694
rect 4958 27746 5010 27758
rect 4958 27682 5010 27694
rect 5854 27746 5906 27758
rect 8990 27746 9042 27758
rect 7746 27694 7758 27746
rect 7810 27694 7822 27746
rect 5854 27682 5906 27694
rect 8990 27682 9042 27694
rect 15710 27746 15762 27758
rect 15710 27682 15762 27694
rect 17726 27746 17778 27758
rect 17726 27682 17778 27694
rect 25566 27746 25618 27758
rect 28702 27746 28754 27758
rect 42142 27746 42194 27758
rect 46958 27746 47010 27758
rect 26786 27694 26798 27746
rect 26850 27694 26862 27746
rect 34178 27694 34190 27746
rect 34242 27694 34254 27746
rect 36866 27694 36878 27746
rect 36930 27694 36942 27746
rect 44034 27694 44046 27746
rect 44098 27694 44110 27746
rect 44482 27694 44494 27746
rect 44546 27694 44558 27746
rect 45938 27694 45950 27746
rect 46002 27694 46014 27746
rect 25566 27682 25618 27694
rect 28702 27682 28754 27694
rect 42142 27682 42194 27694
rect 46958 27682 47010 27694
rect 50542 27746 50594 27758
rect 50542 27682 50594 27694
rect 51214 27746 51266 27758
rect 52210 27694 52222 27746
rect 52274 27694 52286 27746
rect 51214 27682 51266 27694
rect 6302 27634 6354 27646
rect 1810 27582 1822 27634
rect 1874 27631 1886 27634
rect 3266 27631 3278 27634
rect 1874 27585 3278 27631
rect 1874 27582 1886 27585
rect 3266 27582 3278 27585
rect 3330 27582 3342 27634
rect 6302 27570 6354 27582
rect 6638 27634 6690 27646
rect 28142 27634 28194 27646
rect 15138 27582 15150 27634
rect 15202 27631 15214 27634
rect 15922 27631 15934 27634
rect 15202 27585 15934 27631
rect 15202 27582 15214 27585
rect 15922 27582 15934 27585
rect 15986 27582 15998 27634
rect 25442 27582 25454 27634
rect 25506 27631 25518 27634
rect 26002 27631 26014 27634
rect 25506 27585 26014 27631
rect 25506 27582 25518 27585
rect 26002 27582 26014 27585
rect 26066 27582 26078 27634
rect 6638 27570 6690 27582
rect 28142 27570 28194 27582
rect 39342 27634 39394 27646
rect 39342 27570 39394 27582
rect 41918 27634 41970 27646
rect 41918 27570 41970 27582
rect 1344 27466 58576 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 58576 27466
rect 1344 27380 58576 27414
rect 7198 27298 7250 27310
rect 15150 27298 15202 27310
rect 20638 27298 20690 27310
rect 33854 27298 33906 27310
rect 8082 27246 8094 27298
rect 8146 27295 8158 27298
rect 8306 27295 8318 27298
rect 8146 27249 8318 27295
rect 8146 27246 8158 27249
rect 8306 27246 8318 27249
rect 8370 27246 8382 27298
rect 15922 27246 15934 27298
rect 15986 27295 15998 27298
rect 16258 27295 16270 27298
rect 15986 27249 16270 27295
rect 15986 27246 15998 27249
rect 16258 27246 16270 27249
rect 16322 27246 16334 27298
rect 23762 27246 23774 27298
rect 23826 27246 23838 27298
rect 7198 27234 7250 27246
rect 15150 27234 15202 27246
rect 20638 27234 20690 27246
rect 33854 27234 33906 27246
rect 34190 27298 34242 27310
rect 51886 27298 51938 27310
rect 40674 27246 40686 27298
rect 40738 27246 40750 27298
rect 43362 27246 43374 27298
rect 43426 27246 43438 27298
rect 47842 27246 47854 27298
rect 47906 27295 47918 27298
rect 48290 27295 48302 27298
rect 47906 27249 48302 27295
rect 47906 27246 47918 27249
rect 48290 27246 48302 27249
rect 48354 27246 48366 27298
rect 34190 27234 34242 27246
rect 51886 27234 51938 27246
rect 53566 27298 53618 27310
rect 53566 27234 53618 27246
rect 55806 27298 55858 27310
rect 55806 27234 55858 27246
rect 56142 27298 56194 27310
rect 56142 27234 56194 27246
rect 4958 27186 5010 27198
rect 4958 27122 5010 27134
rect 6190 27186 6242 27198
rect 6190 27122 6242 27134
rect 8094 27186 8146 27198
rect 8094 27122 8146 27134
rect 8430 27186 8482 27198
rect 14926 27186 14978 27198
rect 10322 27134 10334 27186
rect 10386 27134 10398 27186
rect 14578 27134 14590 27186
rect 14642 27134 14654 27186
rect 8430 27122 8482 27134
rect 14926 27122 14978 27134
rect 16830 27186 16882 27198
rect 16830 27122 16882 27134
rect 17950 27186 18002 27198
rect 17950 27122 18002 27134
rect 18846 27186 18898 27198
rect 21646 27186 21698 27198
rect 20066 27134 20078 27186
rect 20130 27134 20142 27186
rect 18846 27122 18898 27134
rect 21646 27122 21698 27134
rect 22094 27186 22146 27198
rect 22094 27122 22146 27134
rect 22654 27186 22706 27198
rect 27694 27186 27746 27198
rect 23538 27134 23550 27186
rect 23602 27134 23614 27186
rect 25666 27134 25678 27186
rect 25730 27134 25742 27186
rect 26562 27134 26574 27186
rect 26626 27134 26638 27186
rect 22654 27122 22706 27134
rect 27694 27122 27746 27134
rect 28142 27186 28194 27198
rect 28142 27122 28194 27134
rect 31502 27186 31554 27198
rect 35198 27186 35250 27198
rect 32274 27134 32286 27186
rect 32338 27134 32350 27186
rect 31502 27122 31554 27134
rect 35198 27122 35250 27134
rect 36094 27186 36146 27198
rect 36094 27122 36146 27134
rect 39118 27186 39170 27198
rect 39118 27122 39170 27134
rect 42254 27186 42306 27198
rect 46398 27186 46450 27198
rect 44258 27134 44270 27186
rect 44322 27134 44334 27186
rect 42254 27122 42306 27134
rect 46398 27122 46450 27134
rect 47294 27186 47346 27198
rect 47294 27122 47346 27134
rect 47854 27186 47906 27198
rect 47854 27122 47906 27134
rect 48302 27186 48354 27198
rect 48302 27122 48354 27134
rect 50766 27186 50818 27198
rect 50766 27122 50818 27134
rect 52334 27186 52386 27198
rect 52334 27122 52386 27134
rect 57934 27186 57986 27198
rect 57934 27122 57986 27134
rect 2606 27074 2658 27086
rect 6078 27074 6130 27086
rect 5730 27022 5742 27074
rect 5794 27022 5806 27074
rect 2606 27010 2658 27022
rect 6078 27010 6130 27022
rect 6302 27074 6354 27086
rect 6302 27010 6354 27022
rect 7310 27074 7362 27086
rect 10446 27074 10498 27086
rect 9874 27022 9886 27074
rect 9938 27022 9950 27074
rect 7310 27010 7362 27022
rect 10446 27010 10498 27022
rect 12350 27074 12402 27086
rect 12350 27010 12402 27022
rect 12574 27074 12626 27086
rect 12574 27010 12626 27022
rect 12910 27074 12962 27086
rect 12910 27010 12962 27022
rect 14702 27074 14754 27086
rect 14702 27010 14754 27022
rect 15374 27074 15426 27086
rect 15374 27010 15426 27022
rect 16718 27074 16770 27086
rect 18510 27074 18562 27086
rect 17154 27022 17166 27074
rect 17218 27022 17230 27074
rect 16718 27010 16770 27022
rect 18510 27010 18562 27022
rect 20190 27074 20242 27086
rect 20862 27074 20914 27086
rect 24334 27074 24386 27086
rect 20290 27022 20302 27074
rect 20354 27022 20366 27074
rect 23314 27022 23326 27074
rect 23378 27022 23390 27074
rect 20190 27010 20242 27022
rect 20862 27010 20914 27022
rect 24334 27010 24386 27022
rect 24782 27074 24834 27086
rect 24782 27010 24834 27022
rect 25006 27074 25058 27086
rect 28590 27074 28642 27086
rect 26114 27022 26126 27074
rect 26178 27022 26190 27074
rect 27010 27022 27022 27074
rect 27074 27022 27086 27074
rect 25006 27010 25058 27022
rect 28590 27010 28642 27022
rect 30158 27074 30210 27086
rect 30158 27010 30210 27022
rect 30494 27074 30546 27086
rect 30494 27010 30546 27022
rect 30942 27074 30994 27086
rect 30942 27010 30994 27022
rect 31166 27074 31218 27086
rect 31166 27010 31218 27022
rect 31390 27074 31442 27086
rect 31390 27010 31442 27022
rect 38446 27074 38498 27086
rect 38446 27010 38498 27022
rect 38782 27074 38834 27086
rect 41694 27074 41746 27086
rect 40226 27022 40238 27074
rect 40290 27022 40302 27074
rect 40674 27022 40686 27074
rect 40738 27022 40750 27074
rect 41458 27022 41470 27074
rect 41522 27022 41534 27074
rect 38782 27010 38834 27022
rect 41694 27010 41746 27022
rect 43374 27074 43426 27086
rect 49982 27074 50034 27086
rect 43698 27022 43710 27074
rect 43762 27022 43774 27074
rect 43374 27010 43426 27022
rect 49982 27010 50034 27022
rect 51550 27074 51602 27086
rect 53678 27074 53730 27086
rect 56030 27074 56082 27086
rect 51874 27022 51886 27074
rect 51938 27022 51950 27074
rect 54338 27022 54350 27074
rect 54402 27022 54414 27074
rect 54898 27022 54910 27074
rect 54962 27022 54974 27074
rect 51550 27010 51602 27022
rect 53678 27010 53730 27022
rect 56030 27010 56082 27022
rect 3502 26962 3554 26974
rect 3502 26898 3554 26910
rect 4398 26962 4450 26974
rect 4398 26898 4450 26910
rect 9326 26962 9378 26974
rect 9326 26898 9378 26910
rect 10334 26962 10386 26974
rect 10334 26898 10386 26910
rect 11118 26962 11170 26974
rect 13806 26962 13858 26974
rect 11442 26910 11454 26962
rect 11506 26910 11518 26962
rect 11118 26898 11170 26910
rect 13806 26898 13858 26910
rect 14478 26962 14530 26974
rect 14478 26898 14530 26910
rect 16942 26962 16994 26974
rect 16942 26898 16994 26910
rect 19294 26962 19346 26974
rect 19294 26898 19346 26910
rect 26574 26962 26626 26974
rect 26574 26898 26626 26910
rect 30270 26962 30322 26974
rect 30270 26898 30322 26910
rect 32398 26962 32450 26974
rect 32398 26898 32450 26910
rect 32622 26962 32674 26974
rect 32622 26898 32674 26910
rect 34414 26962 34466 26974
rect 34414 26898 34466 26910
rect 37886 26962 37938 26974
rect 37886 26898 37938 26910
rect 45838 26962 45890 26974
rect 45838 26898 45890 26910
rect 46958 26962 47010 26974
rect 46958 26898 47010 26910
rect 49422 26962 49474 26974
rect 55694 26962 55746 26974
rect 55122 26910 55134 26962
rect 55186 26910 55198 26962
rect 49422 26898 49474 26910
rect 55694 26898 55746 26910
rect 2158 26850 2210 26862
rect 2158 26786 2210 26798
rect 2942 26850 2994 26862
rect 2942 26786 2994 26798
rect 3838 26850 3890 26862
rect 3838 26786 3890 26798
rect 7198 26850 7250 26862
rect 7198 26786 7250 26798
rect 8990 26850 9042 26862
rect 8990 26786 9042 26798
rect 10110 26850 10162 26862
rect 10110 26786 10162 26798
rect 12798 26850 12850 26862
rect 12798 26786 12850 26798
rect 15934 26850 15986 26862
rect 15934 26786 15986 26798
rect 16606 26850 16658 26862
rect 16606 26786 16658 26798
rect 19966 26850 20018 26862
rect 19966 26786 20018 26798
rect 24558 26850 24610 26862
rect 24558 26786 24610 26798
rect 31614 26850 31666 26862
rect 31614 26786 31666 26798
rect 33182 26850 33234 26862
rect 33182 26786 33234 26798
rect 35758 26850 35810 26862
rect 35758 26786 35810 26798
rect 36542 26850 36594 26862
rect 38558 26850 38610 26862
rect 37538 26798 37550 26850
rect 37602 26798 37614 26850
rect 36542 26786 36594 26798
rect 38558 26786 38610 26798
rect 45502 26850 45554 26862
rect 45502 26786 45554 26798
rect 47182 26850 47234 26862
rect 47182 26786 47234 26798
rect 47406 26850 47458 26862
rect 50094 26850 50146 26862
rect 49074 26798 49086 26850
rect 49138 26798 49150 26850
rect 47406 26786 47458 26798
rect 50094 26786 50146 26798
rect 50318 26850 50370 26862
rect 57486 26850 57538 26862
rect 57138 26798 57150 26850
rect 57202 26798 57214 26850
rect 50318 26786 50370 26798
rect 57486 26786 57538 26798
rect 1344 26682 58576 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 58576 26682
rect 1344 26596 58576 26630
rect 2494 26514 2546 26526
rect 3838 26514 3890 26526
rect 3490 26462 3502 26514
rect 3554 26462 3566 26514
rect 2494 26450 2546 26462
rect 3838 26450 3890 26462
rect 7870 26514 7922 26526
rect 7870 26450 7922 26462
rect 9662 26514 9714 26526
rect 9662 26450 9714 26462
rect 10894 26514 10946 26526
rect 10894 26450 10946 26462
rect 12798 26514 12850 26526
rect 12798 26450 12850 26462
rect 12910 26514 12962 26526
rect 12910 26450 12962 26462
rect 14702 26514 14754 26526
rect 14702 26450 14754 26462
rect 16830 26514 16882 26526
rect 16830 26450 16882 26462
rect 17838 26514 17890 26526
rect 17838 26450 17890 26462
rect 19294 26514 19346 26526
rect 19294 26450 19346 26462
rect 25902 26514 25954 26526
rect 28254 26514 28306 26526
rect 27122 26462 27134 26514
rect 27186 26462 27198 26514
rect 25902 26450 25954 26462
rect 28254 26450 28306 26462
rect 34750 26514 34802 26526
rect 34750 26450 34802 26462
rect 35870 26514 35922 26526
rect 35870 26450 35922 26462
rect 39118 26514 39170 26526
rect 39118 26450 39170 26462
rect 40238 26514 40290 26526
rect 40238 26450 40290 26462
rect 43710 26514 43762 26526
rect 43710 26450 43762 26462
rect 44046 26514 44098 26526
rect 44046 26450 44098 26462
rect 44830 26514 44882 26526
rect 49870 26514 49922 26526
rect 46610 26462 46622 26514
rect 46674 26462 46686 26514
rect 44830 26450 44882 26462
rect 49870 26450 49922 26462
rect 50766 26514 50818 26526
rect 50766 26450 50818 26462
rect 52110 26514 52162 26526
rect 52110 26450 52162 26462
rect 52782 26514 52834 26526
rect 52782 26450 52834 26462
rect 4398 26402 4450 26414
rect 4398 26338 4450 26350
rect 4734 26402 4786 26414
rect 4734 26338 4786 26350
rect 5406 26402 5458 26414
rect 5406 26338 5458 26350
rect 7086 26402 7138 26414
rect 7086 26338 7138 26350
rect 9886 26402 9938 26414
rect 9886 26338 9938 26350
rect 10558 26402 10610 26414
rect 10558 26338 10610 26350
rect 13022 26402 13074 26414
rect 13022 26338 13074 26350
rect 13134 26402 13186 26414
rect 14590 26402 14642 26414
rect 13346 26350 13358 26402
rect 13410 26350 13422 26402
rect 13134 26338 13186 26350
rect 14590 26338 14642 26350
rect 15486 26402 15538 26414
rect 15486 26338 15538 26350
rect 15598 26402 15650 26414
rect 29486 26402 29538 26414
rect 34414 26402 34466 26414
rect 20402 26350 20414 26402
rect 20466 26350 20478 26402
rect 22194 26350 22206 26402
rect 22258 26350 22270 26402
rect 23538 26350 23550 26402
rect 23602 26350 23614 26402
rect 31714 26350 31726 26402
rect 31778 26350 31790 26402
rect 32162 26350 32174 26402
rect 32226 26350 32238 26402
rect 15598 26338 15650 26350
rect 29486 26338 29538 26350
rect 34414 26338 34466 26350
rect 35422 26402 35474 26414
rect 35422 26338 35474 26350
rect 37998 26402 38050 26414
rect 37998 26338 38050 26350
rect 39342 26402 39394 26414
rect 39342 26338 39394 26350
rect 41582 26402 41634 26414
rect 41582 26338 41634 26350
rect 42702 26402 42754 26414
rect 42702 26338 42754 26350
rect 43822 26402 43874 26414
rect 43822 26338 43874 26350
rect 44270 26402 44322 26414
rect 44270 26338 44322 26350
rect 45054 26402 45106 26414
rect 45054 26338 45106 26350
rect 45166 26402 45218 26414
rect 50094 26402 50146 26414
rect 47730 26350 47742 26402
rect 47794 26350 47806 26402
rect 45166 26338 45218 26350
rect 50094 26338 50146 26350
rect 6750 26290 6802 26302
rect 6750 26226 6802 26238
rect 7198 26290 7250 26302
rect 7198 26226 7250 26238
rect 8430 26290 8482 26302
rect 8430 26226 8482 26238
rect 9998 26290 10050 26302
rect 9998 26226 10050 26238
rect 10894 26290 10946 26302
rect 10894 26226 10946 26238
rect 11118 26290 11170 26302
rect 11118 26226 11170 26238
rect 16270 26290 16322 26302
rect 16270 26226 16322 26238
rect 16718 26290 16770 26302
rect 16718 26226 16770 26238
rect 16942 26290 16994 26302
rect 16942 26226 16994 26238
rect 17614 26290 17666 26302
rect 17614 26226 17666 26238
rect 17950 26290 18002 26302
rect 17950 26226 18002 26238
rect 19182 26290 19234 26302
rect 19182 26226 19234 26238
rect 19406 26290 19458 26302
rect 25678 26290 25730 26302
rect 20290 26238 20302 26290
rect 20354 26238 20366 26290
rect 22642 26238 22654 26290
rect 22706 26238 22718 26290
rect 24210 26238 24222 26290
rect 24274 26238 24286 26290
rect 19406 26226 19458 26238
rect 25678 26226 25730 26238
rect 25902 26290 25954 26302
rect 25902 26226 25954 26238
rect 26238 26290 26290 26302
rect 26238 26226 26290 26238
rect 28590 26290 28642 26302
rect 34638 26290 34690 26302
rect 31266 26238 31278 26290
rect 31330 26238 31342 26290
rect 32050 26238 32062 26290
rect 32114 26238 32126 26290
rect 28590 26226 28642 26238
rect 34638 26226 34690 26238
rect 34862 26290 34914 26302
rect 34862 26226 34914 26238
rect 35646 26290 35698 26302
rect 35646 26226 35698 26238
rect 36094 26290 36146 26302
rect 36094 26226 36146 26238
rect 36430 26290 36482 26302
rect 38222 26290 38274 26302
rect 37426 26238 37438 26290
rect 37490 26238 37502 26290
rect 37762 26238 37774 26290
rect 37826 26238 37838 26290
rect 36430 26226 36482 26238
rect 38222 26226 38274 26238
rect 38670 26290 38722 26302
rect 38670 26226 38722 26238
rect 40014 26290 40066 26302
rect 41806 26290 41858 26302
rect 40450 26238 40462 26290
rect 40514 26238 40526 26290
rect 40674 26238 40686 26290
rect 40738 26238 40750 26290
rect 40014 26226 40066 26238
rect 41806 26226 41858 26238
rect 42814 26290 42866 26302
rect 42814 26226 42866 26238
rect 43150 26290 43202 26302
rect 48078 26290 48130 26302
rect 46834 26238 46846 26290
rect 46898 26238 46910 26290
rect 43150 26226 43202 26238
rect 48078 26226 48130 26238
rect 49758 26290 49810 26302
rect 49758 26226 49810 26238
rect 50318 26290 50370 26302
rect 50318 26226 50370 26238
rect 52894 26290 52946 26302
rect 52894 26226 52946 26238
rect 54014 26290 54066 26302
rect 54898 26238 54910 26290
rect 54962 26238 54974 26290
rect 54014 26226 54066 26238
rect 2158 26178 2210 26190
rect 2158 26114 2210 26126
rect 2942 26178 2994 26190
rect 2942 26114 2994 26126
rect 5854 26178 5906 26190
rect 5854 26114 5906 26126
rect 6302 26178 6354 26190
rect 6302 26114 6354 26126
rect 6862 26178 6914 26190
rect 6862 26114 6914 26126
rect 11790 26178 11842 26190
rect 11790 26114 11842 26126
rect 12238 26178 12290 26190
rect 12238 26114 12290 26126
rect 14478 26178 14530 26190
rect 14478 26114 14530 26126
rect 18958 26178 19010 26190
rect 18958 26114 19010 26126
rect 24894 26178 24946 26190
rect 24894 26114 24946 26126
rect 27694 26178 27746 26190
rect 27694 26114 27746 26126
rect 29038 26178 29090 26190
rect 29038 26114 29090 26126
rect 30046 26178 30098 26190
rect 30046 26114 30098 26126
rect 31726 26178 31778 26190
rect 31726 26114 31778 26126
rect 33518 26178 33570 26190
rect 33518 26114 33570 26126
rect 36878 26178 36930 26190
rect 39230 26178 39282 26190
rect 45614 26178 45666 26190
rect 37874 26126 37886 26178
rect 37938 26126 37950 26178
rect 40786 26126 40798 26178
rect 40850 26126 40862 26178
rect 36878 26114 36930 26126
rect 39230 26114 39282 26126
rect 45614 26114 45666 26126
rect 46062 26178 46114 26190
rect 46062 26114 46114 26126
rect 48526 26178 48578 26190
rect 48526 26114 48578 26126
rect 51214 26178 51266 26190
rect 51214 26114 51266 26126
rect 51662 26178 51714 26190
rect 51662 26114 51714 26126
rect 53454 26178 53506 26190
rect 56590 26178 56642 26190
rect 56018 26126 56030 26178
rect 56082 26126 56094 26178
rect 53454 26114 53506 26126
rect 56590 26114 56642 26126
rect 58046 26178 58098 26190
rect 58046 26114 58098 26126
rect 8654 26066 8706 26078
rect 15486 26066 15538 26078
rect 5170 26014 5182 26066
rect 5234 26063 5246 26066
rect 5842 26063 5854 26066
rect 5234 26017 5854 26063
rect 5234 26014 5246 26017
rect 5842 26014 5854 26017
rect 5906 26014 5918 26066
rect 8978 26014 8990 26066
rect 9042 26014 9054 26066
rect 8654 26002 8706 26014
rect 15486 26002 15538 26014
rect 18510 26066 18562 26078
rect 18510 26002 18562 26014
rect 18734 26066 18786 26078
rect 18734 26002 18786 26014
rect 27470 26066 27522 26078
rect 27470 26002 27522 26014
rect 42142 26066 42194 26078
rect 42142 26002 42194 26014
rect 43038 26066 43090 26078
rect 52782 26066 52834 26078
rect 51090 26014 51102 26066
rect 51154 26063 51166 26066
rect 51762 26063 51774 26066
rect 51154 26017 51774 26063
rect 51154 26014 51166 26017
rect 51762 26014 51774 26017
rect 51826 26014 51838 26066
rect 43038 26002 43090 26014
rect 52782 26002 52834 26014
rect 57486 26066 57538 26078
rect 57486 26002 57538 26014
rect 57822 26066 57874 26078
rect 57822 26002 57874 26014
rect 1344 25898 58576 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 58576 25898
rect 1344 25812 58576 25846
rect 19854 25730 19906 25742
rect 3602 25678 3614 25730
rect 3666 25727 3678 25730
rect 5170 25727 5182 25730
rect 3666 25681 5182 25727
rect 3666 25678 3678 25681
rect 5170 25678 5182 25681
rect 5234 25678 5246 25730
rect 7186 25678 7198 25730
rect 7250 25678 7262 25730
rect 19854 25666 19906 25678
rect 21534 25730 21586 25742
rect 21534 25666 21586 25678
rect 25454 25730 25506 25742
rect 25454 25666 25506 25678
rect 27694 25730 27746 25742
rect 40574 25730 40626 25742
rect 38322 25678 38334 25730
rect 38386 25678 38398 25730
rect 27694 25666 27746 25678
rect 40574 25666 40626 25678
rect 43934 25730 43986 25742
rect 43934 25666 43986 25678
rect 46622 25730 46674 25742
rect 46622 25666 46674 25678
rect 49198 25730 49250 25742
rect 51650 25678 51662 25730
rect 51714 25727 51726 25730
rect 51986 25727 51998 25730
rect 51714 25681 51998 25727
rect 51714 25678 51726 25681
rect 51986 25678 51998 25681
rect 52050 25678 52062 25730
rect 49198 25666 49250 25678
rect 2270 25618 2322 25630
rect 2270 25554 2322 25566
rect 4958 25618 5010 25630
rect 10110 25618 10162 25630
rect 7298 25566 7310 25618
rect 7362 25566 7374 25618
rect 4958 25554 5010 25566
rect 10110 25554 10162 25566
rect 12574 25618 12626 25630
rect 12574 25554 12626 25566
rect 12910 25618 12962 25630
rect 16942 25618 16994 25630
rect 14466 25566 14478 25618
rect 14530 25566 14542 25618
rect 12910 25554 12962 25566
rect 16942 25554 16994 25566
rect 17614 25618 17666 25630
rect 17614 25554 17666 25566
rect 18398 25618 18450 25630
rect 18398 25554 18450 25566
rect 19518 25618 19570 25630
rect 19518 25554 19570 25566
rect 22654 25618 22706 25630
rect 22654 25554 22706 25566
rect 24334 25618 24386 25630
rect 34526 25618 34578 25630
rect 32050 25566 32062 25618
rect 32114 25566 32126 25618
rect 24334 25554 24386 25566
rect 34526 25554 34578 25566
rect 38782 25618 38834 25630
rect 38782 25554 38834 25566
rect 41470 25618 41522 25630
rect 41470 25554 41522 25566
rect 41918 25618 41970 25630
rect 41918 25554 41970 25566
rect 44494 25618 44546 25630
rect 44494 25554 44546 25566
rect 45614 25618 45666 25630
rect 52334 25618 52386 25630
rect 51090 25566 51102 25618
rect 51154 25566 51166 25618
rect 54562 25566 54574 25618
rect 54626 25566 54638 25618
rect 45614 25554 45666 25566
rect 52334 25554 52386 25566
rect 1934 25506 1986 25518
rect 7982 25506 8034 25518
rect 11454 25506 11506 25518
rect 6850 25454 6862 25506
rect 6914 25454 6926 25506
rect 7186 25454 7198 25506
rect 7250 25454 7262 25506
rect 8418 25454 8430 25506
rect 8482 25454 8494 25506
rect 1934 25442 1986 25454
rect 7982 25442 8034 25454
rect 11454 25442 11506 25454
rect 11566 25506 11618 25518
rect 19742 25506 19794 25518
rect 20862 25506 20914 25518
rect 14354 25454 14366 25506
rect 14418 25454 14430 25506
rect 15250 25454 15262 25506
rect 15314 25454 15326 25506
rect 20066 25454 20078 25506
rect 20130 25454 20142 25506
rect 11566 25442 11618 25454
rect 19742 25442 19794 25454
rect 20862 25442 20914 25454
rect 23438 25506 23490 25518
rect 23438 25442 23490 25454
rect 24446 25506 24498 25518
rect 31278 25506 31330 25518
rect 34414 25506 34466 25518
rect 24770 25454 24782 25506
rect 24834 25454 24846 25506
rect 31938 25454 31950 25506
rect 32002 25454 32014 25506
rect 24446 25442 24498 25454
rect 31278 25442 31330 25454
rect 34414 25442 34466 25454
rect 34862 25506 34914 25518
rect 34862 25442 34914 25454
rect 35086 25506 35138 25518
rect 35086 25442 35138 25454
rect 35870 25506 35922 25518
rect 35870 25442 35922 25454
rect 36430 25506 36482 25518
rect 36430 25442 36482 25454
rect 37774 25506 37826 25518
rect 37774 25442 37826 25454
rect 37886 25506 37938 25518
rect 37886 25442 37938 25454
rect 39566 25506 39618 25518
rect 40798 25506 40850 25518
rect 45726 25506 45778 25518
rect 48078 25506 48130 25518
rect 40114 25454 40126 25506
rect 40178 25454 40190 25506
rect 42578 25454 42590 25506
rect 42642 25454 42654 25506
rect 46610 25454 46622 25506
rect 46674 25454 46686 25506
rect 49970 25454 49982 25506
rect 50034 25454 50046 25506
rect 51202 25454 51214 25506
rect 51266 25454 51278 25506
rect 53666 25454 53678 25506
rect 53730 25454 53742 25506
rect 55234 25454 55246 25506
rect 55298 25454 55310 25506
rect 56578 25454 56590 25506
rect 56642 25454 56654 25506
rect 57922 25454 57934 25506
rect 57986 25454 57998 25506
rect 39566 25442 39618 25454
rect 40798 25442 40850 25454
rect 45726 25442 45778 25454
rect 48078 25442 48130 25454
rect 2830 25394 2882 25406
rect 2830 25330 2882 25342
rect 9998 25394 10050 25406
rect 9998 25330 10050 25342
rect 14030 25394 14082 25406
rect 14030 25330 14082 25342
rect 15038 25394 15090 25406
rect 15038 25330 15090 25342
rect 17502 25394 17554 25406
rect 17502 25330 17554 25342
rect 17726 25394 17778 25406
rect 17726 25330 17778 25342
rect 19406 25394 19458 25406
rect 19406 25330 19458 25342
rect 22094 25394 22146 25406
rect 22094 25330 22146 25342
rect 23102 25394 23154 25406
rect 23102 25330 23154 25342
rect 23214 25394 23266 25406
rect 23214 25330 23266 25342
rect 23662 25394 23714 25406
rect 23662 25330 23714 25342
rect 25566 25394 25618 25406
rect 25566 25330 25618 25342
rect 26014 25394 26066 25406
rect 26014 25330 26066 25342
rect 26238 25394 26290 25406
rect 26238 25330 26290 25342
rect 26350 25394 26402 25406
rect 26350 25330 26402 25342
rect 27694 25394 27746 25406
rect 27694 25330 27746 25342
rect 27806 25394 27858 25406
rect 27806 25330 27858 25342
rect 30942 25394 30994 25406
rect 30942 25330 30994 25342
rect 31390 25394 31442 25406
rect 31390 25330 31442 25342
rect 32286 25394 32338 25406
rect 32286 25330 32338 25342
rect 33742 25394 33794 25406
rect 33742 25330 33794 25342
rect 35534 25394 35586 25406
rect 35534 25330 35586 25342
rect 36654 25394 36706 25406
rect 36654 25330 36706 25342
rect 36766 25394 36818 25406
rect 36766 25330 36818 25342
rect 37662 25394 37714 25406
rect 41022 25394 41074 25406
rect 40338 25342 40350 25394
rect 40402 25342 40414 25394
rect 37662 25330 37714 25342
rect 41022 25330 41074 25342
rect 42926 25394 42978 25406
rect 45502 25394 45554 25406
rect 42926 25330 42978 25342
rect 44046 25338 44098 25350
rect 3278 25282 3330 25294
rect 3278 25218 3330 25230
rect 3726 25282 3778 25294
rect 3726 25218 3778 25230
rect 4174 25282 4226 25294
rect 4174 25218 4226 25230
rect 4622 25282 4674 25294
rect 4622 25218 4674 25230
rect 5742 25282 5794 25294
rect 9438 25282 9490 25294
rect 6066 25230 6078 25282
rect 6130 25230 6142 25282
rect 5742 25218 5794 25230
rect 9438 25218 9490 25230
rect 10222 25282 10274 25294
rect 10222 25218 10274 25230
rect 10446 25282 10498 25294
rect 10446 25218 10498 25230
rect 11230 25282 11282 25294
rect 11230 25218 11282 25230
rect 11678 25282 11730 25294
rect 11678 25218 11730 25230
rect 13694 25282 13746 25294
rect 13694 25218 13746 25230
rect 13918 25282 13970 25294
rect 13918 25218 13970 25230
rect 15486 25282 15538 25294
rect 15486 25218 15538 25230
rect 15598 25282 15650 25294
rect 15598 25218 15650 25230
rect 16046 25282 16098 25294
rect 16046 25218 16098 25230
rect 16382 25282 16434 25294
rect 16382 25218 16434 25230
rect 18958 25282 19010 25294
rect 18958 25218 19010 25230
rect 21646 25282 21698 25294
rect 21646 25218 21698 25230
rect 21870 25282 21922 25294
rect 21870 25218 21922 25230
rect 24222 25282 24274 25294
rect 24222 25218 24274 25230
rect 25454 25282 25506 25294
rect 25454 25218 25506 25230
rect 26798 25282 26850 25294
rect 26798 25218 26850 25230
rect 28254 25282 28306 25294
rect 28254 25218 28306 25230
rect 28814 25282 28866 25294
rect 28814 25218 28866 25230
rect 29486 25282 29538 25294
rect 29486 25218 29538 25230
rect 29934 25282 29986 25294
rect 29934 25218 29986 25230
rect 31166 25282 31218 25294
rect 31166 25218 31218 25230
rect 32734 25282 32786 25294
rect 32734 25218 32786 25230
rect 33406 25282 33458 25294
rect 33406 25218 33458 25230
rect 34638 25282 34690 25294
rect 34638 25218 34690 25230
rect 35758 25282 35810 25294
rect 35758 25218 35810 25230
rect 39454 25282 39506 25294
rect 42814 25282 42866 25294
rect 40450 25230 40462 25282
rect 40514 25230 40526 25282
rect 39454 25218 39506 25230
rect 42814 25218 42866 25230
rect 43038 25282 43090 25294
rect 43038 25218 43090 25230
rect 43150 25282 43202 25294
rect 43150 25218 43202 25230
rect 43934 25282 43986 25294
rect 45502 25330 45554 25342
rect 46062 25394 46114 25406
rect 46062 25330 46114 25342
rect 46958 25394 47010 25406
rect 46958 25330 47010 25342
rect 48974 25394 49026 25406
rect 48974 25330 49026 25342
rect 49086 25394 49138 25406
rect 49086 25330 49138 25342
rect 49758 25394 49810 25406
rect 49758 25330 49810 25342
rect 50766 25394 50818 25406
rect 53778 25342 53790 25394
rect 53842 25342 53854 25394
rect 50766 25330 50818 25342
rect 44046 25274 44098 25286
rect 47406 25282 47458 25294
rect 43934 25218 43986 25230
rect 47406 25218 47458 25230
rect 48190 25282 48242 25294
rect 48190 25218 48242 25230
rect 48414 25282 48466 25294
rect 48414 25218 48466 25230
rect 51886 25282 51938 25294
rect 51886 25218 51938 25230
rect 57710 25282 57762 25294
rect 58594 25230 58606 25282
rect 58658 25279 58670 25282
rect 59602 25279 59614 25282
rect 58658 25233 59614 25279
rect 58658 25230 58670 25233
rect 59602 25230 59614 25233
rect 59666 25230 59678 25282
rect 57710 25218 57762 25230
rect 1344 25114 58576 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 58576 25114
rect 1344 25028 58576 25062
rect 1934 24946 1986 24958
rect 1934 24882 1986 24894
rect 12126 24946 12178 24958
rect 12126 24882 12178 24894
rect 16942 24946 16994 24958
rect 16942 24882 16994 24894
rect 19294 24946 19346 24958
rect 27022 24946 27074 24958
rect 21186 24894 21198 24946
rect 21250 24894 21262 24946
rect 19294 24882 19346 24894
rect 27022 24882 27074 24894
rect 28142 24946 28194 24958
rect 28142 24882 28194 24894
rect 32510 24946 32562 24958
rect 32510 24882 32562 24894
rect 32958 24946 33010 24958
rect 32958 24882 33010 24894
rect 33966 24946 34018 24958
rect 33966 24882 34018 24894
rect 37326 24946 37378 24958
rect 37326 24882 37378 24894
rect 38334 24946 38386 24958
rect 38334 24882 38386 24894
rect 38782 24946 38834 24958
rect 38782 24882 38834 24894
rect 39454 24946 39506 24958
rect 39454 24882 39506 24894
rect 41582 24946 41634 24958
rect 52558 24946 52610 24958
rect 45266 24894 45278 24946
rect 45330 24894 45342 24946
rect 41582 24882 41634 24894
rect 52558 24882 52610 24894
rect 53454 24946 53506 24958
rect 53454 24882 53506 24894
rect 54014 24946 54066 24958
rect 54014 24882 54066 24894
rect 54798 24946 54850 24958
rect 54798 24882 54850 24894
rect 56142 24946 56194 24958
rect 56142 24882 56194 24894
rect 56590 24946 56642 24958
rect 56590 24882 56642 24894
rect 2830 24834 2882 24846
rect 18174 24834 18226 24846
rect 26014 24834 26066 24846
rect 9874 24782 9886 24834
rect 9938 24782 9950 24834
rect 21074 24782 21086 24834
rect 21138 24782 21150 24834
rect 24322 24782 24334 24834
rect 24386 24782 24398 24834
rect 2830 24770 2882 24782
rect 18174 24770 18226 24782
rect 26014 24770 26066 24782
rect 27246 24834 27298 24846
rect 27246 24770 27298 24782
rect 29262 24834 29314 24846
rect 29262 24770 29314 24782
rect 34414 24834 34466 24846
rect 34414 24770 34466 24782
rect 35086 24834 35138 24846
rect 35086 24770 35138 24782
rect 35982 24834 36034 24846
rect 35982 24770 36034 24782
rect 42814 24834 42866 24846
rect 50878 24834 50930 24846
rect 45154 24782 45166 24834
rect 45218 24782 45230 24834
rect 45826 24782 45838 24834
rect 45890 24782 45902 24834
rect 47058 24782 47070 24834
rect 47122 24782 47134 24834
rect 42814 24770 42866 24782
rect 50878 24770 50930 24782
rect 52446 24834 52498 24846
rect 57486 24834 57538 24846
rect 55122 24782 55134 24834
rect 55186 24782 55198 24834
rect 55794 24782 55806 24834
rect 55858 24782 55870 24834
rect 52446 24770 52498 24782
rect 57486 24770 57538 24782
rect 57598 24834 57650 24846
rect 57598 24770 57650 24782
rect 12014 24722 12066 24734
rect 4050 24670 4062 24722
rect 4114 24670 4126 24722
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 5842 24670 5854 24722
rect 5906 24670 5918 24722
rect 6962 24670 6974 24722
rect 7026 24670 7038 24722
rect 8418 24670 8430 24722
rect 8482 24670 8494 24722
rect 10434 24670 10446 24722
rect 10498 24670 10510 24722
rect 10770 24670 10782 24722
rect 10834 24670 10846 24722
rect 12014 24658 12066 24670
rect 12350 24722 12402 24734
rect 13470 24722 13522 24734
rect 12786 24670 12798 24722
rect 12850 24670 12862 24722
rect 12350 24658 12402 24670
rect 13470 24658 13522 24670
rect 14030 24722 14082 24734
rect 14030 24658 14082 24670
rect 17838 24722 17890 24734
rect 26910 24722 26962 24734
rect 19058 24670 19070 24722
rect 19122 24670 19134 24722
rect 20178 24670 20190 24722
rect 20242 24670 20254 24722
rect 21970 24670 21982 24722
rect 22034 24670 22046 24722
rect 23986 24670 23998 24722
rect 24050 24670 24062 24722
rect 25778 24670 25790 24722
rect 25842 24670 25854 24722
rect 17838 24658 17890 24670
rect 2382 24610 2434 24622
rect 9102 24610 9154 24622
rect 11566 24610 11618 24622
rect 6626 24558 6638 24610
rect 6690 24558 6702 24610
rect 10098 24558 10110 24610
rect 10162 24558 10174 24610
rect 2382 24546 2434 24558
rect 9102 24546 9154 24558
rect 11566 24546 11618 24558
rect 14814 24610 14866 24622
rect 14814 24546 14866 24558
rect 15150 24610 15202 24622
rect 15150 24546 15202 24558
rect 15598 24610 15650 24622
rect 15598 24546 15650 24558
rect 16046 24610 16098 24622
rect 16046 24546 16098 24558
rect 16494 24610 16546 24622
rect 16494 24546 16546 24558
rect 18734 24610 18786 24622
rect 18734 24546 18786 24558
rect 3054 24498 3106 24510
rect 3054 24434 3106 24446
rect 3390 24498 3442 24510
rect 3390 24434 3442 24446
rect 12462 24498 12514 24510
rect 18386 24446 18398 24498
rect 18450 24495 18462 24498
rect 19073 24495 19119 24670
rect 26910 24658 26962 24670
rect 27358 24722 27410 24734
rect 27358 24658 27410 24670
rect 28030 24722 28082 24734
rect 28030 24658 28082 24670
rect 28254 24722 28306 24734
rect 37214 24722 37266 24734
rect 28578 24670 28590 24722
rect 28642 24670 28654 24722
rect 28254 24658 28306 24670
rect 37214 24658 37266 24670
rect 37550 24722 37602 24734
rect 39902 24722 39954 24734
rect 37762 24670 37774 24722
rect 37826 24670 37838 24722
rect 37550 24658 37602 24670
rect 39902 24658 39954 24670
rect 43150 24722 43202 24734
rect 47518 24722 47570 24734
rect 49534 24722 49586 24734
rect 51102 24722 51154 24734
rect 52782 24722 52834 24734
rect 44146 24670 44158 24722
rect 44210 24670 44222 24722
rect 45042 24670 45054 24722
rect 45106 24670 45118 24722
rect 45602 24670 45614 24722
rect 45666 24670 45678 24722
rect 46722 24670 46734 24722
rect 46786 24670 46798 24722
rect 47954 24670 47966 24722
rect 48018 24670 48030 24722
rect 49858 24670 49870 24722
rect 49922 24670 49934 24722
rect 50418 24670 50430 24722
rect 50482 24670 50494 24722
rect 51202 24670 51214 24722
rect 51266 24670 51278 24722
rect 43150 24658 43202 24670
rect 47518 24658 47570 24670
rect 49534 24658 49586 24670
rect 51102 24658 51154 24670
rect 52782 24658 52834 24670
rect 53006 24722 53058 24734
rect 53006 24658 53058 24670
rect 53566 24722 53618 24734
rect 53566 24658 53618 24670
rect 53790 24722 53842 24734
rect 53790 24658 53842 24670
rect 54126 24722 54178 24734
rect 54126 24658 54178 24670
rect 57710 24722 57762 24734
rect 58034 24670 58046 24722
rect 58098 24670 58110 24722
rect 57710 24658 57762 24670
rect 19630 24610 19682 24622
rect 19630 24546 19682 24558
rect 24894 24610 24946 24622
rect 29934 24610 29986 24622
rect 29138 24558 29150 24610
rect 29202 24558 29214 24610
rect 24894 24546 24946 24558
rect 29934 24546 29986 24558
rect 30382 24610 30434 24622
rect 30382 24546 30434 24558
rect 30830 24610 30882 24622
rect 30830 24546 30882 24558
rect 31614 24610 31666 24622
rect 31614 24546 31666 24558
rect 33518 24610 33570 24622
rect 33518 24546 33570 24558
rect 35534 24610 35586 24622
rect 35534 24546 35586 24558
rect 36430 24610 36482 24622
rect 40798 24610 40850 24622
rect 37650 24558 37662 24610
rect 37714 24558 37726 24610
rect 36430 24546 36482 24558
rect 40798 24546 40850 24558
rect 41918 24610 41970 24622
rect 48638 24610 48690 24622
rect 46946 24558 46958 24610
rect 47010 24558 47022 24610
rect 41918 24546 41970 24558
rect 48638 24546 48690 24558
rect 29486 24498 29538 24510
rect 40126 24498 40178 24510
rect 19618 24495 19630 24498
rect 18450 24449 19630 24495
rect 18450 24446 18462 24449
rect 19618 24446 19630 24449
rect 19682 24446 19694 24498
rect 35970 24446 35982 24498
rect 36034 24495 36046 24498
rect 36418 24495 36430 24498
rect 36034 24449 36430 24495
rect 36034 24446 36046 24449
rect 36418 24446 36430 24449
rect 36482 24446 36494 24498
rect 12462 24434 12514 24446
rect 29486 24434 29538 24446
rect 40126 24434 40178 24446
rect 40238 24498 40290 24510
rect 48402 24446 48414 24498
rect 48466 24495 48478 24498
rect 48626 24495 48638 24498
rect 48466 24449 48638 24495
rect 48466 24446 48478 24449
rect 48626 24446 48638 24449
rect 48690 24446 48702 24498
rect 40238 24434 40290 24446
rect 1344 24330 58576 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 58576 24330
rect 1344 24244 58576 24278
rect 3166 24162 3218 24174
rect 3166 24098 3218 24110
rect 7982 24162 8034 24174
rect 7982 24098 8034 24110
rect 11566 24162 11618 24174
rect 11566 24098 11618 24110
rect 11790 24162 11842 24174
rect 11790 24098 11842 24110
rect 16382 24162 16434 24174
rect 16382 24098 16434 24110
rect 16942 24162 16994 24174
rect 28590 24162 28642 24174
rect 49310 24162 49362 24174
rect 18386 24110 18398 24162
rect 18450 24110 18462 24162
rect 31154 24110 31166 24162
rect 31218 24110 31230 24162
rect 37650 24110 37662 24162
rect 37714 24159 37726 24162
rect 38322 24159 38334 24162
rect 37714 24113 38334 24159
rect 37714 24110 37726 24113
rect 38322 24110 38334 24113
rect 38386 24110 38398 24162
rect 41122 24110 41134 24162
rect 41186 24159 41198 24162
rect 42018 24159 42030 24162
rect 41186 24113 42030 24159
rect 41186 24110 41198 24113
rect 42018 24110 42030 24113
rect 42082 24110 42094 24162
rect 16942 24098 16994 24110
rect 28590 24098 28642 24110
rect 49310 24098 49362 24110
rect 50766 24162 50818 24174
rect 50766 24098 50818 24110
rect 5966 24050 6018 24062
rect 4498 23998 4510 24050
rect 4562 23998 4574 24050
rect 5966 23986 6018 23998
rect 6974 24050 7026 24062
rect 6974 23986 7026 23998
rect 7870 24050 7922 24062
rect 7870 23986 7922 23998
rect 8878 24050 8930 24062
rect 8878 23986 8930 23998
rect 12014 24050 12066 24062
rect 21646 24050 21698 24062
rect 26798 24050 26850 24062
rect 36206 24050 36258 24062
rect 12338 23998 12350 24050
rect 12402 23998 12414 24050
rect 13794 23998 13806 24050
rect 13858 23998 13870 24050
rect 16594 23998 16606 24050
rect 16658 23998 16670 24050
rect 24098 23998 24110 24050
rect 24162 23998 24174 24050
rect 33058 23998 33070 24050
rect 33122 23998 33134 24050
rect 12014 23986 12066 23998
rect 21646 23986 21698 23998
rect 26798 23986 26850 23998
rect 36206 23986 36258 23998
rect 37438 24050 37490 24062
rect 37438 23986 37490 23998
rect 40238 24050 40290 24062
rect 40238 23986 40290 23998
rect 40686 24050 40738 24062
rect 40686 23986 40738 23998
rect 41246 24050 41298 24062
rect 41246 23986 41298 23998
rect 41694 24050 41746 24062
rect 41694 23986 41746 23998
rect 42030 24050 42082 24062
rect 43598 24050 43650 24062
rect 42690 23998 42702 24050
rect 42754 23998 42766 24050
rect 42030 23986 42082 23998
rect 43598 23986 43650 23998
rect 44494 24050 44546 24062
rect 44494 23986 44546 23998
rect 45614 24050 45666 24062
rect 45614 23986 45666 23998
rect 47182 24050 47234 24062
rect 47182 23986 47234 23998
rect 48526 24050 48578 24062
rect 48526 23986 48578 23998
rect 52334 24050 52386 24062
rect 52334 23986 52386 23998
rect 54462 24050 54514 24062
rect 57822 24050 57874 24062
rect 55906 23998 55918 24050
rect 55970 23998 55982 24050
rect 57138 23998 57150 24050
rect 57202 23998 57214 24050
rect 54462 23986 54514 23998
rect 57822 23986 57874 23998
rect 2158 23938 2210 23950
rect 2158 23874 2210 23886
rect 2494 23938 2546 23950
rect 6526 23938 6578 23950
rect 4834 23886 4846 23938
rect 4898 23886 4910 23938
rect 2494 23874 2546 23886
rect 2270 23826 2322 23838
rect 2930 23830 2942 23882
rect 2994 23830 3006 23882
rect 6526 23874 6578 23886
rect 6750 23938 6802 23950
rect 6750 23874 6802 23886
rect 7198 23938 7250 23950
rect 15374 23938 15426 23950
rect 7410 23886 7422 23938
rect 7474 23886 7486 23938
rect 9650 23886 9662 23938
rect 9714 23886 9726 23938
rect 10210 23886 10222 23938
rect 10274 23886 10286 23938
rect 14690 23886 14702 23938
rect 14754 23886 14766 23938
rect 7198 23874 7250 23886
rect 2270 23762 2322 23774
rect 7425 23714 7471 23886
rect 15374 23874 15426 23886
rect 16494 23938 16546 23950
rect 16494 23874 16546 23886
rect 17166 23938 17218 23950
rect 19630 23938 19682 23950
rect 18498 23886 18510 23938
rect 18562 23886 18574 23938
rect 19282 23886 19294 23938
rect 19346 23886 19358 23938
rect 17166 23874 17218 23886
rect 19630 23874 19682 23886
rect 19742 23938 19794 23950
rect 19742 23874 19794 23886
rect 20526 23938 20578 23950
rect 20526 23874 20578 23886
rect 20862 23938 20914 23950
rect 25342 23938 25394 23950
rect 27694 23938 27746 23950
rect 31502 23938 31554 23950
rect 23202 23886 23214 23938
rect 23266 23886 23278 23938
rect 24210 23886 24222 23938
rect 24274 23886 24286 23938
rect 24770 23886 24782 23938
rect 24834 23886 24846 23938
rect 25442 23886 25454 23938
rect 25506 23886 25518 23938
rect 30930 23886 30942 23938
rect 30994 23886 31006 23938
rect 20862 23874 20914 23886
rect 25342 23874 25394 23886
rect 27694 23874 27746 23886
rect 31502 23874 31554 23886
rect 33854 23938 33906 23950
rect 33854 23874 33906 23886
rect 38894 23938 38946 23950
rect 38894 23874 38946 23886
rect 44046 23938 44098 23950
rect 44046 23874 44098 23886
rect 45726 23938 45778 23950
rect 45726 23874 45778 23886
rect 46174 23938 46226 23950
rect 48750 23938 48802 23950
rect 48178 23886 48190 23938
rect 48242 23886 48254 23938
rect 46174 23874 46226 23886
rect 48750 23874 48802 23886
rect 49982 23938 50034 23950
rect 49982 23874 50034 23886
rect 51550 23938 51602 23950
rect 51550 23874 51602 23886
rect 53454 23938 53506 23950
rect 53454 23874 53506 23886
rect 55246 23938 55298 23950
rect 55246 23874 55298 23886
rect 55582 23938 55634 23950
rect 56578 23886 56590 23938
rect 56642 23886 56654 23938
rect 55582 23874 55634 23886
rect 57038 23882 57090 23894
rect 13806 23826 13858 23838
rect 9762 23774 9774 23826
rect 9826 23774 9838 23826
rect 13806 23762 13858 23774
rect 14030 23826 14082 23838
rect 14030 23762 14082 23774
rect 15710 23826 15762 23838
rect 15710 23762 15762 23774
rect 17838 23826 17890 23838
rect 20078 23826 20130 23838
rect 18050 23774 18062 23826
rect 18114 23774 18126 23826
rect 17838 23762 17890 23774
rect 20078 23762 20130 23774
rect 20750 23826 20802 23838
rect 27246 23826 27298 23838
rect 22306 23774 22318 23826
rect 22370 23774 22382 23826
rect 22866 23774 22878 23826
rect 22930 23774 22942 23826
rect 23762 23774 23774 23826
rect 23826 23774 23838 23826
rect 20750 23762 20802 23774
rect 27246 23762 27298 23774
rect 28030 23826 28082 23838
rect 28030 23762 28082 23774
rect 28702 23826 28754 23838
rect 28702 23762 28754 23774
rect 29934 23826 29986 23838
rect 33518 23826 33570 23838
rect 33282 23774 33294 23826
rect 33346 23774 33358 23826
rect 29934 23762 29986 23774
rect 33518 23762 33570 23774
rect 34302 23826 34354 23838
rect 34302 23762 34354 23774
rect 34638 23826 34690 23838
rect 34638 23762 34690 23774
rect 35646 23826 35698 23838
rect 35646 23762 35698 23774
rect 37886 23826 37938 23838
rect 37886 23762 37938 23774
rect 39342 23826 39394 23838
rect 39342 23762 39394 23774
rect 47294 23826 47346 23838
rect 47294 23762 47346 23774
rect 49422 23826 49474 23838
rect 49422 23762 49474 23774
rect 50542 23826 50594 23838
rect 50542 23762 50594 23774
rect 51886 23826 51938 23838
rect 51886 23762 51938 23774
rect 54014 23826 54066 23838
rect 57038 23818 57090 23830
rect 54014 23762 54066 23774
rect 7758 23714 7810 23726
rect 10558 23714 10610 23726
rect 3490 23662 3502 23714
rect 3554 23662 3566 23714
rect 7410 23662 7422 23714
rect 7474 23662 7486 23714
rect 10434 23662 10446 23714
rect 10498 23662 10510 23714
rect 7758 23650 7810 23662
rect 10558 23650 10610 23662
rect 12238 23714 12290 23726
rect 12238 23650 12290 23662
rect 12462 23714 12514 23726
rect 15598 23714 15650 23726
rect 19294 23714 19346 23726
rect 27918 23714 27970 23726
rect 14914 23662 14926 23714
rect 14978 23662 14990 23714
rect 18274 23662 18286 23714
rect 18338 23662 18350 23714
rect 22418 23662 22430 23714
rect 22482 23662 22494 23714
rect 12462 23650 12514 23662
rect 15598 23650 15650 23662
rect 19294 23650 19346 23662
rect 27918 23650 27970 23662
rect 29486 23714 29538 23726
rect 29486 23650 29538 23662
rect 32510 23714 32562 23726
rect 32510 23650 32562 23662
rect 33630 23714 33682 23726
rect 33630 23650 33682 23662
rect 34526 23714 34578 23726
rect 34526 23650 34578 23662
rect 35310 23714 35362 23726
rect 35310 23650 35362 23662
rect 36542 23714 36594 23726
rect 36542 23650 36594 23662
rect 38334 23714 38386 23726
rect 38334 23650 38386 23662
rect 39790 23714 39842 23726
rect 39790 23650 39842 23662
rect 43150 23714 43202 23726
rect 43150 23650 43202 23662
rect 45502 23714 45554 23726
rect 45502 23650 45554 23662
rect 46846 23714 46898 23726
rect 46846 23650 46898 23662
rect 47070 23714 47122 23726
rect 47070 23650 47122 23662
rect 48414 23714 48466 23726
rect 48414 23650 48466 23662
rect 48638 23714 48690 23726
rect 48638 23650 48690 23662
rect 49646 23714 49698 23726
rect 49646 23650 49698 23662
rect 50654 23714 50706 23726
rect 50654 23650 50706 23662
rect 57150 23714 57202 23726
rect 57150 23650 57202 23662
rect 57374 23714 57426 23726
rect 57374 23650 57426 23662
rect 1344 23546 58576 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 58576 23546
rect 1344 23460 58576 23494
rect 8206 23378 8258 23390
rect 11342 23378 11394 23390
rect 5730 23326 5742 23378
rect 5794 23326 5806 23378
rect 8530 23326 8542 23378
rect 8594 23326 8606 23378
rect 8206 23314 8258 23326
rect 11342 23314 11394 23326
rect 17838 23378 17890 23390
rect 23214 23378 23266 23390
rect 20850 23326 20862 23378
rect 20914 23326 20926 23378
rect 17838 23314 17890 23326
rect 23214 23314 23266 23326
rect 25006 23378 25058 23390
rect 25006 23314 25058 23326
rect 28702 23378 28754 23390
rect 28702 23314 28754 23326
rect 29486 23378 29538 23390
rect 29486 23314 29538 23326
rect 32286 23378 32338 23390
rect 32286 23314 32338 23326
rect 32622 23378 32674 23390
rect 32622 23314 32674 23326
rect 33966 23378 34018 23390
rect 33966 23314 34018 23326
rect 36206 23378 36258 23390
rect 36206 23314 36258 23326
rect 36318 23378 36370 23390
rect 36318 23314 36370 23326
rect 39006 23378 39058 23390
rect 39006 23314 39058 23326
rect 40014 23378 40066 23390
rect 40014 23314 40066 23326
rect 40910 23378 40962 23390
rect 40910 23314 40962 23326
rect 42478 23378 42530 23390
rect 42478 23314 42530 23326
rect 44718 23378 44770 23390
rect 44718 23314 44770 23326
rect 45838 23378 45890 23390
rect 45838 23314 45890 23326
rect 46622 23378 46674 23390
rect 46622 23314 46674 23326
rect 47294 23378 47346 23390
rect 47294 23314 47346 23326
rect 48638 23378 48690 23390
rect 48638 23314 48690 23326
rect 51550 23378 51602 23390
rect 51550 23314 51602 23326
rect 54238 23378 54290 23390
rect 54238 23314 54290 23326
rect 55246 23378 55298 23390
rect 55246 23314 55298 23326
rect 57486 23378 57538 23390
rect 57486 23314 57538 23326
rect 14590 23266 14642 23278
rect 18062 23266 18114 23278
rect 6178 23214 6190 23266
rect 6242 23214 6254 23266
rect 10658 23214 10670 23266
rect 10722 23214 10734 23266
rect 13010 23214 13022 23266
rect 13074 23214 13086 23266
rect 15250 23214 15262 23266
rect 15314 23214 15326 23266
rect 15698 23214 15710 23266
rect 15762 23214 15774 23266
rect 14590 23202 14642 23214
rect 18062 23202 18114 23214
rect 18286 23266 18338 23278
rect 18286 23202 18338 23214
rect 19518 23266 19570 23278
rect 21758 23266 21810 23278
rect 20402 23214 20414 23266
rect 20466 23214 20478 23266
rect 20626 23214 20638 23266
rect 20690 23214 20702 23266
rect 19518 23202 19570 23214
rect 21758 23202 21810 23214
rect 25678 23266 25730 23278
rect 31838 23266 31890 23278
rect 27794 23214 27806 23266
rect 27858 23214 27870 23266
rect 25678 23202 25730 23214
rect 31838 23202 31890 23214
rect 32398 23266 32450 23278
rect 32398 23202 32450 23214
rect 33518 23266 33570 23278
rect 33518 23202 33570 23214
rect 40350 23266 40402 23278
rect 40350 23202 40402 23214
rect 41694 23266 41746 23278
rect 41694 23202 41746 23214
rect 41918 23266 41970 23278
rect 41918 23202 41970 23214
rect 44494 23266 44546 23278
rect 44494 23202 44546 23214
rect 45278 23266 45330 23278
rect 45278 23202 45330 23214
rect 48190 23266 48242 23278
rect 49758 23266 49810 23278
rect 54462 23266 54514 23278
rect 49522 23263 49534 23266
rect 48190 23202 48242 23214
rect 49313 23217 49534 23263
rect 14814 23154 14866 23166
rect 3042 23102 3054 23154
rect 3106 23102 3118 23154
rect 4050 23102 4062 23154
rect 4114 23102 4126 23154
rect 4386 23102 4398 23154
rect 4450 23102 4462 23154
rect 5058 23102 5070 23154
rect 5122 23102 5134 23154
rect 7522 23102 7534 23154
rect 7586 23102 7598 23154
rect 10434 23102 10446 23154
rect 10498 23102 10510 23154
rect 11778 23102 11790 23154
rect 11842 23102 11854 23154
rect 13570 23102 13582 23154
rect 13634 23102 13646 23154
rect 14814 23090 14866 23102
rect 17726 23154 17778 23166
rect 17726 23090 17778 23102
rect 21198 23154 21250 23166
rect 23662 23154 23714 23166
rect 29038 23154 29090 23166
rect 21970 23102 21982 23154
rect 22034 23102 22046 23154
rect 22194 23102 22206 23154
rect 22258 23102 22270 23154
rect 26226 23102 26238 23154
rect 26290 23102 26302 23154
rect 27010 23102 27022 23154
rect 27074 23102 27086 23154
rect 27906 23102 27918 23154
rect 27970 23102 27982 23154
rect 21198 23090 21250 23102
rect 23662 23090 23714 23102
rect 29038 23090 29090 23102
rect 29934 23154 29986 23166
rect 31726 23154 31778 23166
rect 31154 23102 31166 23154
rect 31218 23102 31230 23154
rect 29934 23090 29986 23102
rect 31726 23090 31778 23102
rect 32958 23154 33010 23166
rect 32958 23090 33010 23102
rect 34526 23154 34578 23166
rect 34526 23090 34578 23102
rect 34750 23154 34802 23166
rect 34750 23090 34802 23102
rect 35086 23154 35138 23166
rect 36094 23154 36146 23166
rect 37550 23154 37602 23166
rect 35858 23102 35870 23154
rect 35922 23102 35934 23154
rect 36530 23102 36542 23154
rect 36594 23102 36606 23154
rect 35086 23090 35138 23102
rect 36094 23090 36146 23102
rect 37550 23090 37602 23102
rect 37886 23154 37938 23166
rect 37886 23090 37938 23102
rect 38110 23154 38162 23166
rect 38110 23090 38162 23102
rect 39790 23154 39842 23166
rect 39790 23090 39842 23102
rect 40126 23154 40178 23166
rect 40126 23090 40178 23102
rect 43150 23154 43202 23166
rect 43150 23090 43202 23102
rect 43486 23154 43538 23166
rect 43486 23090 43538 23102
rect 43710 23154 43762 23166
rect 43710 23090 43762 23102
rect 44382 23154 44434 23166
rect 44382 23090 44434 23102
rect 45054 23154 45106 23166
rect 45054 23090 45106 23102
rect 45390 23154 45442 23166
rect 49313 23154 49359 23217
rect 49522 23214 49534 23217
rect 49586 23214 49598 23266
rect 50642 23214 50654 23266
rect 50706 23214 50718 23266
rect 52434 23214 52446 23266
rect 52498 23214 52510 23266
rect 49758 23202 49810 23214
rect 54462 23202 54514 23214
rect 57822 23266 57874 23278
rect 57822 23202 57874 23214
rect 50990 23154 51042 23166
rect 54574 23154 54626 23166
rect 46834 23102 46846 23154
rect 46898 23102 46910 23154
rect 49298 23102 49310 23154
rect 49362 23102 49374 23154
rect 52770 23102 52782 23154
rect 52834 23102 52846 23154
rect 53890 23102 53902 23154
rect 53954 23102 53966 23154
rect 45390 23090 45442 23102
rect 50990 23090 51042 23102
rect 54574 23090 54626 23102
rect 55134 23154 55186 23166
rect 55134 23090 55186 23102
rect 55918 23154 55970 23166
rect 55918 23090 55970 23102
rect 56478 23154 56530 23166
rect 56478 23090 56530 23102
rect 1822 23042 1874 23054
rect 1822 22978 1874 22990
rect 2270 23042 2322 23054
rect 2270 22978 2322 22990
rect 8990 23042 9042 23054
rect 8990 22978 9042 22990
rect 16494 23042 16546 23054
rect 16494 22978 16546 22990
rect 16942 23042 16994 23054
rect 16942 22978 16994 22990
rect 19070 23042 19122 23054
rect 19070 22978 19122 22990
rect 22094 23042 22146 23054
rect 22094 22978 22146 22990
rect 22766 23042 22818 23054
rect 22766 22978 22818 22990
rect 24222 23042 24274 23054
rect 34638 23042 34690 23054
rect 27458 22990 27470 23042
rect 27522 22990 27534 23042
rect 24222 22978 24274 22990
rect 34638 22978 34690 22990
rect 36990 23042 37042 23054
rect 36990 22978 37042 22990
rect 37662 23042 37714 23054
rect 37662 22978 37714 22990
rect 38558 23042 38610 23054
rect 43262 23042 43314 23054
rect 41570 22990 41582 23042
rect 41634 22990 41646 23042
rect 38558 22978 38610 22990
rect 43262 22978 43314 22990
rect 47742 23042 47794 23054
rect 47742 22978 47794 22990
rect 51886 23042 51938 23054
rect 53218 22990 53230 23042
rect 53282 22990 53294 23042
rect 51886 22978 51938 22990
rect 25790 22930 25842 22942
rect 25790 22866 25842 22878
rect 26014 22930 26066 22942
rect 26014 22866 26066 22878
rect 46510 22930 46562 22942
rect 49646 22930 49698 22942
rect 47506 22878 47518 22930
rect 47570 22927 47582 22930
rect 48626 22927 48638 22930
rect 47570 22881 48638 22927
rect 47570 22878 47582 22881
rect 48626 22878 48638 22881
rect 48690 22878 48702 22930
rect 46510 22866 46562 22878
rect 49646 22866 49698 22878
rect 49982 22930 50034 22942
rect 49982 22866 50034 22878
rect 55246 22930 55298 22942
rect 55246 22866 55298 22878
rect 1344 22762 58576 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 58576 22762
rect 1344 22676 58576 22710
rect 9214 22594 9266 22606
rect 9214 22530 9266 22542
rect 10782 22594 10834 22606
rect 10782 22530 10834 22542
rect 16046 22594 16098 22606
rect 29934 22594 29986 22606
rect 26786 22542 26798 22594
rect 26850 22542 26862 22594
rect 16046 22530 16098 22542
rect 29934 22530 29986 22542
rect 34526 22594 34578 22606
rect 34526 22530 34578 22542
rect 35758 22594 35810 22606
rect 35758 22530 35810 22542
rect 42814 22594 42866 22606
rect 42814 22530 42866 22542
rect 46958 22594 47010 22606
rect 46958 22530 47010 22542
rect 51326 22594 51378 22606
rect 51326 22530 51378 22542
rect 56590 22594 56642 22606
rect 56590 22530 56642 22542
rect 3726 22482 3778 22494
rect 1922 22430 1934 22482
rect 1986 22430 1998 22482
rect 3726 22418 3778 22430
rect 7534 22482 7586 22494
rect 7534 22418 7586 22430
rect 8542 22482 8594 22494
rect 8542 22418 8594 22430
rect 11790 22482 11842 22494
rect 11790 22418 11842 22430
rect 12574 22482 12626 22494
rect 12574 22418 12626 22430
rect 13022 22482 13074 22494
rect 13022 22418 13074 22430
rect 13806 22482 13858 22494
rect 13806 22418 13858 22430
rect 18734 22482 18786 22494
rect 18734 22418 18786 22430
rect 18958 22482 19010 22494
rect 18958 22418 19010 22430
rect 21646 22482 21698 22494
rect 29598 22482 29650 22494
rect 25554 22430 25566 22482
rect 25618 22430 25630 22482
rect 21646 22418 21698 22430
rect 29598 22418 29650 22430
rect 31390 22482 31442 22494
rect 40126 22482 40178 22494
rect 31938 22430 31950 22482
rect 32002 22430 32014 22482
rect 37986 22430 37998 22482
rect 38050 22430 38062 22482
rect 38994 22430 39006 22482
rect 39058 22430 39070 22482
rect 31390 22418 31442 22430
rect 40126 22418 40178 22430
rect 41022 22482 41074 22494
rect 41022 22418 41074 22430
rect 41470 22482 41522 22494
rect 41470 22418 41522 22430
rect 47294 22482 47346 22494
rect 47294 22418 47346 22430
rect 48862 22482 48914 22494
rect 55794 22430 55806 22482
rect 55858 22430 55870 22482
rect 48862 22418 48914 22430
rect 3614 22370 3666 22382
rect 2818 22318 2830 22370
rect 2882 22318 2894 22370
rect 3614 22306 3666 22318
rect 4286 22370 4338 22382
rect 4286 22306 4338 22318
rect 4958 22370 5010 22382
rect 4958 22306 5010 22318
rect 6302 22370 6354 22382
rect 6302 22306 6354 22318
rect 6638 22370 6690 22382
rect 6638 22306 6690 22318
rect 6974 22370 7026 22382
rect 6974 22306 7026 22318
rect 7422 22370 7474 22382
rect 7422 22306 7474 22318
rect 9326 22370 9378 22382
rect 9326 22306 9378 22318
rect 10110 22370 10162 22382
rect 16606 22370 16658 22382
rect 14242 22318 14254 22370
rect 14306 22318 14318 22370
rect 15362 22318 15374 22370
rect 15426 22318 15438 22370
rect 10110 22306 10162 22318
rect 16606 22306 16658 22318
rect 16942 22370 16994 22382
rect 16942 22306 16994 22318
rect 18174 22370 18226 22382
rect 18174 22306 18226 22318
rect 18622 22370 18674 22382
rect 18622 22306 18674 22318
rect 19182 22370 19234 22382
rect 19182 22306 19234 22318
rect 20078 22370 20130 22382
rect 20078 22306 20130 22318
rect 20638 22370 20690 22382
rect 26350 22370 26402 22382
rect 28590 22370 28642 22382
rect 32286 22370 32338 22382
rect 22866 22318 22878 22370
rect 22930 22318 22942 22370
rect 25666 22318 25678 22370
rect 25730 22318 25742 22370
rect 27458 22318 27470 22370
rect 27522 22318 27534 22370
rect 31826 22318 31838 22370
rect 31890 22318 31902 22370
rect 20638 22306 20690 22318
rect 26350 22306 26402 22318
rect 28590 22306 28642 22318
rect 32286 22306 32338 22318
rect 35870 22370 35922 22382
rect 36542 22370 36594 22382
rect 36418 22318 36430 22370
rect 36482 22318 36494 22370
rect 35870 22306 35922 22318
rect 36542 22306 36594 22318
rect 40014 22370 40066 22382
rect 40014 22306 40066 22318
rect 42478 22370 42530 22382
rect 42478 22306 42530 22318
rect 43038 22370 43090 22382
rect 43038 22306 43090 22318
rect 47070 22370 47122 22382
rect 48974 22370 49026 22382
rect 51438 22370 51490 22382
rect 47506 22318 47518 22370
rect 47570 22318 47582 22370
rect 49746 22318 49758 22370
rect 49810 22318 49822 22370
rect 50194 22318 50206 22370
rect 50258 22318 50270 22370
rect 47070 22306 47122 22318
rect 48974 22306 49026 22318
rect 51438 22306 51490 22318
rect 52110 22370 52162 22382
rect 55022 22370 55074 22382
rect 52322 22318 52334 22370
rect 52386 22318 52398 22370
rect 52110 22306 52162 22318
rect 55022 22306 55074 22318
rect 55246 22370 55298 22382
rect 55246 22306 55298 22318
rect 55470 22370 55522 22382
rect 55470 22306 55522 22318
rect 55694 22370 55746 22382
rect 57586 22318 57598 22370
rect 57650 22318 57662 22370
rect 55694 22306 55746 22318
rect 3838 22258 3890 22270
rect 3838 22194 3890 22206
rect 5854 22258 5906 22270
rect 5854 22194 5906 22206
rect 6414 22258 6466 22270
rect 6414 22194 6466 22206
rect 9214 22258 9266 22270
rect 9214 22194 9266 22206
rect 10670 22258 10722 22270
rect 15934 22258 15986 22270
rect 28254 22258 28306 22270
rect 14578 22206 14590 22258
rect 14642 22206 14654 22258
rect 21970 22206 21982 22258
rect 22034 22206 22046 22258
rect 22754 22206 22766 22258
rect 22818 22206 22830 22258
rect 23538 22206 23550 22258
rect 23602 22206 23614 22258
rect 10670 22194 10722 22206
rect 15934 22194 15986 22206
rect 28254 22194 28306 22206
rect 28478 22258 28530 22270
rect 28478 22194 28530 22206
rect 30158 22258 30210 22270
rect 30158 22194 30210 22206
rect 30606 22258 30658 22270
rect 30606 22194 30658 22206
rect 32510 22258 32562 22270
rect 32510 22194 32562 22206
rect 33518 22258 33570 22270
rect 33518 22194 33570 22206
rect 34302 22258 34354 22270
rect 34302 22194 34354 22206
rect 36654 22258 36706 22270
rect 37998 22258 38050 22270
rect 37874 22206 37886 22258
rect 37938 22206 37950 22258
rect 36654 22194 36706 22206
rect 37998 22194 38050 22206
rect 40462 22258 40514 22270
rect 40462 22194 40514 22206
rect 42254 22258 42306 22270
rect 42254 22194 42306 22206
rect 44046 22258 44098 22270
rect 44046 22194 44098 22206
rect 45838 22258 45890 22270
rect 45838 22194 45890 22206
rect 46174 22258 46226 22270
rect 46174 22194 46226 22206
rect 46398 22258 46450 22270
rect 46398 22194 46450 22206
rect 48414 22258 48466 22270
rect 48414 22194 48466 22206
rect 48638 22258 48690 22270
rect 53454 22258 53506 22270
rect 50754 22206 50766 22258
rect 50818 22206 50830 22258
rect 51986 22206 51998 22258
rect 52050 22206 52062 22258
rect 48638 22194 48690 22206
rect 53454 22194 53506 22206
rect 56926 22258 56978 22270
rect 56926 22194 56978 22206
rect 57822 22258 57874 22270
rect 57822 22194 57874 22206
rect 7646 22146 7698 22158
rect 7646 22082 7698 22094
rect 8094 22146 8146 22158
rect 8094 22082 8146 22094
rect 10446 22146 10498 22158
rect 10446 22082 10498 22094
rect 11230 22146 11282 22158
rect 16046 22146 16098 22158
rect 15138 22094 15150 22146
rect 15202 22094 15214 22146
rect 11230 22082 11282 22094
rect 16046 22082 16098 22094
rect 16830 22146 16882 22158
rect 16830 22082 16882 22094
rect 17838 22146 17890 22158
rect 17838 22082 17890 22094
rect 19294 22146 19346 22158
rect 19294 22082 19346 22094
rect 23886 22146 23938 22158
rect 23886 22082 23938 22094
rect 32062 22146 32114 22158
rect 32062 22082 32114 22094
rect 33182 22146 33234 22158
rect 33182 22082 33234 22094
rect 34414 22146 34466 22158
rect 34414 22082 34466 22094
rect 34974 22146 35026 22158
rect 34974 22082 35026 22094
rect 36206 22146 36258 22158
rect 36206 22082 36258 22094
rect 38110 22146 38162 22158
rect 38110 22082 38162 22094
rect 38334 22146 38386 22158
rect 38334 22082 38386 22094
rect 39454 22146 39506 22158
rect 39454 22082 39506 22094
rect 40238 22146 40290 22158
rect 40238 22082 40290 22094
rect 43150 22146 43202 22158
rect 43150 22082 43202 22094
rect 43710 22146 43762 22158
rect 43710 22082 43762 22094
rect 44494 22146 44546 22158
rect 44494 22082 44546 22094
rect 46062 22146 46114 22158
rect 51774 22146 51826 22158
rect 49746 22094 49758 22146
rect 49810 22094 49822 22146
rect 46062 22082 46114 22094
rect 51774 22082 51826 22094
rect 53790 22146 53842 22158
rect 53790 22082 53842 22094
rect 54238 22146 54290 22158
rect 54238 22082 54290 22094
rect 55918 22146 55970 22158
rect 55918 22082 55970 22094
rect 56702 22146 56754 22158
rect 56702 22082 56754 22094
rect 1344 21978 58576 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 58576 21978
rect 1344 21892 58576 21926
rect 2158 21810 2210 21822
rect 2158 21746 2210 21758
rect 3838 21810 3890 21822
rect 6638 21810 6690 21822
rect 5506 21758 5518 21810
rect 5570 21758 5582 21810
rect 3838 21746 3890 21758
rect 6638 21746 6690 21758
rect 7982 21810 8034 21822
rect 7982 21746 8034 21758
rect 10558 21810 10610 21822
rect 16830 21810 16882 21822
rect 12674 21758 12686 21810
rect 12738 21758 12750 21810
rect 10558 21746 10610 21758
rect 16830 21746 16882 21758
rect 17838 21810 17890 21822
rect 17838 21746 17890 21758
rect 19182 21810 19234 21822
rect 19182 21746 19234 21758
rect 20078 21810 20130 21822
rect 20078 21746 20130 21758
rect 21646 21810 21698 21822
rect 21646 21746 21698 21758
rect 22542 21810 22594 21822
rect 22542 21746 22594 21758
rect 26014 21810 26066 21822
rect 26014 21746 26066 21758
rect 27694 21810 27746 21822
rect 27694 21746 27746 21758
rect 30830 21810 30882 21822
rect 30830 21746 30882 21758
rect 35422 21810 35474 21822
rect 35422 21746 35474 21758
rect 36654 21810 36706 21822
rect 36654 21746 36706 21758
rect 37662 21810 37714 21822
rect 37662 21746 37714 21758
rect 40126 21810 40178 21822
rect 40126 21746 40178 21758
rect 41470 21810 41522 21822
rect 41470 21746 41522 21758
rect 41918 21810 41970 21822
rect 49422 21810 49474 21822
rect 47506 21758 47518 21810
rect 47570 21758 47582 21810
rect 41918 21746 41970 21758
rect 49422 21746 49474 21758
rect 50542 21810 50594 21822
rect 50542 21746 50594 21758
rect 54350 21810 54402 21822
rect 54350 21746 54402 21758
rect 57486 21810 57538 21822
rect 57486 21746 57538 21758
rect 10110 21698 10162 21710
rect 15822 21698 15874 21710
rect 2818 21646 2830 21698
rect 2882 21646 2894 21698
rect 3266 21646 3278 21698
rect 3330 21646 3342 21698
rect 4946 21646 4958 21698
rect 5010 21646 5022 21698
rect 12226 21646 12238 21698
rect 12290 21646 12302 21698
rect 12898 21646 12910 21698
rect 12962 21646 12974 21698
rect 10110 21634 10162 21646
rect 15822 21634 15874 21646
rect 16158 21698 16210 21710
rect 16158 21634 16210 21646
rect 17054 21698 17106 21710
rect 17054 21634 17106 21646
rect 17950 21698 18002 21710
rect 17950 21634 18002 21646
rect 18062 21698 18114 21710
rect 22094 21698 22146 21710
rect 18162 21646 18174 21698
rect 18226 21646 18238 21698
rect 20850 21646 20862 21698
rect 20914 21646 20926 21698
rect 18062 21634 18114 21646
rect 22094 21634 22146 21646
rect 22318 21698 22370 21710
rect 22318 21634 22370 21646
rect 23438 21698 23490 21710
rect 23438 21634 23490 21646
rect 23662 21698 23714 21710
rect 23662 21634 23714 21646
rect 26686 21698 26738 21710
rect 30046 21698 30098 21710
rect 27794 21646 27806 21698
rect 27858 21646 27870 21698
rect 26686 21634 26738 21646
rect 30046 21634 30098 21646
rect 32510 21698 32562 21710
rect 32510 21634 32562 21646
rect 32846 21698 32898 21710
rect 36206 21698 36258 21710
rect 47966 21698 48018 21710
rect 34066 21646 34078 21698
rect 34130 21646 34142 21698
rect 42466 21646 42478 21698
rect 42530 21646 42542 21698
rect 44930 21646 44942 21698
rect 44994 21646 45006 21698
rect 45826 21646 45838 21698
rect 45890 21646 45902 21698
rect 47730 21646 47742 21698
rect 47794 21646 47806 21698
rect 32846 21634 32898 21646
rect 36206 21634 36258 21646
rect 47966 21634 48018 21646
rect 51662 21698 51714 21710
rect 51662 21634 51714 21646
rect 55582 21698 55634 21710
rect 56354 21646 56366 21698
rect 56418 21646 56430 21698
rect 55582 21634 55634 21646
rect 7870 21586 7922 21598
rect 4498 21534 4510 21586
rect 4562 21534 4574 21586
rect 5394 21534 5406 21586
rect 5458 21534 5470 21586
rect 6402 21534 6414 21586
rect 6466 21534 6478 21586
rect 7870 21522 7922 21534
rect 8094 21586 8146 21598
rect 14702 21586 14754 21598
rect 10322 21534 10334 21586
rect 10386 21534 10398 21586
rect 11106 21534 11118 21586
rect 11170 21534 11182 21586
rect 12114 21534 12126 21586
rect 12178 21534 12190 21586
rect 13010 21534 13022 21586
rect 13074 21534 13086 21586
rect 8094 21522 8146 21534
rect 14702 21522 14754 21534
rect 14926 21586 14978 21598
rect 14926 21522 14978 21534
rect 15374 21586 15426 21598
rect 15374 21522 15426 21534
rect 16718 21586 16770 21598
rect 16718 21522 16770 21534
rect 17726 21586 17778 21598
rect 20526 21586 20578 21598
rect 19394 21534 19406 21586
rect 19458 21534 19470 21586
rect 17726 21522 17778 21534
rect 20526 21522 20578 21534
rect 21310 21586 21362 21598
rect 21310 21522 21362 21534
rect 21534 21586 21586 21598
rect 21534 21522 21586 21534
rect 22654 21586 22706 21598
rect 22654 21522 22706 21534
rect 23326 21586 23378 21598
rect 23326 21522 23378 21534
rect 24446 21586 24498 21598
rect 24446 21522 24498 21534
rect 26574 21586 26626 21598
rect 26574 21522 26626 21534
rect 27022 21586 27074 21598
rect 27022 21522 27074 21534
rect 27582 21586 27634 21598
rect 28926 21586 28978 21598
rect 31278 21586 31330 21598
rect 40014 21586 40066 21598
rect 28354 21534 28366 21586
rect 28418 21534 28430 21586
rect 30258 21534 30270 21586
rect 30322 21534 30334 21586
rect 33954 21534 33966 21586
rect 34018 21534 34030 21586
rect 34514 21534 34526 21586
rect 34578 21534 34590 21586
rect 35410 21534 35422 21586
rect 35474 21534 35486 21586
rect 35970 21534 35982 21586
rect 36034 21534 36046 21586
rect 27582 21522 27634 21534
rect 28926 21522 28978 21534
rect 31278 21522 31330 21534
rect 40014 21522 40066 21534
rect 40350 21586 40402 21598
rect 40350 21522 40402 21534
rect 40574 21586 40626 21598
rect 47518 21586 47570 21598
rect 42690 21534 42702 21586
rect 42754 21534 42766 21586
rect 44146 21534 44158 21586
rect 44210 21534 44222 21586
rect 46386 21534 46398 21586
rect 46450 21534 46462 21586
rect 47394 21534 47406 21586
rect 47458 21534 47470 21586
rect 40574 21522 40626 21534
rect 47518 21522 47570 21534
rect 50318 21586 50370 21598
rect 50318 21522 50370 21534
rect 50542 21586 50594 21598
rect 50542 21522 50594 21534
rect 50878 21586 50930 21598
rect 50878 21522 50930 21534
rect 51886 21586 51938 21598
rect 53790 21586 53842 21598
rect 52210 21534 52222 21586
rect 52274 21534 52286 21586
rect 51886 21522 51938 21534
rect 53790 21522 53842 21534
rect 55246 21586 55298 21598
rect 55246 21522 55298 21534
rect 56702 21586 56754 21598
rect 57698 21534 57710 21586
rect 57762 21534 57774 21586
rect 56702 21522 56754 21534
rect 3502 21474 3554 21486
rect 3502 21410 3554 21422
rect 7646 21474 7698 21486
rect 7646 21410 7698 21422
rect 9102 21474 9154 21486
rect 14142 21474 14194 21486
rect 10546 21422 10558 21474
rect 10610 21422 10622 21474
rect 9102 21410 9154 21422
rect 14142 21410 14194 21422
rect 14814 21474 14866 21486
rect 14814 21410 14866 21422
rect 19070 21474 19122 21486
rect 19070 21410 19122 21422
rect 23998 21474 24050 21486
rect 23998 21410 24050 21422
rect 24894 21474 24946 21486
rect 24894 21410 24946 21422
rect 26910 21474 26962 21486
rect 26910 21410 26962 21422
rect 28030 21474 28082 21486
rect 28030 21410 28082 21422
rect 31950 21474 32002 21486
rect 37102 21474 37154 21486
rect 34178 21422 34190 21474
rect 34242 21422 34254 21474
rect 31950 21410 32002 21422
rect 37102 21410 37154 21422
rect 38110 21474 38162 21486
rect 38110 21410 38162 21422
rect 38558 21474 38610 21486
rect 38558 21410 38610 21422
rect 39006 21474 39058 21486
rect 39006 21410 39058 21422
rect 39454 21474 39506 21486
rect 39454 21410 39506 21422
rect 48414 21474 48466 21486
rect 48414 21410 48466 21422
rect 51774 21474 51826 21486
rect 51774 21410 51826 21422
rect 52670 21474 52722 21486
rect 54686 21474 54738 21486
rect 53330 21422 53342 21474
rect 53394 21422 53406 21474
rect 52670 21410 52722 21422
rect 54686 21410 54738 21422
rect 7198 21362 7250 21374
rect 7198 21298 7250 21310
rect 7422 21362 7474 21374
rect 21086 21362 21138 21374
rect 14242 21310 14254 21362
rect 14306 21359 14318 21362
rect 14466 21359 14478 21362
rect 14306 21313 14478 21359
rect 14306 21310 14318 21313
rect 14466 21310 14478 21313
rect 14530 21310 14542 21362
rect 7422 21298 7474 21310
rect 21086 21298 21138 21310
rect 29150 21362 29202 21374
rect 35758 21362 35810 21374
rect 29474 21310 29486 21362
rect 29538 21310 29550 21362
rect 37314 21310 37326 21362
rect 37378 21359 37390 21362
rect 37874 21359 37886 21362
rect 37378 21313 37886 21359
rect 37378 21310 37390 21313
rect 37874 21310 37886 21313
rect 37938 21359 37950 21362
rect 38546 21359 38558 21362
rect 37938 21313 38558 21359
rect 37938 21310 37950 21313
rect 38546 21310 38558 21313
rect 38610 21310 38622 21362
rect 41458 21310 41470 21362
rect 41522 21359 41534 21362
rect 41906 21359 41918 21362
rect 41522 21313 41918 21359
rect 41522 21310 41534 21313
rect 41906 21310 41918 21313
rect 41970 21310 41982 21362
rect 29150 21298 29202 21310
rect 35758 21298 35810 21310
rect 1344 21194 58576 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 58576 21194
rect 1344 21108 58576 21142
rect 20078 21026 20130 21038
rect 18834 20974 18846 21026
rect 18898 21023 18910 21026
rect 19842 21023 19854 21026
rect 18898 20977 19854 21023
rect 18898 20974 18910 20977
rect 19842 20974 19854 20977
rect 19906 20974 19918 21026
rect 20078 20962 20130 20974
rect 23102 21026 23154 21038
rect 23102 20962 23154 20974
rect 23774 21026 23826 21038
rect 37662 21026 37714 21038
rect 31938 20974 31950 21026
rect 32002 21023 32014 21026
rect 32610 21023 32622 21026
rect 32002 20977 32622 21023
rect 32002 20974 32014 20977
rect 32610 20974 32622 20977
rect 32674 20974 32686 21026
rect 34290 20974 34302 21026
rect 34354 21023 34366 21026
rect 34850 21023 34862 21026
rect 34354 20977 34862 21023
rect 34354 20974 34366 20977
rect 34850 20974 34862 20977
rect 34914 20974 34926 21026
rect 23774 20962 23826 20974
rect 37662 20962 37714 20974
rect 40462 21026 40514 21038
rect 40462 20962 40514 20974
rect 41470 21026 41522 21038
rect 42478 21026 42530 21038
rect 41794 20974 41806 21026
rect 41858 20974 41870 21026
rect 41470 20962 41522 20974
rect 42478 20962 42530 20974
rect 46622 21026 46674 21038
rect 46622 20962 46674 20974
rect 47742 21026 47794 21038
rect 57262 21026 57314 21038
rect 47954 20974 47966 21026
rect 48018 21023 48030 21026
rect 48626 21023 48638 21026
rect 48018 20977 48638 21023
rect 48018 20974 48030 20977
rect 48626 20974 48638 20977
rect 48690 20974 48702 21026
rect 48962 20974 48974 21026
rect 49026 21023 49038 21026
rect 49410 21023 49422 21026
rect 49026 20977 49422 21023
rect 49026 20974 49038 20977
rect 49410 20974 49422 20977
rect 49474 20974 49486 21026
rect 50418 21023 50430 21026
rect 50321 20977 50430 21023
rect 47742 20962 47794 20974
rect 1934 20914 1986 20926
rect 1934 20850 1986 20862
rect 2382 20914 2434 20926
rect 2382 20850 2434 20862
rect 2830 20914 2882 20926
rect 2830 20850 2882 20862
rect 4174 20914 4226 20926
rect 4174 20850 4226 20862
rect 6078 20914 6130 20926
rect 12462 20914 12514 20926
rect 8306 20862 8318 20914
rect 8370 20862 8382 20914
rect 6078 20850 6130 20862
rect 12462 20850 12514 20862
rect 13582 20914 13634 20926
rect 15374 20914 15426 20926
rect 14242 20862 14254 20914
rect 14306 20862 14318 20914
rect 13582 20850 13634 20862
rect 15374 20850 15426 20862
rect 15822 20914 15874 20926
rect 15822 20850 15874 20862
rect 16494 20914 16546 20926
rect 16494 20850 16546 20862
rect 18622 20914 18674 20926
rect 18622 20850 18674 20862
rect 20638 20914 20690 20926
rect 25342 20914 25394 20926
rect 24658 20862 24670 20914
rect 24722 20862 24734 20914
rect 20638 20850 20690 20862
rect 25342 20850 25394 20862
rect 26462 20914 26514 20926
rect 29486 20914 29538 20926
rect 27570 20862 27582 20914
rect 27634 20862 27646 20914
rect 26462 20850 26514 20862
rect 29486 20850 29538 20862
rect 32286 20914 32338 20926
rect 32286 20850 32338 20862
rect 32734 20914 32786 20926
rect 32734 20850 32786 20862
rect 33070 20914 33122 20926
rect 33070 20850 33122 20862
rect 34862 20914 34914 20926
rect 34862 20850 34914 20862
rect 36654 20914 36706 20926
rect 36654 20850 36706 20862
rect 38894 20914 38946 20926
rect 38894 20850 38946 20862
rect 45390 20914 45442 20926
rect 45390 20850 45442 20862
rect 48190 20914 48242 20926
rect 48190 20850 48242 20862
rect 6302 20802 6354 20814
rect 12350 20802 12402 20814
rect 6626 20750 6638 20802
rect 6690 20750 6702 20802
rect 7634 20750 7646 20802
rect 7698 20750 7710 20802
rect 8978 20750 8990 20802
rect 9042 20750 9054 20802
rect 10322 20750 10334 20802
rect 10386 20750 10398 20802
rect 6302 20738 6354 20750
rect 12350 20738 12402 20750
rect 14590 20802 14642 20814
rect 18174 20802 18226 20814
rect 16930 20750 16942 20802
rect 16994 20750 17006 20802
rect 14590 20738 14642 20750
rect 18174 20738 18226 20750
rect 20302 20802 20354 20814
rect 20302 20738 20354 20750
rect 22878 20802 22930 20814
rect 22878 20738 22930 20750
rect 23326 20802 23378 20814
rect 23326 20738 23378 20750
rect 24334 20802 24386 20814
rect 24334 20738 24386 20750
rect 25118 20802 25170 20814
rect 25118 20738 25170 20750
rect 25566 20802 25618 20814
rect 30830 20802 30882 20814
rect 27682 20750 27694 20802
rect 27746 20750 27758 20802
rect 28130 20750 28142 20802
rect 28194 20750 28206 20802
rect 30258 20750 30270 20802
rect 30322 20750 30334 20802
rect 25566 20738 25618 20750
rect 30830 20738 30882 20750
rect 33406 20802 33458 20814
rect 33406 20738 33458 20750
rect 33854 20802 33906 20814
rect 33854 20738 33906 20750
rect 35870 20802 35922 20814
rect 35870 20738 35922 20750
rect 37774 20802 37826 20814
rect 37774 20738 37826 20750
rect 38110 20802 38162 20814
rect 38110 20738 38162 20750
rect 38334 20802 38386 20814
rect 41246 20802 41298 20814
rect 40114 20750 40126 20802
rect 40178 20750 40190 20802
rect 38334 20738 38386 20750
rect 41246 20738 41298 20750
rect 42814 20802 42866 20814
rect 42814 20738 42866 20750
rect 43038 20802 43090 20814
rect 43038 20738 43090 20750
rect 4622 20690 4674 20702
rect 12798 20690 12850 20702
rect 7522 20638 7534 20690
rect 7586 20638 7598 20690
rect 4622 20626 4674 20638
rect 12798 20626 12850 20638
rect 14254 20690 14306 20702
rect 14254 20626 14306 20638
rect 14814 20690 14866 20702
rect 14814 20626 14866 20638
rect 17726 20690 17778 20702
rect 17726 20626 17778 20638
rect 19182 20690 19234 20702
rect 19182 20626 19234 20638
rect 19518 20690 19570 20702
rect 19518 20626 19570 20638
rect 25790 20690 25842 20702
rect 33182 20690 33234 20702
rect 27122 20638 27134 20690
rect 27186 20638 27198 20690
rect 28690 20638 28702 20690
rect 28754 20638 28766 20690
rect 25790 20626 25842 20638
rect 33182 20626 33234 20638
rect 37550 20690 37602 20702
rect 37550 20626 37602 20638
rect 39902 20690 39954 20702
rect 39902 20626 39954 20638
rect 43598 20690 43650 20702
rect 43598 20626 43650 20638
rect 46622 20690 46674 20702
rect 46622 20626 46674 20638
rect 46734 20690 46786 20702
rect 46734 20626 46786 20638
rect 47406 20690 47458 20702
rect 50321 20690 50367 20977
rect 50418 20974 50430 20977
rect 50482 20974 50494 21026
rect 57262 20962 57314 20974
rect 50878 20914 50930 20926
rect 50878 20850 50930 20862
rect 53342 20914 53394 20926
rect 53342 20850 53394 20862
rect 56590 20914 56642 20926
rect 56590 20850 56642 20862
rect 57822 20914 57874 20926
rect 57822 20850 57874 20862
rect 54014 20802 54066 20814
rect 57374 20802 57426 20814
rect 55010 20750 55022 20802
rect 55074 20750 55086 20802
rect 54014 20738 54066 20750
rect 57374 20738 57426 20750
rect 51550 20690 51602 20702
rect 50306 20638 50318 20690
rect 50370 20638 50382 20690
rect 47406 20626 47458 20638
rect 51550 20626 51602 20638
rect 51886 20690 51938 20702
rect 51886 20626 51938 20638
rect 54350 20690 54402 20702
rect 56018 20638 56030 20690
rect 56082 20638 56094 20690
rect 54350 20626 54402 20638
rect 3278 20578 3330 20590
rect 3278 20514 3330 20526
rect 3726 20578 3778 20590
rect 3726 20514 3778 20526
rect 5070 20578 5122 20590
rect 5070 20514 5122 20526
rect 11566 20578 11618 20590
rect 11566 20514 11618 20526
rect 12238 20578 12290 20590
rect 12238 20514 12290 20526
rect 12574 20578 12626 20590
rect 12574 20514 12626 20526
rect 14366 20578 14418 20590
rect 14366 20514 14418 20526
rect 16382 20578 16434 20590
rect 16382 20514 16434 20526
rect 16606 20578 16658 20590
rect 16606 20514 16658 20526
rect 20526 20578 20578 20590
rect 20526 20514 20578 20526
rect 20750 20578 20802 20590
rect 20750 20514 20802 20526
rect 21870 20578 21922 20590
rect 21870 20514 21922 20526
rect 22318 20578 22370 20590
rect 22318 20514 22370 20526
rect 24558 20578 24610 20590
rect 31838 20578 31890 20590
rect 30034 20526 30046 20578
rect 30098 20526 30110 20578
rect 24558 20514 24610 20526
rect 31838 20514 31890 20526
rect 33630 20578 33682 20590
rect 33630 20514 33682 20526
rect 34302 20578 34354 20590
rect 34302 20514 34354 20526
rect 35310 20578 35362 20590
rect 35310 20514 35362 20526
rect 36206 20578 36258 20590
rect 36206 20514 36258 20526
rect 39342 20578 39394 20590
rect 39342 20514 39394 20526
rect 40350 20578 40402 20590
rect 40350 20514 40402 20526
rect 43934 20578 43986 20590
rect 43934 20514 43986 20526
rect 44382 20578 44434 20590
rect 44382 20514 44434 20526
rect 45838 20578 45890 20590
rect 45838 20514 45890 20526
rect 47630 20578 47682 20590
rect 47630 20514 47682 20526
rect 48638 20578 48690 20590
rect 48638 20514 48690 20526
rect 49086 20578 49138 20590
rect 49086 20514 49138 20526
rect 49534 20578 49586 20590
rect 49534 20514 49586 20526
rect 49982 20578 50034 20590
rect 49982 20514 50034 20526
rect 50430 20578 50482 20590
rect 50430 20514 50482 20526
rect 51774 20578 51826 20590
rect 51774 20514 51826 20526
rect 52334 20578 52386 20590
rect 52334 20514 52386 20526
rect 54238 20578 54290 20590
rect 54238 20514 54290 20526
rect 1344 20410 58576 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 58576 20410
rect 1344 20324 58576 20358
rect 12350 20242 12402 20254
rect 3042 20190 3054 20242
rect 3106 20190 3118 20242
rect 4274 20190 4286 20242
rect 4338 20190 4350 20242
rect 12350 20178 12402 20190
rect 18510 20242 18562 20254
rect 27358 20242 27410 20254
rect 20178 20190 20190 20242
rect 20242 20190 20254 20242
rect 23650 20190 23662 20242
rect 23714 20190 23726 20242
rect 26226 20190 26238 20242
rect 26290 20190 26302 20242
rect 18510 20178 18562 20190
rect 27358 20178 27410 20190
rect 29934 20242 29986 20254
rect 29934 20178 29986 20190
rect 33630 20242 33682 20254
rect 33630 20178 33682 20190
rect 35758 20242 35810 20254
rect 35758 20178 35810 20190
rect 38446 20242 38498 20254
rect 38446 20178 38498 20190
rect 39566 20242 39618 20254
rect 39566 20178 39618 20190
rect 40126 20242 40178 20254
rect 48526 20242 48578 20254
rect 53566 20242 53618 20254
rect 44258 20190 44270 20242
rect 44322 20190 44334 20242
rect 45826 20190 45838 20242
rect 45890 20190 45902 20242
rect 51538 20190 51550 20242
rect 51602 20190 51614 20242
rect 40126 20178 40178 20190
rect 48526 20178 48578 20190
rect 53566 20178 53618 20190
rect 54574 20242 54626 20254
rect 54574 20178 54626 20190
rect 55582 20242 55634 20254
rect 55582 20178 55634 20190
rect 57822 20242 57874 20254
rect 57822 20178 57874 20190
rect 2158 20130 2210 20142
rect 12238 20130 12290 20142
rect 10658 20078 10670 20130
rect 10722 20078 10734 20130
rect 2158 20066 2210 20078
rect 12238 20066 12290 20078
rect 15038 20130 15090 20142
rect 15038 20066 15090 20078
rect 16158 20130 16210 20142
rect 29038 20130 29090 20142
rect 19842 20078 19854 20130
rect 19906 20078 19918 20130
rect 22418 20078 22430 20130
rect 22482 20078 22494 20130
rect 23762 20078 23774 20130
rect 23826 20078 23838 20130
rect 24322 20078 24334 20130
rect 24386 20078 24398 20130
rect 16158 20066 16210 20078
rect 29038 20066 29090 20078
rect 32510 20130 32562 20142
rect 32510 20066 32562 20078
rect 34078 20130 34130 20142
rect 35198 20130 35250 20142
rect 34850 20078 34862 20130
rect 34914 20078 34926 20130
rect 34078 20066 34130 20078
rect 35198 20066 35250 20078
rect 36766 20130 36818 20142
rect 36766 20066 36818 20078
rect 36990 20130 37042 20142
rect 36990 20066 37042 20078
rect 41582 20130 41634 20142
rect 41582 20066 41634 20078
rect 42814 20130 42866 20142
rect 42814 20066 42866 20078
rect 43038 20130 43090 20142
rect 48414 20130 48466 20142
rect 45266 20078 45278 20130
rect 45330 20078 45342 20130
rect 43038 20066 43090 20078
rect 48414 20066 48466 20078
rect 53006 20130 53058 20142
rect 53006 20066 53058 20078
rect 56702 20130 56754 20142
rect 56702 20066 56754 20078
rect 57486 20130 57538 20142
rect 57486 20066 57538 20078
rect 3390 20018 3442 20030
rect 4958 20018 5010 20030
rect 8430 20018 8482 20030
rect 11790 20018 11842 20030
rect 4498 19966 4510 20018
rect 4562 19966 4574 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 8082 19966 8094 20018
rect 8146 19966 8158 20018
rect 9650 19966 9662 20018
rect 9714 19966 9726 20018
rect 10434 19966 10446 20018
rect 10498 19966 10510 20018
rect 3390 19954 3442 19966
rect 4958 19954 5010 19966
rect 8430 19954 8482 19966
rect 11790 19954 11842 19966
rect 12462 20018 12514 20030
rect 19070 20018 19122 20030
rect 23550 20018 23602 20030
rect 26014 20018 26066 20030
rect 26462 20018 26514 20030
rect 14018 19966 14030 20018
rect 14082 19966 14094 20018
rect 19730 19966 19742 20018
rect 19794 19966 19806 20018
rect 20962 19966 20974 20018
rect 21026 19966 21038 20018
rect 25890 19966 25902 20018
rect 25954 19966 25966 20018
rect 26226 19966 26238 20018
rect 26290 19966 26302 20018
rect 12462 19954 12514 19966
rect 19070 19954 19122 19966
rect 23550 19954 23602 19966
rect 26014 19954 26066 19966
rect 26462 19954 26514 19966
rect 28142 20018 28194 20030
rect 28142 19954 28194 19966
rect 29710 20018 29762 20030
rect 29710 19954 29762 19966
rect 30158 20018 30210 20030
rect 30158 19954 30210 19966
rect 30382 20018 30434 20030
rect 36094 20018 36146 20030
rect 33842 19966 33854 20018
rect 33906 19966 33918 20018
rect 30382 19954 30434 19966
rect 36094 19954 36146 19966
rect 37550 20018 37602 20030
rect 41806 20018 41858 20030
rect 39106 19966 39118 20018
rect 39170 19966 39182 20018
rect 39330 19966 39342 20018
rect 39394 19966 39406 20018
rect 37550 19954 37602 19966
rect 41806 19954 41858 19966
rect 42030 20018 42082 20030
rect 46174 20018 46226 20030
rect 44258 19966 44270 20018
rect 44322 19966 44334 20018
rect 45154 19966 45166 20018
rect 45218 19966 45230 20018
rect 42030 19954 42082 19966
rect 46174 19954 46226 19966
rect 46734 20018 46786 20030
rect 48302 20018 48354 20030
rect 47170 19966 47182 20018
rect 47234 19966 47246 20018
rect 46734 19954 46786 19966
rect 48302 19954 48354 19966
rect 48862 20018 48914 20030
rect 51886 20018 51938 20030
rect 49746 19966 49758 20018
rect 49810 19966 49822 20018
rect 50306 19966 50318 20018
rect 50370 19966 50382 20018
rect 48862 19954 48914 19966
rect 51886 19954 51938 19966
rect 52782 20018 52834 20030
rect 52782 19954 52834 19966
rect 53230 20018 53282 20030
rect 53230 19954 53282 19966
rect 53454 20018 53506 20030
rect 54338 19966 54350 20018
rect 54402 19966 54414 20018
rect 55458 19966 55470 20018
rect 55522 19966 55534 20018
rect 53454 19954 53506 19966
rect 2606 19906 2658 19918
rect 5742 19906 5794 19918
rect 4722 19854 4734 19906
rect 4786 19854 4798 19906
rect 2606 19842 2658 19854
rect 5742 19842 5794 19854
rect 6078 19906 6130 19918
rect 8990 19906 9042 19918
rect 13694 19906 13746 19918
rect 7186 19854 7198 19906
rect 7250 19854 7262 19906
rect 7634 19854 7646 19906
rect 7698 19854 7710 19906
rect 10322 19854 10334 19906
rect 10386 19854 10398 19906
rect 6078 19842 6130 19854
rect 8990 19842 9042 19854
rect 13694 19842 13746 19854
rect 13806 19906 13858 19918
rect 17950 19906 18002 19918
rect 16594 19854 16606 19906
rect 16658 19854 16670 19906
rect 13806 19842 13858 19854
rect 17950 19842 18002 19854
rect 20526 19906 20578 19918
rect 20526 19842 20578 19854
rect 21870 19906 21922 19918
rect 21870 19842 21922 19854
rect 22990 19906 23042 19918
rect 22990 19842 23042 19854
rect 26910 19906 26962 19918
rect 26910 19842 26962 19854
rect 28590 19906 28642 19918
rect 28590 19842 28642 19854
rect 30830 19906 30882 19918
rect 30830 19842 30882 19854
rect 31278 19906 31330 19918
rect 31278 19842 31330 19854
rect 31726 19906 31778 19918
rect 31726 19842 31778 19854
rect 32958 19906 33010 19918
rect 32958 19842 33010 19854
rect 37998 19906 38050 19918
rect 37998 19842 38050 19854
rect 39230 19906 39282 19918
rect 39230 19842 39282 19854
rect 40574 19906 40626 19918
rect 40574 19842 40626 19854
rect 41694 19906 41746 19918
rect 41694 19842 41746 19854
rect 43486 19906 43538 19918
rect 43486 19842 43538 19854
rect 47406 19906 47458 19918
rect 56590 19906 56642 19918
rect 50530 19854 50542 19906
rect 50594 19854 50606 19906
rect 47406 19842 47458 19854
rect 56590 19842 56642 19854
rect 22766 19794 22818 19806
rect 33518 19794 33570 19806
rect 26898 19742 26910 19794
rect 26962 19791 26974 19794
rect 27234 19791 27246 19794
rect 26962 19745 27246 19791
rect 26962 19742 26974 19745
rect 27234 19742 27246 19745
rect 27298 19742 27310 19794
rect 30482 19742 30494 19794
rect 30546 19791 30558 19794
rect 30818 19791 30830 19794
rect 30546 19745 30830 19791
rect 30546 19742 30558 19745
rect 30818 19742 30830 19745
rect 30882 19742 30894 19794
rect 22766 19730 22818 19742
rect 33518 19730 33570 19742
rect 37102 19794 37154 19806
rect 37102 19730 37154 19742
rect 42702 19794 42754 19806
rect 42702 19730 42754 19742
rect 47518 19794 47570 19806
rect 55694 19794 55746 19806
rect 50642 19742 50654 19794
rect 50706 19742 50718 19794
rect 47518 19730 47570 19742
rect 55694 19730 55746 19742
rect 55918 19794 55970 19806
rect 55918 19730 55970 19742
rect 1344 19626 58576 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 58576 19626
rect 1344 19540 58576 19574
rect 5742 19458 5794 19470
rect 5742 19394 5794 19406
rect 12350 19458 12402 19470
rect 12350 19394 12402 19406
rect 12686 19458 12738 19470
rect 12686 19394 12738 19406
rect 14254 19458 14306 19470
rect 14254 19394 14306 19406
rect 15486 19458 15538 19470
rect 15486 19394 15538 19406
rect 21646 19458 21698 19470
rect 21646 19394 21698 19406
rect 21982 19458 22034 19470
rect 27358 19458 27410 19470
rect 23986 19406 23998 19458
rect 24050 19455 24062 19458
rect 24210 19455 24222 19458
rect 24050 19409 24222 19455
rect 24050 19406 24062 19409
rect 24210 19406 24222 19409
rect 24274 19406 24286 19458
rect 21982 19394 22034 19406
rect 27358 19394 27410 19406
rect 35982 19458 36034 19470
rect 35982 19394 36034 19406
rect 36430 19458 36482 19470
rect 36430 19394 36482 19406
rect 45614 19458 45666 19470
rect 45614 19394 45666 19406
rect 46174 19458 46226 19470
rect 46174 19394 46226 19406
rect 53454 19458 53506 19470
rect 53454 19394 53506 19406
rect 54126 19458 54178 19470
rect 54126 19394 54178 19406
rect 7758 19346 7810 19358
rect 13918 19346 13970 19358
rect 10322 19294 10334 19346
rect 10386 19294 10398 19346
rect 7758 19282 7810 19294
rect 13918 19282 13970 19294
rect 15374 19346 15426 19358
rect 15374 19282 15426 19294
rect 16158 19346 16210 19358
rect 16158 19282 16210 19294
rect 16606 19346 16658 19358
rect 16606 19282 16658 19294
rect 17166 19346 17218 19358
rect 17166 19282 17218 19294
rect 18062 19346 18114 19358
rect 22990 19346 23042 19358
rect 19618 19294 19630 19346
rect 19682 19294 19694 19346
rect 20738 19294 20750 19346
rect 20802 19294 20814 19346
rect 18062 19282 18114 19294
rect 22990 19282 23042 19294
rect 23550 19346 23602 19358
rect 23550 19282 23602 19294
rect 24894 19346 24946 19358
rect 24894 19282 24946 19294
rect 25342 19346 25394 19358
rect 25342 19282 25394 19294
rect 25790 19346 25842 19358
rect 25790 19282 25842 19294
rect 31166 19346 31218 19358
rect 31166 19282 31218 19294
rect 33406 19346 33458 19358
rect 33406 19282 33458 19294
rect 33854 19346 33906 19358
rect 33854 19282 33906 19294
rect 34302 19346 34354 19358
rect 34302 19282 34354 19294
rect 41470 19346 41522 19358
rect 41470 19282 41522 19294
rect 42590 19346 42642 19358
rect 42590 19282 42642 19294
rect 42926 19346 42978 19358
rect 48974 19346 49026 19358
rect 44146 19294 44158 19346
rect 44210 19294 44222 19346
rect 45938 19294 45950 19346
rect 46002 19294 46014 19346
rect 47842 19294 47854 19346
rect 47906 19294 47918 19346
rect 42926 19282 42978 19294
rect 48974 19282 49026 19294
rect 50654 19346 50706 19358
rect 54014 19346 54066 19358
rect 51650 19294 51662 19346
rect 51714 19294 51726 19346
rect 50654 19282 50706 19294
rect 54014 19282 54066 19294
rect 57710 19346 57762 19358
rect 57710 19282 57762 19294
rect 2382 19234 2434 19246
rect 2382 19170 2434 19182
rect 3614 19234 3666 19246
rect 8990 19234 9042 19246
rect 12462 19234 12514 19246
rect 13806 19234 13858 19246
rect 6850 19182 6862 19234
rect 6914 19182 6926 19234
rect 10210 19182 10222 19234
rect 10274 19182 10286 19234
rect 10882 19182 10894 19234
rect 10946 19182 10958 19234
rect 12898 19182 12910 19234
rect 12962 19182 12974 19234
rect 3614 19170 3666 19182
rect 8990 19170 9042 19182
rect 12462 19170 12514 19182
rect 13806 19170 13858 19182
rect 14142 19234 14194 19246
rect 14142 19170 14194 19182
rect 17614 19234 17666 19246
rect 17614 19170 17666 19182
rect 18286 19234 18338 19246
rect 23326 19234 23378 19246
rect 19506 19182 19518 19234
rect 19570 19182 19582 19234
rect 20290 19182 20302 19234
rect 20354 19182 20366 19234
rect 18286 19170 18338 19182
rect 23326 19170 23378 19182
rect 26350 19234 26402 19246
rect 26350 19170 26402 19182
rect 26574 19234 26626 19246
rect 26574 19170 26626 19182
rect 27022 19234 27074 19246
rect 27022 19170 27074 19182
rect 28030 19234 28082 19246
rect 28030 19170 28082 19182
rect 30718 19234 30770 19246
rect 30718 19170 30770 19182
rect 32958 19234 33010 19246
rect 32958 19170 33010 19182
rect 34750 19234 34802 19246
rect 34750 19170 34802 19182
rect 35310 19234 35362 19246
rect 35310 19170 35362 19182
rect 36094 19234 36146 19246
rect 36094 19170 36146 19182
rect 36654 19234 36706 19246
rect 36654 19170 36706 19182
rect 37662 19234 37714 19246
rect 37662 19170 37714 19182
rect 38334 19234 38386 19246
rect 40014 19234 40066 19246
rect 38882 19182 38894 19234
rect 38946 19182 38958 19234
rect 38334 19170 38386 19182
rect 40014 19170 40066 19182
rect 42030 19234 42082 19246
rect 46398 19234 46450 19246
rect 43810 19182 43822 19234
rect 43874 19182 43886 19234
rect 44034 19182 44046 19234
rect 44098 19182 44110 19234
rect 42030 19170 42082 19182
rect 46398 19170 46450 19182
rect 48750 19234 48802 19246
rect 48750 19170 48802 19182
rect 49086 19234 49138 19246
rect 49086 19170 49138 19182
rect 49870 19234 49922 19246
rect 53566 19234 53618 19246
rect 51426 19182 51438 19234
rect 51490 19182 51502 19234
rect 52210 19182 52222 19234
rect 52274 19182 52286 19234
rect 49870 19170 49922 19182
rect 53566 19170 53618 19182
rect 53790 19234 53842 19246
rect 53790 19170 53842 19182
rect 3278 19122 3330 19134
rect 3278 19058 3330 19070
rect 4062 19122 4114 19134
rect 15262 19122 15314 19134
rect 4946 19070 4958 19122
rect 5010 19070 5022 19122
rect 6626 19070 6638 19122
rect 6690 19070 6702 19122
rect 8642 19070 8654 19122
rect 8706 19070 8718 19122
rect 9650 19070 9662 19122
rect 9714 19070 9726 19122
rect 4062 19058 4114 19070
rect 15262 19058 15314 19070
rect 17838 19122 17890 19134
rect 27470 19122 27522 19134
rect 19282 19070 19294 19122
rect 19346 19070 19358 19122
rect 17838 19058 17890 19070
rect 27470 19058 27522 19070
rect 27694 19122 27746 19134
rect 27694 19058 27746 19070
rect 28478 19122 28530 19134
rect 28478 19058 28530 19070
rect 28814 19122 28866 19134
rect 28814 19058 28866 19070
rect 29598 19122 29650 19134
rect 29598 19058 29650 19070
rect 29934 19122 29986 19134
rect 29934 19058 29986 19070
rect 30606 19122 30658 19134
rect 30606 19058 30658 19070
rect 34862 19122 34914 19134
rect 34862 19058 34914 19070
rect 35086 19122 35138 19134
rect 35870 19122 35922 19134
rect 35522 19070 35534 19122
rect 35586 19119 35598 19122
rect 35746 19119 35758 19122
rect 35586 19073 35758 19119
rect 35586 19070 35598 19073
rect 35746 19070 35758 19073
rect 35810 19070 35822 19122
rect 35086 19058 35138 19070
rect 35870 19058 35922 19070
rect 37886 19122 37938 19134
rect 40462 19122 40514 19134
rect 45838 19122 45890 19134
rect 55806 19122 55858 19134
rect 39106 19070 39118 19122
rect 39170 19070 39182 19122
rect 39666 19070 39678 19122
rect 39730 19070 39742 19122
rect 40786 19070 40798 19122
rect 40850 19070 40862 19122
rect 47618 19070 47630 19122
rect 47682 19070 47694 19122
rect 52098 19070 52110 19122
rect 52162 19070 52174 19122
rect 37886 19058 37938 19070
rect 40462 19058 40514 19070
rect 45838 19058 45890 19070
rect 55806 19058 55858 19070
rect 56926 19122 56978 19134
rect 56926 19058 56978 19070
rect 57262 19122 57314 19134
rect 57262 19058 57314 19070
rect 1934 19010 1986 19022
rect 1934 18946 1986 18958
rect 2830 19010 2882 19022
rect 2830 18946 2882 18958
rect 4622 19010 4674 19022
rect 4622 18946 4674 18958
rect 5854 19010 5906 19022
rect 5854 18946 5906 18958
rect 5966 19010 6018 19022
rect 5966 18946 6018 18958
rect 8094 19010 8146 19022
rect 8094 18946 8146 18958
rect 11342 19010 11394 19022
rect 11342 18946 11394 18958
rect 11790 19010 11842 19022
rect 11790 18946 11842 18958
rect 18622 19010 18674 19022
rect 18622 18946 18674 18958
rect 21758 19010 21810 19022
rect 21758 18946 21810 18958
rect 22878 19010 22930 19022
rect 22878 18946 22930 18958
rect 23102 19010 23154 19022
rect 23102 18946 23154 18958
rect 24222 19010 24274 19022
rect 24222 18946 24274 18958
rect 26462 19010 26514 19022
rect 26462 18946 26514 18958
rect 30382 19010 30434 19022
rect 30382 18946 30434 18958
rect 31838 19010 31890 19022
rect 31838 18946 31890 18958
rect 32510 19010 32562 19022
rect 32510 18946 32562 18958
rect 37774 19010 37826 19022
rect 46958 19010 47010 19022
rect 54686 19010 54738 19022
rect 44706 18958 44718 19010
rect 44770 18958 44782 19010
rect 50194 18958 50206 19010
rect 50258 18958 50270 19010
rect 37774 18946 37826 18958
rect 46958 18946 47010 18958
rect 54686 18946 54738 18958
rect 55470 19010 55522 19022
rect 55470 18946 55522 18958
rect 56254 19010 56306 19022
rect 56254 18946 56306 18958
rect 1344 18842 58576 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 58576 18842
rect 1344 18756 58576 18790
rect 3614 18674 3666 18686
rect 3614 18610 3666 18622
rect 3726 18674 3778 18686
rect 3726 18610 3778 18622
rect 4958 18674 5010 18686
rect 4958 18610 5010 18622
rect 5966 18674 6018 18686
rect 5966 18610 6018 18622
rect 6078 18674 6130 18686
rect 13918 18674 13970 18686
rect 8530 18622 8542 18674
rect 8594 18622 8606 18674
rect 6078 18610 6130 18622
rect 13918 18610 13970 18622
rect 14702 18674 14754 18686
rect 20750 18674 20802 18686
rect 14702 18610 14754 18622
rect 14814 18618 14866 18630
rect 6190 18562 6242 18574
rect 7870 18562 7922 18574
rect 6962 18510 6974 18562
rect 7026 18510 7038 18562
rect 6190 18498 6242 18510
rect 7870 18498 7922 18510
rect 8094 18562 8146 18574
rect 8094 18498 8146 18510
rect 13806 18562 13858 18574
rect 20750 18610 20802 18622
rect 20862 18674 20914 18686
rect 20862 18610 20914 18622
rect 21982 18674 22034 18686
rect 21982 18610 22034 18622
rect 23998 18674 24050 18686
rect 23998 18610 24050 18622
rect 24110 18674 24162 18686
rect 24110 18610 24162 18622
rect 24894 18674 24946 18686
rect 27022 18674 27074 18686
rect 30158 18674 30210 18686
rect 26226 18622 26238 18674
rect 26290 18622 26302 18674
rect 27570 18622 27582 18674
rect 27634 18622 27646 18674
rect 29698 18622 29710 18674
rect 29762 18622 29774 18674
rect 24894 18610 24946 18622
rect 27022 18610 27074 18622
rect 30158 18610 30210 18622
rect 31278 18674 31330 18686
rect 31278 18610 31330 18622
rect 31502 18674 31554 18686
rect 31502 18610 31554 18622
rect 34302 18674 34354 18686
rect 34302 18610 34354 18622
rect 35870 18674 35922 18686
rect 35870 18610 35922 18622
rect 37438 18674 37490 18686
rect 37438 18610 37490 18622
rect 38222 18674 38274 18686
rect 38222 18610 38274 18622
rect 38782 18674 38834 18686
rect 38782 18610 38834 18622
rect 39566 18674 39618 18686
rect 39566 18610 39618 18622
rect 40686 18674 40738 18686
rect 40686 18610 40738 18622
rect 42030 18674 42082 18686
rect 42030 18610 42082 18622
rect 45614 18674 45666 18686
rect 45614 18610 45666 18622
rect 46622 18674 46674 18686
rect 46622 18610 46674 18622
rect 48526 18674 48578 18686
rect 49870 18674 49922 18686
rect 49522 18622 49534 18674
rect 49586 18622 49598 18674
rect 48526 18610 48578 18622
rect 49870 18610 49922 18622
rect 50318 18674 50370 18686
rect 54798 18674 54850 18686
rect 57822 18674 57874 18686
rect 51538 18622 51550 18674
rect 51602 18622 51614 18674
rect 52770 18622 52782 18674
rect 52834 18622 52846 18674
rect 56466 18622 56478 18674
rect 56530 18622 56542 18674
rect 50318 18610 50370 18622
rect 54798 18610 54850 18622
rect 57822 18610 57874 18622
rect 14814 18554 14866 18566
rect 15374 18562 15426 18574
rect 13806 18498 13858 18510
rect 15374 18498 15426 18510
rect 15598 18562 15650 18574
rect 15598 18498 15650 18510
rect 15710 18562 15762 18574
rect 21870 18562 21922 18574
rect 15922 18510 15934 18562
rect 15986 18510 15998 18562
rect 15710 18498 15762 18510
rect 21870 18498 21922 18510
rect 24222 18562 24274 18574
rect 24222 18498 24274 18510
rect 32174 18562 32226 18574
rect 32174 18498 32226 18510
rect 32510 18562 32562 18574
rect 32510 18498 32562 18510
rect 35982 18562 36034 18574
rect 37102 18562 37154 18574
rect 36866 18510 36878 18562
rect 36930 18510 36942 18562
rect 35982 18498 36034 18510
rect 37102 18498 37154 18510
rect 37214 18562 37266 18574
rect 37214 18498 37266 18510
rect 37326 18562 37378 18574
rect 37326 18498 37378 18510
rect 39118 18562 39170 18574
rect 39118 18498 39170 18510
rect 40574 18562 40626 18574
rect 40574 18498 40626 18510
rect 40798 18562 40850 18574
rect 42254 18562 42306 18574
rect 41010 18510 41022 18562
rect 41074 18510 41086 18562
rect 40798 18498 40850 18510
rect 3054 18450 3106 18462
rect 3054 18386 3106 18398
rect 3502 18450 3554 18462
rect 3502 18386 3554 18398
rect 4622 18450 4674 18462
rect 4622 18386 4674 18398
rect 5518 18450 5570 18462
rect 5518 18386 5570 18398
rect 7310 18450 7362 18462
rect 7310 18386 7362 18398
rect 8318 18450 8370 18462
rect 8318 18386 8370 18398
rect 8542 18450 8594 18462
rect 8542 18386 8594 18398
rect 8990 18450 9042 18462
rect 8990 18386 9042 18398
rect 9774 18450 9826 18462
rect 9774 18386 9826 18398
rect 10782 18450 10834 18462
rect 10782 18386 10834 18398
rect 12350 18450 12402 18462
rect 12350 18386 12402 18398
rect 14142 18450 14194 18462
rect 19182 18450 19234 18462
rect 20638 18450 20690 18462
rect 18050 18398 18062 18450
rect 18114 18398 18126 18450
rect 18274 18398 18286 18450
rect 18338 18398 18350 18450
rect 19394 18398 19406 18450
rect 19458 18398 19470 18450
rect 14142 18386 14194 18398
rect 19182 18386 19234 18398
rect 20638 18386 20690 18398
rect 21310 18450 21362 18462
rect 21310 18386 21362 18398
rect 23550 18450 23602 18462
rect 26574 18450 26626 18462
rect 23874 18398 23886 18450
rect 23938 18398 23950 18450
rect 23550 18386 23602 18398
rect 26574 18386 26626 18398
rect 27918 18450 27970 18462
rect 27918 18386 27970 18398
rect 28366 18450 28418 18462
rect 28366 18386 28418 18398
rect 28926 18450 28978 18462
rect 28926 18386 28978 18398
rect 29374 18450 29426 18462
rect 32622 18450 32674 18462
rect 31154 18398 31166 18450
rect 31218 18398 31230 18450
rect 29374 18386 29426 18398
rect 32622 18386 32674 18398
rect 35646 18450 35698 18462
rect 35646 18386 35698 18398
rect 40126 18450 40178 18462
rect 40126 18386 40178 18398
rect 1822 18338 1874 18350
rect 1822 18274 1874 18286
rect 2270 18338 2322 18350
rect 2270 18274 2322 18286
rect 2718 18338 2770 18350
rect 11454 18338 11506 18350
rect 4834 18286 4846 18338
rect 4898 18286 4910 18338
rect 10322 18286 10334 18338
rect 10386 18286 10398 18338
rect 2718 18274 2770 18286
rect 11454 18274 11506 18286
rect 11902 18338 11954 18350
rect 11902 18274 11954 18286
rect 12798 18338 12850 18350
rect 12798 18274 12850 18286
rect 13358 18338 13410 18350
rect 17054 18338 17106 18350
rect 22878 18338 22930 18350
rect 16146 18286 16158 18338
rect 16210 18286 16222 18338
rect 18162 18286 18174 18338
rect 18226 18286 18238 18338
rect 13358 18274 13410 18286
rect 17054 18274 17106 18286
rect 22878 18274 22930 18286
rect 25678 18338 25730 18350
rect 25678 18274 25730 18286
rect 31390 18338 31442 18350
rect 31390 18274 31442 18286
rect 32286 18338 32338 18350
rect 32286 18274 32338 18286
rect 34862 18338 34914 18350
rect 41025 18338 41071 18510
rect 42254 18498 42306 18510
rect 42478 18562 42530 18574
rect 42478 18498 42530 18510
rect 44158 18562 44210 18574
rect 44158 18498 44210 18510
rect 44270 18562 44322 18574
rect 44270 18498 44322 18510
rect 46062 18562 46114 18574
rect 46062 18498 46114 18510
rect 46958 18562 47010 18574
rect 46958 18498 47010 18510
rect 48638 18562 48690 18574
rect 48638 18498 48690 18510
rect 51886 18562 51938 18574
rect 51886 18498 51938 18510
rect 52446 18562 52498 18574
rect 52446 18498 52498 18510
rect 54910 18562 54962 18574
rect 55906 18510 55918 18562
rect 55970 18510 55982 18562
rect 57474 18510 57486 18562
rect 57538 18510 57550 18562
rect 54910 18498 54962 18510
rect 41806 18450 41858 18462
rect 41806 18386 41858 18398
rect 44718 18450 44770 18462
rect 44718 18386 44770 18398
rect 45390 18450 45442 18462
rect 45390 18386 45442 18398
rect 45726 18450 45778 18462
rect 45726 18386 45778 18398
rect 47630 18450 47682 18462
rect 47630 18386 47682 18398
rect 54238 18450 54290 18462
rect 54238 18386 54290 18398
rect 54686 18450 54738 18462
rect 55794 18398 55806 18450
rect 55858 18398 55870 18450
rect 56354 18398 56366 18450
rect 56418 18398 56430 18450
rect 54686 18386 54738 18398
rect 43038 18338 43090 18350
rect 41010 18286 41022 18338
rect 41074 18286 41086 18338
rect 34862 18274 34914 18286
rect 43038 18274 43090 18286
rect 43374 18338 43426 18350
rect 43374 18274 43426 18286
rect 50766 18338 50818 18350
rect 50766 18274 50818 18286
rect 53342 18338 53394 18350
rect 53342 18274 53394 18286
rect 53790 18338 53842 18350
rect 53790 18274 53842 18286
rect 14702 18226 14754 18238
rect 22094 18226 22146 18238
rect 1698 18174 1710 18226
rect 1762 18223 1774 18226
rect 2706 18223 2718 18226
rect 1762 18177 2718 18223
rect 1762 18174 1774 18177
rect 2706 18174 2718 18177
rect 2770 18174 2782 18226
rect 12898 18174 12910 18226
rect 12962 18223 12974 18226
rect 13234 18223 13246 18226
rect 12962 18177 13246 18223
rect 12962 18174 12974 18177
rect 13234 18174 13246 18177
rect 13298 18174 13310 18226
rect 18722 18174 18734 18226
rect 18786 18174 18798 18226
rect 14702 18162 14754 18174
rect 22094 18162 22146 18174
rect 23326 18226 23378 18238
rect 23326 18162 23378 18174
rect 30830 18226 30882 18238
rect 30830 18162 30882 18174
rect 33742 18226 33794 18238
rect 33742 18162 33794 18174
rect 33966 18226 34018 18238
rect 33966 18162 34018 18174
rect 34190 18226 34242 18238
rect 34190 18162 34242 18174
rect 34302 18226 34354 18238
rect 34302 18162 34354 18174
rect 41918 18226 41970 18238
rect 41918 18162 41970 18174
rect 44158 18226 44210 18238
rect 44158 18162 44210 18174
rect 48414 18226 48466 18238
rect 48414 18162 48466 18174
rect 1344 18058 58576 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 58576 18058
rect 1344 17972 58576 18006
rect 7534 17890 7586 17902
rect 3938 17838 3950 17890
rect 4002 17887 4014 17890
rect 4834 17887 4846 17890
rect 4002 17841 4846 17887
rect 4002 17838 4014 17841
rect 4834 17838 4846 17841
rect 4898 17838 4910 17890
rect 7534 17826 7586 17838
rect 9214 17890 9266 17902
rect 11678 17890 11730 17902
rect 10210 17838 10222 17890
rect 10274 17838 10286 17890
rect 9214 17826 9266 17838
rect 11678 17826 11730 17838
rect 17950 17890 18002 17902
rect 27246 17890 27298 17902
rect 18274 17838 18286 17890
rect 18338 17838 18350 17890
rect 25442 17838 25454 17890
rect 25506 17887 25518 17890
rect 25666 17887 25678 17890
rect 25506 17841 25678 17887
rect 25506 17838 25518 17841
rect 25666 17838 25678 17841
rect 25730 17838 25742 17890
rect 17950 17826 18002 17838
rect 27246 17826 27298 17838
rect 31166 17890 31218 17902
rect 35534 17890 35586 17902
rect 40350 17890 40402 17902
rect 55582 17890 55634 17902
rect 34850 17838 34862 17890
rect 34914 17887 34926 17890
rect 35074 17887 35086 17890
rect 34914 17841 35086 17887
rect 34914 17838 34926 17841
rect 35074 17838 35086 17841
rect 35138 17838 35150 17890
rect 36082 17838 36094 17890
rect 36146 17887 36158 17890
rect 36642 17887 36654 17890
rect 36146 17841 36654 17887
rect 36146 17838 36158 17841
rect 36642 17838 36654 17841
rect 36706 17838 36718 17890
rect 42466 17838 42478 17890
rect 42530 17838 42542 17890
rect 46050 17838 46062 17890
rect 46114 17887 46126 17890
rect 46722 17887 46734 17890
rect 46114 17841 46734 17887
rect 46114 17838 46126 17841
rect 46722 17838 46734 17841
rect 46786 17838 46798 17890
rect 50306 17838 50318 17890
rect 50370 17887 50382 17890
rect 51314 17887 51326 17890
rect 50370 17841 51326 17887
rect 50370 17838 50382 17841
rect 51314 17838 51326 17841
rect 51378 17838 51390 17890
rect 31166 17826 31218 17838
rect 35534 17826 35586 17838
rect 40350 17826 40402 17838
rect 55582 17826 55634 17838
rect 56814 17890 56866 17902
rect 56814 17826 56866 17838
rect 6526 17778 6578 17790
rect 3042 17726 3054 17778
rect 3106 17726 3118 17778
rect 6526 17714 6578 17726
rect 8206 17778 8258 17790
rect 8206 17714 8258 17726
rect 9662 17778 9714 17790
rect 9662 17714 9714 17726
rect 12462 17778 12514 17790
rect 12462 17714 12514 17726
rect 12910 17778 12962 17790
rect 17278 17778 17330 17790
rect 15474 17726 15486 17778
rect 15538 17726 15550 17778
rect 16258 17726 16270 17778
rect 16322 17726 16334 17778
rect 12910 17714 12962 17726
rect 17278 17714 17330 17726
rect 20414 17778 20466 17790
rect 20414 17714 20466 17726
rect 24446 17778 24498 17790
rect 24446 17714 24498 17726
rect 32510 17778 32562 17790
rect 32510 17714 32562 17726
rect 33966 17778 34018 17790
rect 33966 17714 34018 17726
rect 34638 17778 34690 17790
rect 34638 17714 34690 17726
rect 36430 17778 36482 17790
rect 36430 17714 36482 17726
rect 36878 17778 36930 17790
rect 36878 17714 36930 17726
rect 37438 17778 37490 17790
rect 37438 17714 37490 17726
rect 39006 17778 39058 17790
rect 39006 17714 39058 17726
rect 39678 17778 39730 17790
rect 39678 17714 39730 17726
rect 40798 17778 40850 17790
rect 42142 17778 42194 17790
rect 41010 17726 41022 17778
rect 41074 17726 41086 17778
rect 40798 17714 40850 17726
rect 42142 17714 42194 17726
rect 42926 17778 42978 17790
rect 42926 17714 42978 17726
rect 46734 17778 46786 17790
rect 46734 17714 46786 17726
rect 47182 17778 47234 17790
rect 47182 17714 47234 17726
rect 48750 17778 48802 17790
rect 48750 17714 48802 17726
rect 49198 17778 49250 17790
rect 49198 17714 49250 17726
rect 49646 17778 49698 17790
rect 49646 17714 49698 17726
rect 50878 17778 50930 17790
rect 50878 17714 50930 17726
rect 52334 17778 52386 17790
rect 52334 17714 52386 17726
rect 52670 17778 52722 17790
rect 52670 17714 52722 17726
rect 9886 17666 9938 17678
rect 11006 17666 11058 17678
rect 11790 17666 11842 17678
rect 7634 17614 7646 17666
rect 7698 17614 7710 17666
rect 8754 17614 8766 17666
rect 8818 17614 8830 17666
rect 10770 17614 10782 17666
rect 10834 17614 10846 17666
rect 11106 17614 11118 17666
rect 11170 17614 11182 17666
rect 9886 17602 9938 17614
rect 11006 17602 11058 17614
rect 11790 17602 11842 17614
rect 13806 17666 13858 17678
rect 13806 17602 13858 17614
rect 14030 17666 14082 17678
rect 17726 17666 17778 17678
rect 14354 17614 14366 17666
rect 14418 17614 14430 17666
rect 15138 17614 15150 17666
rect 15202 17614 15214 17666
rect 16146 17614 16158 17666
rect 16210 17614 16222 17666
rect 14030 17602 14082 17614
rect 17726 17602 17778 17614
rect 19742 17666 19794 17678
rect 19742 17602 19794 17614
rect 21982 17666 22034 17678
rect 21982 17602 22034 17614
rect 23326 17666 23378 17678
rect 25006 17666 25058 17678
rect 23874 17614 23886 17666
rect 23938 17614 23950 17666
rect 23326 17602 23378 17614
rect 25006 17602 25058 17614
rect 25342 17666 25394 17678
rect 25342 17602 25394 17614
rect 27358 17666 27410 17678
rect 27358 17602 27410 17614
rect 28254 17666 28306 17678
rect 28254 17602 28306 17614
rect 29822 17666 29874 17678
rect 29822 17602 29874 17614
rect 32734 17666 32786 17678
rect 32734 17602 32786 17614
rect 33518 17666 33570 17678
rect 35758 17666 35810 17678
rect 35298 17614 35310 17666
rect 35362 17614 35374 17666
rect 33518 17602 33570 17614
rect 35758 17602 35810 17614
rect 38110 17666 38162 17678
rect 38110 17602 38162 17614
rect 40574 17666 40626 17678
rect 40574 17602 40626 17614
rect 41918 17666 41970 17678
rect 44718 17666 44770 17678
rect 44258 17614 44270 17666
rect 44322 17614 44334 17666
rect 41918 17602 41970 17614
rect 44718 17602 44770 17614
rect 53454 17666 53506 17678
rect 53454 17602 53506 17614
rect 56478 17666 56530 17678
rect 56478 17602 56530 17614
rect 8542 17554 8594 17566
rect 19854 17554 19906 17566
rect 2034 17502 2046 17554
rect 2098 17502 2110 17554
rect 7522 17502 7534 17554
rect 7586 17502 7598 17554
rect 8306 17502 8318 17554
rect 8370 17502 8382 17554
rect 16482 17502 16494 17554
rect 16546 17502 16558 17554
rect 19170 17502 19182 17554
rect 19234 17502 19246 17554
rect 8542 17490 8594 17502
rect 19854 17490 19906 17502
rect 21646 17554 21698 17566
rect 21646 17490 21698 17502
rect 23214 17554 23266 17566
rect 23214 17490 23266 17502
rect 23438 17554 23490 17566
rect 23438 17490 23490 17502
rect 25118 17554 25170 17566
rect 25118 17490 25170 17502
rect 26238 17554 26290 17566
rect 26238 17490 26290 17502
rect 26462 17554 26514 17566
rect 26462 17490 26514 17502
rect 26574 17554 26626 17566
rect 26574 17490 26626 17502
rect 31166 17554 31218 17566
rect 31166 17490 31218 17502
rect 31278 17554 31330 17566
rect 31278 17490 31330 17502
rect 32062 17554 32114 17566
rect 32062 17490 32114 17502
rect 32286 17554 32338 17566
rect 32286 17490 32338 17502
rect 38446 17554 38498 17566
rect 38446 17490 38498 17502
rect 41022 17554 41074 17566
rect 41022 17490 41074 17502
rect 53790 17554 53842 17566
rect 53790 17490 53842 17502
rect 55694 17554 55746 17566
rect 55694 17490 55746 17502
rect 56254 17554 56306 17566
rect 57362 17502 57374 17554
rect 57426 17502 57438 17554
rect 56254 17490 56306 17502
rect 4174 17442 4226 17454
rect 4174 17378 4226 17390
rect 4622 17442 4674 17454
rect 4622 17378 4674 17390
rect 4958 17442 5010 17454
rect 4958 17378 5010 17390
rect 5966 17442 6018 17454
rect 5966 17378 6018 17390
rect 11342 17442 11394 17454
rect 11342 17378 11394 17390
rect 18846 17442 18898 17454
rect 18846 17378 18898 17390
rect 20078 17442 20130 17454
rect 20078 17378 20130 17390
rect 20862 17442 20914 17454
rect 20862 17378 20914 17390
rect 21758 17442 21810 17454
rect 21758 17378 21810 17390
rect 22542 17442 22594 17454
rect 22542 17378 22594 17390
rect 25678 17442 25730 17454
rect 25678 17378 25730 17390
rect 27246 17442 27298 17454
rect 27246 17378 27298 17390
rect 27918 17442 27970 17454
rect 27918 17378 27970 17390
rect 28814 17442 28866 17454
rect 28814 17378 28866 17390
rect 29486 17442 29538 17454
rect 29486 17378 29538 17390
rect 29710 17442 29762 17454
rect 29710 17378 29762 17390
rect 30494 17442 30546 17454
rect 30494 17378 30546 17390
rect 33182 17442 33234 17454
rect 33182 17378 33234 17390
rect 35422 17442 35474 17454
rect 35422 17378 35474 17390
rect 38334 17442 38386 17454
rect 38334 17378 38386 17390
rect 41246 17442 41298 17454
rect 41246 17378 41298 17390
rect 43374 17442 43426 17454
rect 45838 17442 45890 17454
rect 45490 17390 45502 17442
rect 45554 17390 45566 17442
rect 43374 17378 43426 17390
rect 45838 17378 45890 17390
rect 46286 17442 46338 17454
rect 48302 17442 48354 17454
rect 47954 17390 47966 17442
rect 48018 17390 48030 17442
rect 46286 17378 46338 17390
rect 48302 17378 48354 17390
rect 50430 17442 50482 17454
rect 50430 17378 50482 17390
rect 51326 17442 51378 17454
rect 51326 17378 51378 17390
rect 51774 17442 51826 17454
rect 51774 17378 51826 17390
rect 54574 17442 54626 17454
rect 55582 17442 55634 17454
rect 54898 17390 54910 17442
rect 54962 17390 54974 17442
rect 54574 17378 54626 17390
rect 55582 17378 55634 17390
rect 57710 17442 57762 17454
rect 57710 17378 57762 17390
rect 1344 17274 58576 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 58576 17274
rect 1344 17188 58576 17222
rect 2158 17106 2210 17118
rect 2158 17042 2210 17054
rect 2494 17106 2546 17118
rect 2494 17042 2546 17054
rect 2942 17106 2994 17118
rect 9102 17106 9154 17118
rect 11902 17106 11954 17118
rect 5618 17054 5630 17106
rect 5682 17054 5694 17106
rect 10098 17054 10110 17106
rect 10162 17054 10174 17106
rect 10994 17054 11006 17106
rect 11058 17054 11070 17106
rect 2942 17042 2994 17054
rect 9102 17042 9154 17054
rect 11902 17042 11954 17054
rect 15038 17106 15090 17118
rect 16606 17106 16658 17118
rect 15362 17054 15374 17106
rect 15426 17054 15438 17106
rect 15038 17042 15090 17054
rect 16606 17042 16658 17054
rect 17054 17106 17106 17118
rect 17054 17042 17106 17054
rect 18174 17106 18226 17118
rect 18174 17042 18226 17054
rect 20190 17106 20242 17118
rect 20190 17042 20242 17054
rect 25566 17106 25618 17118
rect 25566 17042 25618 17054
rect 28142 17106 28194 17118
rect 28142 17042 28194 17054
rect 28590 17106 28642 17118
rect 28590 17042 28642 17054
rect 29934 17106 29986 17118
rect 29934 17042 29986 17054
rect 30718 17106 30770 17118
rect 30718 17042 30770 17054
rect 31726 17106 31778 17118
rect 33966 17106 34018 17118
rect 32162 17054 32174 17106
rect 32226 17054 32238 17106
rect 31726 17042 31778 17054
rect 33966 17042 34018 17054
rect 34750 17106 34802 17118
rect 34750 17042 34802 17054
rect 36318 17106 36370 17118
rect 36318 17042 36370 17054
rect 36654 17106 36706 17118
rect 36654 17042 36706 17054
rect 37102 17106 37154 17118
rect 37102 17042 37154 17054
rect 37550 17106 37602 17118
rect 37550 17042 37602 17054
rect 39118 17106 39170 17118
rect 39118 17042 39170 17054
rect 41918 17106 41970 17118
rect 41918 17042 41970 17054
rect 42366 17106 42418 17118
rect 42366 17042 42418 17054
rect 43374 17106 43426 17118
rect 43374 17042 43426 17054
rect 44270 17106 44322 17118
rect 51998 17106 52050 17118
rect 54910 17106 54962 17118
rect 45714 17054 45726 17106
rect 45778 17054 45790 17106
rect 46834 17054 46846 17106
rect 46898 17054 46910 17106
rect 53554 17054 53566 17106
rect 53618 17054 53630 17106
rect 44270 17042 44322 17054
rect 51998 17042 52050 17054
rect 54910 17042 54962 17054
rect 56702 17106 56754 17118
rect 56702 17042 56754 17054
rect 6974 16994 7026 17006
rect 4386 16942 4398 16994
rect 4450 16942 4462 16994
rect 5730 16942 5742 16994
rect 5794 16942 5806 16994
rect 6066 16942 6078 16994
rect 6130 16942 6142 16994
rect 6974 16930 7026 16942
rect 7310 16994 7362 17006
rect 7310 16930 7362 16942
rect 12238 16994 12290 17006
rect 12238 16930 12290 16942
rect 13582 16994 13634 17006
rect 13582 16930 13634 16942
rect 14478 16994 14530 17006
rect 14478 16930 14530 16942
rect 17726 16994 17778 17006
rect 17726 16930 17778 16942
rect 19966 16994 20018 17006
rect 19966 16930 20018 16942
rect 26574 16994 26626 17006
rect 26574 16930 26626 16942
rect 29150 16994 29202 17006
rect 29150 16930 29202 16942
rect 34414 16994 34466 17006
rect 34414 16930 34466 16942
rect 35534 16994 35586 17006
rect 35534 16930 35586 16942
rect 45390 16994 45442 17006
rect 51550 16994 51602 17006
rect 47842 16942 47854 16994
rect 47906 16942 47918 16994
rect 49634 16942 49646 16994
rect 49698 16942 49710 16994
rect 45390 16930 45442 16942
rect 51550 16930 51602 16942
rect 54462 16994 54514 17006
rect 54462 16930 54514 16942
rect 54686 16994 54738 17006
rect 54686 16930 54738 16942
rect 55918 16994 55970 17006
rect 57474 16942 57486 16994
rect 57538 16942 57550 16994
rect 55918 16930 55970 16942
rect 3390 16882 3442 16894
rect 7198 16882 7250 16894
rect 4610 16830 4622 16882
rect 4674 16830 4686 16882
rect 6402 16830 6414 16882
rect 6466 16830 6478 16882
rect 3390 16818 3442 16830
rect 7198 16818 7250 16830
rect 8654 16882 8706 16894
rect 8654 16818 8706 16830
rect 9774 16882 9826 16894
rect 9774 16818 9826 16830
rect 10670 16882 10722 16894
rect 10670 16818 10722 16830
rect 12798 16882 12850 16894
rect 18846 16882 18898 16894
rect 20750 16882 20802 16894
rect 13234 16830 13246 16882
rect 13298 16830 13310 16882
rect 13906 16830 13918 16882
rect 13970 16830 13982 16882
rect 17938 16830 17950 16882
rect 18002 16830 18014 16882
rect 19394 16830 19406 16882
rect 19458 16830 19470 16882
rect 19730 16830 19742 16882
rect 19794 16830 19806 16882
rect 12798 16818 12850 16830
rect 18846 16818 18898 16830
rect 20750 16818 20802 16830
rect 21310 16882 21362 16894
rect 21310 16818 21362 16830
rect 21646 16882 21698 16894
rect 21646 16818 21698 16830
rect 21870 16882 21922 16894
rect 23102 16882 23154 16894
rect 26462 16882 26514 16894
rect 22642 16830 22654 16882
rect 22706 16830 22718 16882
rect 23762 16830 23774 16882
rect 23826 16830 23838 16882
rect 21870 16818 21922 16830
rect 23102 16818 23154 16830
rect 26462 16818 26514 16830
rect 27694 16882 27746 16894
rect 27694 16818 27746 16830
rect 29486 16882 29538 16894
rect 29486 16818 29538 16830
rect 32510 16882 32562 16894
rect 32510 16818 32562 16830
rect 32734 16882 32786 16894
rect 32734 16818 32786 16830
rect 35646 16882 35698 16894
rect 35646 16818 35698 16830
rect 36094 16882 36146 16894
rect 36094 16818 36146 16830
rect 37998 16882 38050 16894
rect 40350 16882 40402 16894
rect 38882 16830 38894 16882
rect 38946 16830 38958 16882
rect 40002 16830 40014 16882
rect 40066 16830 40078 16882
rect 37998 16818 38050 16830
rect 40350 16818 40402 16830
rect 41470 16882 41522 16894
rect 41470 16818 41522 16830
rect 42814 16882 42866 16894
rect 42814 16818 42866 16830
rect 44606 16882 44658 16894
rect 44606 16818 44658 16830
rect 46174 16882 46226 16894
rect 46174 16818 46226 16830
rect 47182 16882 47234 16894
rect 47182 16818 47234 16830
rect 48190 16882 48242 16894
rect 48190 16818 48242 16830
rect 48414 16882 48466 16894
rect 55022 16882 55074 16894
rect 49970 16830 49982 16882
rect 50034 16830 50046 16882
rect 50530 16830 50542 16882
rect 50594 16830 50606 16882
rect 52994 16830 53006 16882
rect 53058 16830 53070 16882
rect 53218 16830 53230 16882
rect 53282 16830 53294 16882
rect 48414 16818 48466 16830
rect 55022 16818 55074 16830
rect 56254 16882 56306 16894
rect 57698 16830 57710 16882
rect 57762 16830 57774 16882
rect 56254 16818 56306 16830
rect 3950 16770 4002 16782
rect 3950 16706 4002 16718
rect 7534 16770 7586 16782
rect 7534 16706 7586 16718
rect 16046 16770 16098 16782
rect 16046 16706 16098 16718
rect 18286 16770 18338 16782
rect 21422 16770 21474 16782
rect 24894 16770 24946 16782
rect 19842 16718 19854 16770
rect 19906 16718 19918 16770
rect 23650 16718 23662 16770
rect 23714 16718 23726 16770
rect 18286 16706 18338 16718
rect 21422 16706 21474 16718
rect 24894 16706 24946 16718
rect 27358 16770 27410 16782
rect 27358 16706 27410 16718
rect 35310 16770 35362 16782
rect 35310 16706 35362 16718
rect 40574 16770 40626 16782
rect 50318 16770 50370 16782
rect 49746 16718 49758 16770
rect 49810 16718 49822 16770
rect 53554 16718 53566 16770
rect 53618 16718 53630 16770
rect 40574 16706 40626 16718
rect 50318 16706 50370 16718
rect 7758 16658 7810 16670
rect 26574 16658 26626 16670
rect 2146 16606 2158 16658
rect 2210 16655 2222 16658
rect 2930 16655 2942 16658
rect 2210 16609 2942 16655
rect 2210 16606 2222 16609
rect 2930 16606 2942 16609
rect 2994 16606 3006 16658
rect 23426 16606 23438 16658
rect 23490 16606 23502 16658
rect 7758 16594 7810 16606
rect 26574 16594 26626 16606
rect 1344 16490 58576 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 58576 16490
rect 1344 16404 58576 16438
rect 23774 16322 23826 16334
rect 12114 16270 12126 16322
rect 12178 16319 12190 16322
rect 12562 16319 12574 16322
rect 12178 16273 12574 16319
rect 12178 16270 12190 16273
rect 12562 16270 12574 16273
rect 12626 16270 12638 16322
rect 23774 16258 23826 16270
rect 33630 16322 33682 16334
rect 33630 16258 33682 16270
rect 40910 16322 40962 16334
rect 40910 16258 40962 16270
rect 41022 16322 41074 16334
rect 41022 16258 41074 16270
rect 41358 16322 41410 16334
rect 45490 16270 45502 16322
rect 45554 16270 45566 16322
rect 54114 16270 54126 16322
rect 54178 16270 54190 16322
rect 41358 16258 41410 16270
rect 3278 16210 3330 16222
rect 3278 16146 3330 16158
rect 3614 16210 3666 16222
rect 3614 16146 3666 16158
rect 4622 16210 4674 16222
rect 4622 16146 4674 16158
rect 6526 16210 6578 16222
rect 8430 16210 8482 16222
rect 7858 16158 7870 16210
rect 7922 16158 7934 16210
rect 6526 16146 6578 16158
rect 8430 16146 8482 16158
rect 10334 16210 10386 16222
rect 10334 16146 10386 16158
rect 12910 16210 12962 16222
rect 12910 16146 12962 16158
rect 14478 16210 14530 16222
rect 14478 16146 14530 16158
rect 15374 16210 15426 16222
rect 20974 16210 21026 16222
rect 17490 16158 17502 16210
rect 17554 16158 17566 16210
rect 18162 16158 18174 16210
rect 18226 16158 18238 16210
rect 15374 16146 15426 16158
rect 20974 16146 21026 16158
rect 23214 16210 23266 16222
rect 23214 16146 23266 16158
rect 26126 16210 26178 16222
rect 26126 16146 26178 16158
rect 27022 16210 27074 16222
rect 28814 16210 28866 16222
rect 28242 16158 28254 16210
rect 28306 16158 28318 16210
rect 27022 16146 27074 16158
rect 28814 16146 28866 16158
rect 30830 16210 30882 16222
rect 30830 16146 30882 16158
rect 33518 16210 33570 16222
rect 33518 16146 33570 16158
rect 34526 16210 34578 16222
rect 34526 16146 34578 16158
rect 35534 16210 35586 16222
rect 35534 16146 35586 16158
rect 44158 16210 44210 16222
rect 44158 16146 44210 16158
rect 44494 16210 44546 16222
rect 44494 16146 44546 16158
rect 48302 16210 48354 16222
rect 48302 16146 48354 16158
rect 50206 16210 50258 16222
rect 54686 16210 54738 16222
rect 52210 16158 52222 16210
rect 52274 16158 52286 16210
rect 50206 16146 50258 16158
rect 54686 16146 54738 16158
rect 57374 16210 57426 16222
rect 57374 16146 57426 16158
rect 4174 16098 4226 16110
rect 4174 16034 4226 16046
rect 5070 16098 5122 16110
rect 11118 16098 11170 16110
rect 19070 16098 19122 16110
rect 9538 16046 9550 16098
rect 9602 16046 9614 16098
rect 15810 16046 15822 16098
rect 15874 16046 15886 16098
rect 16034 16046 16046 16098
rect 16098 16046 16110 16098
rect 17042 16046 17054 16098
rect 17106 16046 17118 16098
rect 18274 16046 18286 16098
rect 18338 16046 18350 16098
rect 5070 16034 5122 16046
rect 11118 16034 11170 16046
rect 19070 16034 19122 16046
rect 20526 16098 20578 16110
rect 24558 16098 24610 16110
rect 23426 16046 23438 16098
rect 23490 16046 23502 16098
rect 20526 16034 20578 16046
rect 24558 16034 24610 16046
rect 25118 16098 25170 16110
rect 25118 16034 25170 16046
rect 26350 16098 26402 16110
rect 26350 16034 26402 16046
rect 26574 16098 26626 16110
rect 29934 16098 29986 16110
rect 27906 16046 27918 16098
rect 27970 16046 27982 16098
rect 26574 16034 26626 16046
rect 29934 16034 29986 16046
rect 30382 16098 30434 16110
rect 30382 16034 30434 16046
rect 32062 16098 32114 16110
rect 32062 16034 32114 16046
rect 35086 16098 35138 16110
rect 35086 16034 35138 16046
rect 35310 16098 35362 16110
rect 35310 16034 35362 16046
rect 35758 16098 35810 16110
rect 35758 16034 35810 16046
rect 37998 16098 38050 16110
rect 37998 16034 38050 16046
rect 38110 16098 38162 16110
rect 39118 16098 39170 16110
rect 38434 16046 38446 16098
rect 38498 16046 38510 16098
rect 38110 16034 38162 16046
rect 39118 16034 39170 16046
rect 41246 16098 41298 16110
rect 43598 16098 43650 16110
rect 42242 16046 42254 16098
rect 42306 16046 42318 16098
rect 41246 16034 41298 16046
rect 43598 16034 43650 16046
rect 45838 16098 45890 16110
rect 45838 16034 45890 16046
rect 46062 16098 46114 16110
rect 49646 16098 49698 16110
rect 47618 16046 47630 16098
rect 47682 16046 47694 16098
rect 49298 16046 49310 16098
rect 49362 16046 49374 16098
rect 46062 16034 46114 16046
rect 49646 16034 49698 16046
rect 50766 16098 50818 16110
rect 55806 16098 55858 16110
rect 51202 16046 51214 16098
rect 51266 16046 51278 16098
rect 52098 16046 52110 16098
rect 52162 16046 52174 16098
rect 53666 16046 53678 16098
rect 53730 16046 53742 16098
rect 54114 16046 54126 16098
rect 54178 16046 54190 16098
rect 55458 16046 55470 16098
rect 55522 16046 55534 16098
rect 50766 16034 50818 16046
rect 55806 16034 55858 16046
rect 7310 15986 7362 15998
rect 5730 15934 5742 15986
rect 5794 15934 5806 15986
rect 7310 15922 7362 15934
rect 7422 15986 7474 15998
rect 13918 15986 13970 15998
rect 7522 15934 7534 15986
rect 7586 15934 7598 15986
rect 9314 15934 9326 15986
rect 9378 15934 9390 15986
rect 7422 15922 7474 15934
rect 13918 15922 13970 15934
rect 16270 15986 16322 15998
rect 16270 15922 16322 15934
rect 16382 15986 16434 15998
rect 16382 15922 16434 15934
rect 17838 15986 17890 15998
rect 17838 15922 17890 15934
rect 21758 15986 21810 15998
rect 21758 15922 21810 15934
rect 21982 15986 22034 15998
rect 21982 15922 22034 15934
rect 22318 15986 22370 15998
rect 22318 15922 22370 15934
rect 25454 15986 25506 15998
rect 25454 15922 25506 15934
rect 26014 15986 26066 15998
rect 26014 15922 26066 15934
rect 29598 15986 29650 15998
rect 29598 15922 29650 15934
rect 31950 15986 32002 15998
rect 31950 15922 32002 15934
rect 32622 15986 32674 15998
rect 32622 15922 32674 15934
rect 32958 15986 33010 15998
rect 32958 15922 33010 15934
rect 34078 15986 34130 15998
rect 34078 15922 34130 15934
rect 36318 15986 36370 15998
rect 36318 15922 36370 15934
rect 36430 15986 36482 15998
rect 36430 15922 36482 15934
rect 36654 15986 36706 15998
rect 36654 15922 36706 15934
rect 37662 15986 37714 15998
rect 37662 15922 37714 15934
rect 39454 15986 39506 15998
rect 39454 15922 39506 15934
rect 42030 15986 42082 15998
rect 42030 15922 42082 15934
rect 46622 15986 46674 15998
rect 46622 15922 46674 15934
rect 46958 15986 47010 15998
rect 47842 15934 47854 15986
rect 47906 15934 47918 15986
rect 52546 15934 52558 15986
rect 52610 15934 52622 15986
rect 56578 15934 56590 15986
rect 56642 15934 56654 15986
rect 46958 15922 47010 15934
rect 1934 15874 1986 15886
rect 1934 15810 1986 15822
rect 2382 15874 2434 15886
rect 2382 15810 2434 15822
rect 2830 15874 2882 15886
rect 2830 15810 2882 15822
rect 6078 15874 6130 15886
rect 6078 15810 6130 15822
rect 7086 15874 7138 15886
rect 7086 15810 7138 15822
rect 8878 15874 8930 15886
rect 8878 15810 8930 15822
rect 10894 15874 10946 15886
rect 10894 15810 10946 15822
rect 11006 15874 11058 15886
rect 11006 15810 11058 15822
rect 11342 15874 11394 15886
rect 11342 15810 11394 15822
rect 12014 15874 12066 15886
rect 12014 15810 12066 15822
rect 12574 15874 12626 15886
rect 12574 15810 12626 15822
rect 13582 15874 13634 15886
rect 13582 15810 13634 15822
rect 13806 15874 13858 15886
rect 13806 15810 13858 15822
rect 19182 15874 19234 15886
rect 19182 15810 19234 15822
rect 19294 15874 19346 15886
rect 19294 15810 19346 15822
rect 19518 15874 19570 15886
rect 19518 15810 19570 15822
rect 22094 15874 22146 15886
rect 22094 15810 22146 15822
rect 23102 15874 23154 15886
rect 23102 15810 23154 15822
rect 23326 15874 23378 15886
rect 23326 15810 23378 15822
rect 31278 15874 31330 15886
rect 31278 15810 31330 15822
rect 31726 15874 31778 15886
rect 31726 15810 31778 15822
rect 37774 15874 37826 15886
rect 37774 15810 37826 15822
rect 39902 15874 39954 15886
rect 39902 15810 39954 15822
rect 43262 15874 43314 15886
rect 43262 15810 43314 15822
rect 48974 15874 49026 15886
rect 48974 15810 49026 15822
rect 49086 15874 49138 15886
rect 49086 15810 49138 15822
rect 50094 15874 50146 15886
rect 50094 15810 50146 15822
rect 50318 15874 50370 15886
rect 50318 15810 50370 15822
rect 55358 15874 55410 15886
rect 55358 15810 55410 15822
rect 56926 15874 56978 15886
rect 56926 15810 56978 15822
rect 57822 15874 57874 15886
rect 57822 15810 57874 15822
rect 1344 15706 58576 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 58576 15706
rect 1344 15620 58576 15654
rect 2158 15538 2210 15550
rect 2158 15474 2210 15486
rect 2606 15538 2658 15550
rect 5406 15538 5458 15550
rect 8654 15538 8706 15550
rect 3378 15486 3390 15538
rect 3442 15486 3454 15538
rect 3938 15486 3950 15538
rect 4002 15486 4014 15538
rect 6738 15486 6750 15538
rect 6802 15486 6814 15538
rect 2606 15474 2658 15486
rect 5406 15474 5458 15486
rect 8654 15474 8706 15486
rect 9662 15538 9714 15550
rect 9662 15474 9714 15486
rect 11454 15538 11506 15550
rect 16158 15538 16210 15550
rect 13010 15486 13022 15538
rect 13074 15486 13086 15538
rect 11454 15474 11506 15486
rect 16158 15474 16210 15486
rect 16942 15538 16994 15550
rect 16942 15474 16994 15486
rect 18174 15538 18226 15550
rect 18174 15474 18226 15486
rect 22430 15538 22482 15550
rect 22430 15474 22482 15486
rect 22990 15538 23042 15550
rect 22990 15474 23042 15486
rect 23774 15538 23826 15550
rect 23774 15474 23826 15486
rect 24558 15538 24610 15550
rect 24558 15474 24610 15486
rect 24782 15538 24834 15550
rect 24782 15474 24834 15486
rect 25790 15538 25842 15550
rect 25790 15474 25842 15486
rect 28030 15538 28082 15550
rect 28030 15474 28082 15486
rect 29262 15538 29314 15550
rect 29262 15474 29314 15486
rect 29934 15538 29986 15550
rect 29934 15474 29986 15486
rect 31726 15538 31778 15550
rect 31726 15474 31778 15486
rect 32510 15538 32562 15550
rect 32510 15474 32562 15486
rect 33742 15538 33794 15550
rect 33742 15474 33794 15486
rect 34302 15538 34354 15550
rect 34302 15474 34354 15486
rect 34862 15538 34914 15550
rect 34862 15474 34914 15486
rect 35422 15538 35474 15550
rect 35422 15474 35474 15486
rect 36206 15538 36258 15550
rect 36206 15474 36258 15486
rect 36990 15538 37042 15550
rect 36990 15474 37042 15486
rect 38110 15538 38162 15550
rect 38110 15474 38162 15486
rect 38670 15538 38722 15550
rect 38670 15474 38722 15486
rect 39230 15538 39282 15550
rect 39230 15474 39282 15486
rect 39566 15538 39618 15550
rect 39566 15474 39618 15486
rect 40014 15538 40066 15550
rect 40014 15474 40066 15486
rect 40686 15538 40738 15550
rect 40686 15474 40738 15486
rect 41582 15538 41634 15550
rect 41582 15474 41634 15486
rect 44382 15538 44434 15550
rect 44382 15474 44434 15486
rect 45054 15538 45106 15550
rect 45054 15474 45106 15486
rect 45950 15538 46002 15550
rect 46846 15538 46898 15550
rect 46274 15486 46286 15538
rect 46338 15486 46350 15538
rect 45950 15474 46002 15486
rect 46846 15474 46898 15486
rect 51326 15538 51378 15550
rect 53790 15538 53842 15550
rect 51874 15486 51886 15538
rect 51938 15486 51950 15538
rect 53330 15486 53342 15538
rect 53394 15486 53406 15538
rect 51326 15474 51378 15486
rect 53790 15474 53842 15486
rect 54574 15538 54626 15550
rect 54574 15474 54626 15486
rect 56590 15538 56642 15550
rect 56590 15474 56642 15486
rect 57486 15538 57538 15550
rect 57486 15474 57538 15486
rect 9886 15426 9938 15438
rect 9886 15362 9938 15374
rect 10558 15426 10610 15438
rect 10558 15362 10610 15374
rect 10782 15426 10834 15438
rect 10782 15362 10834 15374
rect 16046 15426 16098 15438
rect 16046 15362 16098 15374
rect 16382 15426 16434 15438
rect 16382 15362 16434 15374
rect 17950 15426 18002 15438
rect 26462 15426 26514 15438
rect 21634 15374 21646 15426
rect 21698 15374 21710 15426
rect 17950 15362 18002 15374
rect 26462 15362 26514 15374
rect 26686 15426 26738 15438
rect 26686 15362 26738 15374
rect 33854 15426 33906 15438
rect 33854 15362 33906 15374
rect 35870 15426 35922 15438
rect 35870 15362 35922 15374
rect 37886 15426 37938 15438
rect 42366 15426 42418 15438
rect 42130 15374 42142 15426
rect 42194 15374 42206 15426
rect 37886 15362 37938 15374
rect 42366 15362 42418 15374
rect 45390 15426 45442 15438
rect 45390 15362 45442 15374
rect 46958 15426 47010 15438
rect 46958 15362 47010 15374
rect 48190 15426 48242 15438
rect 48190 15362 48242 15374
rect 48526 15426 48578 15438
rect 48526 15362 48578 15374
rect 53006 15426 53058 15438
rect 53006 15362 53058 15374
rect 54686 15426 54738 15438
rect 54686 15362 54738 15374
rect 54910 15426 54962 15438
rect 54910 15362 54962 15374
rect 55470 15426 55522 15438
rect 55470 15362 55522 15374
rect 3054 15314 3106 15326
rect 4846 15314 4898 15326
rect 4162 15262 4174 15314
rect 4226 15262 4238 15314
rect 3054 15250 3106 15262
rect 4846 15250 4898 15262
rect 5742 15314 5794 15326
rect 8094 15314 8146 15326
rect 6850 15262 6862 15314
rect 6914 15262 6926 15314
rect 7186 15262 7198 15314
rect 7250 15262 7262 15314
rect 5742 15250 5794 15262
rect 8094 15250 8146 15262
rect 9998 15314 10050 15326
rect 13694 15314 13746 15326
rect 15934 15314 15986 15326
rect 12338 15262 12350 15314
rect 12402 15262 12414 15314
rect 12898 15262 12910 15314
rect 12962 15262 12974 15314
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 15026 15262 15038 15314
rect 15090 15262 15102 15314
rect 9998 15250 10050 15262
rect 13694 15250 13746 15262
rect 15934 15250 15986 15262
rect 18398 15314 18450 15326
rect 18398 15250 18450 15262
rect 18510 15314 18562 15326
rect 23326 15314 23378 15326
rect 19506 15262 19518 15314
rect 19570 15262 19582 15314
rect 19842 15262 19854 15314
rect 19906 15262 19918 15314
rect 20514 15262 20526 15314
rect 20578 15262 20590 15314
rect 21074 15262 21086 15314
rect 21138 15262 21150 15314
rect 18510 15250 18562 15262
rect 23326 15250 23378 15262
rect 24894 15314 24946 15326
rect 24894 15250 24946 15262
rect 27246 15314 27298 15326
rect 28814 15314 28866 15326
rect 27794 15262 27806 15314
rect 27858 15262 27870 15314
rect 27246 15250 27298 15262
rect 28814 15250 28866 15262
rect 30158 15314 30210 15326
rect 30158 15250 30210 15262
rect 30382 15314 30434 15326
rect 30382 15250 30434 15262
rect 30606 15314 30658 15326
rect 30606 15250 30658 15262
rect 32286 15314 32338 15326
rect 32286 15250 32338 15262
rect 32958 15314 33010 15326
rect 32958 15250 33010 15262
rect 33518 15314 33570 15326
rect 33518 15250 33570 15262
rect 36094 15314 36146 15326
rect 36094 15250 36146 15262
rect 36542 15314 36594 15326
rect 37998 15314 38050 15326
rect 37202 15262 37214 15314
rect 37266 15262 37278 15314
rect 36542 15250 36594 15262
rect 37998 15250 38050 15262
rect 42030 15314 42082 15326
rect 43486 15314 43538 15326
rect 42690 15262 42702 15314
rect 42754 15262 42766 15314
rect 42030 15250 42082 15262
rect 43486 15250 43538 15262
rect 43710 15314 43762 15326
rect 52222 15314 52274 15326
rect 50418 15262 50430 15314
rect 50482 15262 50494 15314
rect 43710 15250 43762 15262
rect 52222 15250 52274 15262
rect 54238 15314 54290 15326
rect 54238 15250 54290 15262
rect 55918 15314 55970 15326
rect 57698 15262 57710 15314
rect 57762 15262 57774 15314
rect 55918 15250 55970 15262
rect 8990 15202 9042 15214
rect 7298 15150 7310 15202
rect 7362 15150 7374 15202
rect 8990 15138 9042 15150
rect 11118 15202 11170 15214
rect 11118 15138 11170 15150
rect 12014 15202 12066 15214
rect 31278 15202 31330 15214
rect 20962 15150 20974 15202
rect 21026 15150 21038 15202
rect 26338 15150 26350 15202
rect 26402 15150 26414 15202
rect 30034 15150 30046 15202
rect 30098 15150 30110 15202
rect 12014 15138 12066 15150
rect 31278 15138 31330 15150
rect 32398 15202 32450 15214
rect 32398 15138 32450 15150
rect 43038 15202 43090 15214
rect 43038 15138 43090 15150
rect 43934 15202 43986 15214
rect 43934 15138 43986 15150
rect 47406 15202 47458 15214
rect 47406 15138 47458 15150
rect 49422 15202 49474 15214
rect 50878 15202 50930 15214
rect 50194 15150 50206 15202
rect 50258 15150 50270 15202
rect 49422 15138 49474 15150
rect 50878 15138 50930 15150
rect 52446 15202 52498 15214
rect 52446 15138 52498 15150
rect 56142 15202 56194 15214
rect 56142 15138 56194 15150
rect 11342 15090 11394 15102
rect 11342 15026 11394 15038
rect 18062 15090 18114 15102
rect 30830 15090 30882 15102
rect 25554 15038 25566 15090
rect 25618 15087 25630 15090
rect 26114 15087 26126 15090
rect 25618 15041 26126 15087
rect 25618 15038 25630 15041
rect 26114 15038 26126 15041
rect 26178 15038 26190 15090
rect 18062 15026 18114 15038
rect 30830 15026 30882 15038
rect 55694 15090 55746 15102
rect 55694 15026 55746 15038
rect 1344 14922 58576 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 58576 14922
rect 1344 14836 58576 14870
rect 9550 14754 9602 14766
rect 1810 14702 1822 14754
rect 1874 14751 1886 14754
rect 2258 14751 2270 14754
rect 1874 14705 2270 14751
rect 1874 14702 1886 14705
rect 2258 14702 2270 14705
rect 2322 14702 2334 14754
rect 4162 14702 4174 14754
rect 4226 14751 4238 14754
rect 4946 14751 4958 14754
rect 4226 14705 4958 14751
rect 4226 14702 4238 14705
rect 4946 14702 4958 14705
rect 5010 14702 5022 14754
rect 9550 14690 9602 14702
rect 12126 14754 12178 14766
rect 12126 14690 12178 14702
rect 12910 14754 12962 14766
rect 26238 14754 26290 14766
rect 17042 14702 17054 14754
rect 17106 14751 17118 14754
rect 17378 14751 17390 14754
rect 17106 14705 17390 14751
rect 17106 14702 17118 14705
rect 17378 14702 17390 14705
rect 17442 14702 17454 14754
rect 20402 14702 20414 14754
rect 20466 14751 20478 14754
rect 20962 14751 20974 14754
rect 20466 14705 20974 14751
rect 20466 14702 20478 14705
rect 20962 14702 20974 14705
rect 21026 14702 21038 14754
rect 12910 14690 12962 14702
rect 26238 14690 26290 14702
rect 36094 14754 36146 14766
rect 45938 14702 45950 14754
rect 46002 14751 46014 14754
rect 46274 14751 46286 14754
rect 46002 14705 46286 14751
rect 46002 14702 46014 14705
rect 46274 14702 46286 14705
rect 46338 14702 46350 14754
rect 47842 14702 47854 14754
rect 47906 14751 47918 14754
rect 48066 14751 48078 14754
rect 47906 14705 48078 14751
rect 47906 14702 47918 14705
rect 48066 14702 48078 14705
rect 48130 14702 48142 14754
rect 36094 14690 36146 14702
rect 1934 14642 1986 14654
rect 1934 14578 1986 14590
rect 3614 14642 3666 14654
rect 3614 14578 3666 14590
rect 4062 14642 4114 14654
rect 4062 14578 4114 14590
rect 5854 14642 5906 14654
rect 5854 14578 5906 14590
rect 7646 14642 7698 14654
rect 7646 14578 7698 14590
rect 15598 14642 15650 14654
rect 15598 14578 15650 14590
rect 17054 14642 17106 14654
rect 17054 14578 17106 14590
rect 18062 14642 18114 14654
rect 18062 14578 18114 14590
rect 19070 14642 19122 14654
rect 19070 14578 19122 14590
rect 19854 14642 19906 14654
rect 19854 14578 19906 14590
rect 21870 14642 21922 14654
rect 21870 14578 21922 14590
rect 23102 14642 23154 14654
rect 23102 14578 23154 14590
rect 25230 14642 25282 14654
rect 25230 14578 25282 14590
rect 29598 14642 29650 14654
rect 29598 14578 29650 14590
rect 30270 14642 30322 14654
rect 30270 14578 30322 14590
rect 31278 14642 31330 14654
rect 31278 14578 31330 14590
rect 34638 14642 34690 14654
rect 34638 14578 34690 14590
rect 38446 14642 38498 14654
rect 38446 14578 38498 14590
rect 39790 14642 39842 14654
rect 39790 14578 39842 14590
rect 41246 14642 41298 14654
rect 47182 14642 47234 14654
rect 42914 14590 42926 14642
rect 42978 14590 42990 14642
rect 41246 14578 41298 14590
rect 47182 14578 47234 14590
rect 48190 14642 48242 14654
rect 48190 14578 48242 14590
rect 48750 14642 48802 14654
rect 48750 14578 48802 14590
rect 50318 14642 50370 14654
rect 50318 14578 50370 14590
rect 51102 14642 51154 14654
rect 52210 14590 52222 14642
rect 52274 14590 52286 14642
rect 55346 14590 55358 14642
rect 55410 14590 55422 14642
rect 51102 14578 51154 14590
rect 4510 14530 4562 14542
rect 4510 14466 4562 14478
rect 6862 14530 6914 14542
rect 6862 14466 6914 14478
rect 7758 14530 7810 14542
rect 7758 14466 7810 14478
rect 8654 14530 8706 14542
rect 8654 14466 8706 14478
rect 9102 14530 9154 14542
rect 9102 14466 9154 14478
rect 9326 14530 9378 14542
rect 11454 14530 11506 14542
rect 13694 14530 13746 14542
rect 10322 14478 10334 14530
rect 10386 14478 10398 14530
rect 11778 14478 11790 14530
rect 11842 14478 11854 14530
rect 12898 14478 12910 14530
rect 12962 14478 12974 14530
rect 9326 14466 9378 14478
rect 11454 14466 11506 14478
rect 13694 14466 13746 14478
rect 17390 14530 17442 14542
rect 17390 14466 17442 14478
rect 19630 14530 19682 14542
rect 30046 14530 30098 14542
rect 23762 14478 23774 14530
rect 23826 14478 23838 14530
rect 19630 14466 19682 14478
rect 30046 14466 30098 14478
rect 35534 14530 35586 14542
rect 35534 14466 35586 14478
rect 35982 14530 36034 14542
rect 35982 14466 36034 14478
rect 36318 14530 36370 14542
rect 36318 14466 36370 14478
rect 40462 14530 40514 14542
rect 57934 14530 57986 14542
rect 43138 14478 43150 14530
rect 43202 14478 43214 14530
rect 52322 14478 52334 14530
rect 52386 14478 52398 14530
rect 56018 14478 56030 14530
rect 56082 14478 56094 14530
rect 40462 14466 40514 14478
rect 57934 14466 57986 14478
rect 6414 14418 6466 14430
rect 6414 14354 6466 14366
rect 6638 14418 6690 14430
rect 6638 14354 6690 14366
rect 6974 14418 7026 14430
rect 6974 14354 7026 14366
rect 7534 14418 7586 14430
rect 7534 14354 7586 14366
rect 8094 14418 8146 14430
rect 8094 14354 8146 14366
rect 9774 14418 9826 14430
rect 12014 14418 12066 14430
rect 10434 14366 10446 14418
rect 10498 14366 10510 14418
rect 10994 14366 11006 14418
rect 11058 14366 11070 14418
rect 9774 14354 9826 14366
rect 12014 14354 12066 14366
rect 12574 14418 12626 14430
rect 16046 14418 16098 14430
rect 13906 14366 13918 14418
rect 13970 14366 13982 14418
rect 14466 14366 14478 14418
rect 14530 14366 14542 14418
rect 12574 14354 12626 14366
rect 16046 14354 16098 14366
rect 18734 14418 18786 14430
rect 18734 14354 18786 14366
rect 20078 14418 20130 14430
rect 20078 14354 20130 14366
rect 20302 14418 20354 14430
rect 20302 14354 20354 14366
rect 23326 14418 23378 14430
rect 25566 14418 25618 14430
rect 24658 14366 24670 14418
rect 24722 14366 24734 14418
rect 23326 14354 23378 14366
rect 25566 14354 25618 14366
rect 26574 14418 26626 14430
rect 36542 14418 36594 14430
rect 28802 14366 28814 14418
rect 28866 14366 28878 14418
rect 26574 14354 26626 14366
rect 36542 14354 36594 14366
rect 37550 14418 37602 14430
rect 37550 14354 37602 14366
rect 37886 14418 37938 14430
rect 37886 14354 37938 14366
rect 39006 14418 39058 14430
rect 39006 14354 39058 14366
rect 41694 14418 41746 14430
rect 41694 14354 41746 14366
rect 42478 14418 42530 14430
rect 42478 14354 42530 14366
rect 42926 14418 42978 14430
rect 42926 14354 42978 14366
rect 43710 14418 43762 14430
rect 43710 14354 43762 14366
rect 44046 14418 44098 14430
rect 44046 14354 44098 14366
rect 45502 14418 45554 14430
rect 45502 14354 45554 14366
rect 45614 14418 45666 14430
rect 45614 14354 45666 14366
rect 49422 14418 49474 14430
rect 51774 14418 51826 14430
rect 51314 14366 51326 14418
rect 51378 14415 51390 14418
rect 51650 14415 51662 14418
rect 51378 14369 51662 14415
rect 51378 14366 51390 14369
rect 51650 14366 51662 14369
rect 51714 14366 51726 14418
rect 49422 14354 49474 14366
rect 51774 14354 51826 14366
rect 53902 14418 53954 14430
rect 53902 14354 53954 14366
rect 56702 14418 56754 14430
rect 56702 14354 56754 14366
rect 57038 14418 57090 14430
rect 57038 14354 57090 14366
rect 57598 14418 57650 14430
rect 57598 14354 57650 14366
rect 2382 14306 2434 14318
rect 2382 14242 2434 14254
rect 2830 14306 2882 14318
rect 2830 14242 2882 14254
rect 3278 14306 3330 14318
rect 3278 14242 3330 14254
rect 4958 14306 5010 14318
rect 16382 14306 16434 14318
rect 13794 14254 13806 14306
rect 13858 14254 13870 14306
rect 4958 14242 5010 14254
rect 16382 14242 16434 14254
rect 18958 14306 19010 14318
rect 18958 14242 19010 14254
rect 19182 14306 19234 14318
rect 19182 14242 19234 14254
rect 20862 14306 20914 14318
rect 20862 14242 20914 14254
rect 22430 14306 22482 14318
rect 22430 14242 22482 14254
rect 22990 14306 23042 14318
rect 22990 14242 23042 14254
rect 23214 14306 23266 14318
rect 23214 14242 23266 14254
rect 24334 14306 24386 14318
rect 24334 14242 24386 14254
rect 26350 14306 26402 14318
rect 26350 14242 26402 14254
rect 27022 14306 27074 14318
rect 27918 14306 27970 14318
rect 27570 14254 27582 14306
rect 27634 14254 27646 14306
rect 27022 14242 27074 14254
rect 27918 14242 27970 14254
rect 28478 14306 28530 14318
rect 28478 14242 28530 14254
rect 30494 14306 30546 14318
rect 30494 14242 30546 14254
rect 30606 14306 30658 14318
rect 30606 14242 30658 14254
rect 30718 14306 30770 14318
rect 30718 14242 30770 14254
rect 31726 14306 31778 14318
rect 31726 14242 31778 14254
rect 34302 14306 34354 14318
rect 34302 14242 34354 14254
rect 35086 14306 35138 14318
rect 35086 14242 35138 14254
rect 36654 14306 36706 14318
rect 36654 14242 36706 14254
rect 39342 14306 39394 14318
rect 39342 14242 39394 14254
rect 40798 14306 40850 14318
rect 40798 14242 40850 14254
rect 42702 14306 42754 14318
rect 42702 14242 42754 14254
rect 44494 14306 44546 14318
rect 44494 14242 44546 14254
rect 45838 14306 45890 14318
rect 45838 14242 45890 14254
rect 46286 14306 46338 14318
rect 46286 14242 46338 14254
rect 46734 14306 46786 14318
rect 46734 14242 46786 14254
rect 47630 14306 47682 14318
rect 47630 14242 47682 14254
rect 49534 14306 49586 14318
rect 49534 14242 49586 14254
rect 49646 14306 49698 14318
rect 49646 14242 49698 14254
rect 50654 14306 50706 14318
rect 50654 14242 50706 14254
rect 53566 14306 53618 14318
rect 53566 14242 53618 14254
rect 54350 14306 54402 14318
rect 54350 14242 54402 14254
rect 1344 14138 58576 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 58576 14138
rect 1344 14052 58576 14086
rect 1822 13970 1874 13982
rect 1822 13906 1874 13918
rect 2270 13970 2322 13982
rect 2270 13906 2322 13918
rect 2718 13970 2770 13982
rect 2718 13906 2770 13918
rect 3166 13970 3218 13982
rect 3166 13906 3218 13918
rect 3614 13970 3666 13982
rect 3614 13906 3666 13918
rect 4510 13970 4562 13982
rect 4510 13906 4562 13918
rect 6750 13970 6802 13982
rect 6750 13906 6802 13918
rect 14702 13970 14754 13982
rect 14702 13906 14754 13918
rect 16494 13970 16546 13982
rect 16494 13906 16546 13918
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 18174 13970 18226 13982
rect 18174 13906 18226 13918
rect 19518 13970 19570 13982
rect 22654 13970 22706 13982
rect 24782 13970 24834 13982
rect 21186 13918 21198 13970
rect 21250 13918 21262 13970
rect 24210 13918 24222 13970
rect 24274 13918 24286 13970
rect 19518 13906 19570 13918
rect 22654 13906 22706 13918
rect 24782 13906 24834 13918
rect 30158 13970 30210 13982
rect 30158 13906 30210 13918
rect 30942 13970 30994 13982
rect 30942 13906 30994 13918
rect 33630 13970 33682 13982
rect 33630 13906 33682 13918
rect 34414 13970 34466 13982
rect 34414 13906 34466 13918
rect 35758 13970 35810 13982
rect 35758 13906 35810 13918
rect 37662 13970 37714 13982
rect 37662 13906 37714 13918
rect 38222 13970 38274 13982
rect 38222 13906 38274 13918
rect 40126 13970 40178 13982
rect 40126 13906 40178 13918
rect 40350 13970 40402 13982
rect 40350 13906 40402 13918
rect 43038 13970 43090 13982
rect 43038 13906 43090 13918
rect 43486 13970 43538 13982
rect 43486 13906 43538 13918
rect 44270 13970 44322 13982
rect 44270 13906 44322 13918
rect 46510 13970 46562 13982
rect 46510 13906 46562 13918
rect 47070 13970 47122 13982
rect 47070 13906 47122 13918
rect 47854 13970 47906 13982
rect 47854 13906 47906 13918
rect 48414 13970 48466 13982
rect 48414 13906 48466 13918
rect 51326 13970 51378 13982
rect 51326 13906 51378 13918
rect 57486 13970 57538 13982
rect 57486 13906 57538 13918
rect 6190 13858 6242 13870
rect 5842 13806 5854 13858
rect 5906 13806 5918 13858
rect 6190 13794 6242 13806
rect 7870 13858 7922 13870
rect 9774 13858 9826 13870
rect 8866 13806 8878 13858
rect 8930 13806 8942 13858
rect 7870 13794 7922 13806
rect 9774 13794 9826 13806
rect 18734 13858 18786 13870
rect 41806 13858 41858 13870
rect 53230 13858 53282 13870
rect 23426 13806 23438 13858
rect 23490 13806 23502 13858
rect 25890 13806 25902 13858
rect 25954 13806 25966 13858
rect 33954 13806 33966 13858
rect 34018 13806 34030 13858
rect 37538 13806 37550 13858
rect 37602 13806 37614 13858
rect 45378 13806 45390 13858
rect 45442 13806 45454 13858
rect 18734 13794 18786 13806
rect 7758 13746 7810 13758
rect 7758 13682 7810 13694
rect 8094 13746 8146 13758
rect 8094 13682 8146 13694
rect 8542 13746 8594 13758
rect 15262 13746 15314 13758
rect 16382 13746 16434 13758
rect 11218 13694 11230 13746
rect 11282 13694 11294 13746
rect 12114 13694 12126 13746
rect 12178 13694 12190 13746
rect 13458 13694 13470 13746
rect 13522 13694 13534 13746
rect 14130 13694 14142 13746
rect 14194 13694 14206 13746
rect 15810 13694 15822 13746
rect 15874 13694 15886 13746
rect 8542 13682 8594 13694
rect 15262 13682 15314 13694
rect 16382 13682 16434 13694
rect 16606 13746 16658 13758
rect 28478 13746 28530 13758
rect 21186 13694 21198 13746
rect 21250 13694 21262 13746
rect 21522 13694 21534 13746
rect 21586 13694 21598 13746
rect 23762 13694 23774 13746
rect 23826 13694 23838 13746
rect 24098 13694 24110 13746
rect 24162 13694 24174 13746
rect 27346 13694 27358 13746
rect 27410 13694 27422 13746
rect 28242 13694 28254 13746
rect 28306 13694 28318 13746
rect 16606 13682 16658 13694
rect 28478 13682 28530 13694
rect 29486 13746 29538 13758
rect 29486 13682 29538 13694
rect 30382 13746 30434 13758
rect 30382 13682 30434 13694
rect 35310 13746 35362 13758
rect 35310 13682 35362 13694
rect 36318 13746 36370 13758
rect 36530 13694 36542 13746
rect 36594 13694 36606 13746
rect 36318 13682 36370 13694
rect 4062 13634 4114 13646
rect 4062 13570 4114 13582
rect 4846 13634 4898 13646
rect 4846 13570 4898 13582
rect 5294 13634 5346 13646
rect 5294 13570 5346 13582
rect 7310 13634 7362 13646
rect 7310 13570 7362 13582
rect 17726 13634 17778 13646
rect 17726 13570 17778 13582
rect 19182 13634 19234 13646
rect 19182 13570 19234 13582
rect 20302 13634 20354 13646
rect 29934 13634 29986 13646
rect 31390 13634 31442 13646
rect 21074 13582 21086 13634
rect 21138 13582 21150 13634
rect 25554 13582 25566 13634
rect 25618 13631 25630 13634
rect 25778 13631 25790 13634
rect 25618 13585 25790 13631
rect 25618 13582 25630 13585
rect 25778 13582 25790 13585
rect 25842 13582 25854 13634
rect 30258 13582 30270 13634
rect 30322 13582 30334 13634
rect 20302 13570 20354 13582
rect 29934 13570 29986 13582
rect 31390 13570 31442 13582
rect 37214 13634 37266 13646
rect 37214 13570 37266 13582
rect 15486 13522 15538 13534
rect 29710 13522 29762 13534
rect 37553 13522 37599 13806
rect 41806 13794 41858 13806
rect 53230 13794 53282 13806
rect 38670 13746 38722 13758
rect 38670 13682 38722 13694
rect 38894 13746 38946 13758
rect 38894 13682 38946 13694
rect 39342 13746 39394 13758
rect 48750 13746 48802 13758
rect 50542 13746 50594 13758
rect 52782 13746 52834 13758
rect 42018 13694 42030 13746
rect 42082 13694 42094 13746
rect 45602 13694 45614 13746
rect 45666 13694 45678 13746
rect 47618 13694 47630 13746
rect 47682 13694 47694 13746
rect 49970 13694 49982 13746
rect 50034 13694 50046 13746
rect 52322 13694 52334 13746
rect 52386 13694 52398 13746
rect 39342 13682 39394 13694
rect 48750 13682 48802 13694
rect 50542 13682 50594 13694
rect 52782 13682 52834 13694
rect 54462 13746 54514 13758
rect 57822 13746 57874 13758
rect 54898 13694 54910 13746
rect 54962 13694 54974 13746
rect 55682 13694 55694 13746
rect 55746 13694 55758 13746
rect 54462 13682 54514 13694
rect 57822 13682 57874 13694
rect 38782 13634 38834 13646
rect 38782 13570 38834 13582
rect 40238 13634 40290 13646
rect 40238 13570 40290 13582
rect 40574 13634 40626 13646
rect 40574 13570 40626 13582
rect 42702 13634 42754 13646
rect 42702 13570 42754 13582
rect 44718 13634 44770 13646
rect 51662 13634 51714 13646
rect 49634 13582 49646 13634
rect 49698 13582 49710 13634
rect 44718 13570 44770 13582
rect 51662 13570 51714 13582
rect 54238 13634 54290 13646
rect 56018 13582 56030 13634
rect 56082 13582 56094 13634
rect 54238 13570 54290 13582
rect 40798 13522 40850 13534
rect 2258 13470 2270 13522
rect 2322 13519 2334 13522
rect 3042 13519 3054 13522
rect 2322 13473 3054 13519
rect 2322 13470 2334 13473
rect 3042 13470 3054 13473
rect 3106 13470 3118 13522
rect 10322 13470 10334 13522
rect 10386 13470 10398 13522
rect 26338 13470 26350 13522
rect 26402 13470 26414 13522
rect 28242 13470 28254 13522
rect 28306 13470 28318 13522
rect 37538 13470 37550 13522
rect 37602 13470 37614 13522
rect 53890 13470 53902 13522
rect 53954 13470 53966 13522
rect 55570 13470 55582 13522
rect 55634 13470 55646 13522
rect 15486 13458 15538 13470
rect 29710 13458 29762 13470
rect 40798 13458 40850 13470
rect 1344 13354 58576 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 58576 13354
rect 1344 13268 58576 13302
rect 16494 13186 16546 13198
rect 16494 13122 16546 13134
rect 16830 13186 16882 13198
rect 16830 13122 16882 13134
rect 22430 13186 22482 13198
rect 28366 13186 28418 13198
rect 24658 13134 24670 13186
rect 24722 13183 24734 13186
rect 24882 13183 24894 13186
rect 24722 13137 24894 13183
rect 24722 13134 24734 13137
rect 24882 13134 24894 13137
rect 24946 13134 24958 13186
rect 27346 13134 27358 13186
rect 27410 13183 27422 13186
rect 28130 13183 28142 13186
rect 27410 13137 28142 13183
rect 27410 13134 27422 13137
rect 28130 13134 28142 13137
rect 28194 13134 28206 13186
rect 22430 13122 22482 13134
rect 28366 13122 28418 13134
rect 40910 13186 40962 13198
rect 55134 13186 55186 13198
rect 48290 13134 48302 13186
rect 48354 13134 48366 13186
rect 40910 13122 40962 13134
rect 55134 13122 55186 13134
rect 1934 13074 1986 13086
rect 1934 13010 1986 13022
rect 4622 13074 4674 13086
rect 4622 13010 4674 13022
rect 7758 13074 7810 13086
rect 7758 13010 7810 13022
rect 10110 13074 10162 13086
rect 10110 13010 10162 13022
rect 15038 13074 15090 13086
rect 21534 13074 21586 13086
rect 18610 13022 18622 13074
rect 18674 13022 18686 13074
rect 20178 13022 20190 13074
rect 20242 13022 20254 13074
rect 15038 13010 15090 13022
rect 21534 13010 21586 13022
rect 22318 13074 22370 13086
rect 22318 13010 22370 13022
rect 22990 13074 23042 13086
rect 22990 13010 23042 13022
rect 27358 13074 27410 13086
rect 27358 13010 27410 13022
rect 29598 13074 29650 13086
rect 29598 13010 29650 13022
rect 30382 13074 30434 13086
rect 30382 13010 30434 13022
rect 30830 13074 30882 13086
rect 30830 13010 30882 13022
rect 32846 13074 32898 13086
rect 32846 13010 32898 13022
rect 35198 13074 35250 13086
rect 35198 13010 35250 13022
rect 36318 13074 36370 13086
rect 36318 13010 36370 13022
rect 36766 13074 36818 13086
rect 36766 13010 36818 13022
rect 38558 13074 38610 13086
rect 44158 13074 44210 13086
rect 41794 13022 41806 13074
rect 41858 13022 41870 13074
rect 38558 13010 38610 13022
rect 44158 13010 44210 13022
rect 44606 13074 44658 13086
rect 44606 13010 44658 13022
rect 45502 13074 45554 13086
rect 45502 13010 45554 13022
rect 48974 13074 49026 13086
rect 48974 13010 49026 13022
rect 49534 13074 49586 13086
rect 49534 13010 49586 13022
rect 53342 13074 53394 13086
rect 53342 13010 53394 13022
rect 55694 13074 55746 13086
rect 55694 13010 55746 13022
rect 56142 13074 56194 13086
rect 56142 13010 56194 13022
rect 57822 13074 57874 13086
rect 57822 13010 57874 13022
rect 2382 12962 2434 12974
rect 16046 12962 16098 12974
rect 6066 12910 6078 12962
rect 6130 12910 6142 12962
rect 7186 12910 7198 12962
rect 7250 12910 7262 12962
rect 9090 12910 9102 12962
rect 9154 12910 9166 12962
rect 11554 12910 11566 12962
rect 11618 12910 11630 12962
rect 12898 12910 12910 12962
rect 12962 12910 12974 12962
rect 2382 12898 2434 12910
rect 16046 12898 16098 12910
rect 16606 12962 16658 12974
rect 16606 12898 16658 12910
rect 16942 12962 16994 12974
rect 16942 12898 16994 12910
rect 17950 12962 18002 12974
rect 17950 12898 18002 12910
rect 18734 12962 18786 12974
rect 18734 12898 18786 12910
rect 19070 12962 19122 12974
rect 31278 12962 31330 12974
rect 19730 12910 19742 12962
rect 19794 12910 19806 12962
rect 20850 12910 20862 12962
rect 20914 12910 20926 12962
rect 22082 12910 22094 12962
rect 22146 12910 22158 12962
rect 25330 12910 25342 12962
rect 25394 12910 25406 12962
rect 26450 12910 26462 12962
rect 26514 12910 26526 12962
rect 19070 12898 19122 12910
rect 31278 12898 31330 12910
rect 33294 12962 33346 12974
rect 33294 12898 33346 12910
rect 33630 12962 33682 12974
rect 39118 12962 39170 12974
rect 37762 12910 37774 12962
rect 37826 12910 37838 12962
rect 33630 12898 33682 12910
rect 39118 12898 39170 12910
rect 39902 12962 39954 12974
rect 39902 12898 39954 12910
rect 40238 12962 40290 12974
rect 40238 12898 40290 12910
rect 41022 12962 41074 12974
rect 46398 12962 46450 12974
rect 42018 12910 42030 12962
rect 42082 12910 42094 12962
rect 46162 12910 46174 12962
rect 46226 12910 46238 12962
rect 41022 12898 41074 12910
rect 46398 12898 46450 12910
rect 47742 12962 47794 12974
rect 47742 12898 47794 12910
rect 47966 12962 48018 12974
rect 47966 12898 48018 12910
rect 49198 12962 49250 12974
rect 49198 12898 49250 12910
rect 51774 12962 51826 12974
rect 51774 12898 51826 12910
rect 14254 12850 14306 12862
rect 3602 12798 3614 12850
rect 3666 12798 3678 12850
rect 8754 12798 8766 12850
rect 8818 12798 8830 12850
rect 10882 12798 10894 12850
rect 10946 12798 10958 12850
rect 12786 12798 12798 12850
rect 12850 12798 12862 12850
rect 14254 12786 14306 12798
rect 14590 12850 14642 12862
rect 14590 12786 14642 12798
rect 17614 12850 17666 12862
rect 23662 12850 23714 12862
rect 20738 12798 20750 12850
rect 20802 12798 20814 12850
rect 17614 12786 17666 12798
rect 23662 12786 23714 12798
rect 23998 12850 24050 12862
rect 28478 12850 28530 12862
rect 25554 12798 25566 12850
rect 25618 12798 25630 12850
rect 23998 12786 24050 12798
rect 28478 12786 28530 12798
rect 33966 12850 34018 12862
rect 33966 12786 34018 12798
rect 34526 12850 34578 12862
rect 34526 12786 34578 12798
rect 34638 12850 34690 12862
rect 34638 12786 34690 12798
rect 39454 12850 39506 12862
rect 39454 12786 39506 12798
rect 40910 12850 40962 12862
rect 40910 12786 40962 12798
rect 42590 12850 42642 12862
rect 42590 12786 42642 12798
rect 43262 12850 43314 12862
rect 43262 12786 43314 12798
rect 49646 12850 49698 12862
rect 52334 12850 52386 12862
rect 51426 12798 51438 12850
rect 51490 12798 51502 12850
rect 49646 12786 49698 12798
rect 52334 12786 52386 12798
rect 52670 12850 52722 12862
rect 52670 12786 52722 12798
rect 54126 12850 54178 12862
rect 54126 12786 54178 12798
rect 54462 12850 54514 12862
rect 54462 12786 54514 12798
rect 55134 12850 55186 12862
rect 55134 12786 55186 12798
rect 55246 12850 55298 12862
rect 55246 12786 55298 12798
rect 57038 12850 57090 12862
rect 57038 12786 57090 12798
rect 57374 12850 57426 12862
rect 57374 12786 57426 12798
rect 2718 12738 2770 12750
rect 2718 12674 2770 12686
rect 3950 12738 4002 12750
rect 3950 12674 4002 12686
rect 5070 12738 5122 12750
rect 5070 12674 5122 12686
rect 13806 12738 13858 12750
rect 13806 12674 13858 12686
rect 15598 12738 15650 12750
rect 15598 12674 15650 12686
rect 18622 12738 18674 12750
rect 18622 12674 18674 12686
rect 18958 12738 19010 12750
rect 18958 12674 19010 12686
rect 24670 12738 24722 12750
rect 24670 12674 24722 12686
rect 26686 12738 26738 12750
rect 26686 12674 26738 12686
rect 27806 12738 27858 12750
rect 27806 12674 27858 12686
rect 29934 12738 29986 12750
rect 29934 12674 29986 12686
rect 33630 12738 33682 12750
rect 33630 12674 33682 12686
rect 34862 12738 34914 12750
rect 34862 12674 34914 12686
rect 35646 12738 35698 12750
rect 35646 12674 35698 12686
rect 37998 12738 38050 12750
rect 37998 12674 38050 12686
rect 40126 12738 40178 12750
rect 40126 12674 40178 12686
rect 43598 12738 43650 12750
rect 43598 12674 43650 12686
rect 47070 12738 47122 12750
rect 47070 12674 47122 12686
rect 49422 12738 49474 12750
rect 49422 12674 49474 12686
rect 50318 12738 50370 12750
rect 50642 12686 50654 12738
rect 50706 12686 50718 12738
rect 50318 12674 50370 12686
rect 1344 12570 58576 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 58576 12570
rect 1344 12484 58576 12518
rect 4398 12402 4450 12414
rect 6190 12402 6242 12414
rect 6066 12350 6078 12402
rect 6130 12350 6142 12402
rect 4398 12338 4450 12350
rect 6190 12338 6242 12350
rect 8654 12402 8706 12414
rect 8654 12338 8706 12350
rect 11678 12402 11730 12414
rect 11678 12338 11730 12350
rect 12238 12402 12290 12414
rect 13134 12402 13186 12414
rect 15150 12402 15202 12414
rect 12562 12350 12574 12402
rect 12626 12350 12638 12402
rect 14018 12350 14030 12402
rect 14082 12350 14094 12402
rect 12238 12338 12290 12350
rect 13134 12338 13186 12350
rect 15150 12338 15202 12350
rect 15710 12402 15762 12414
rect 15710 12338 15762 12350
rect 16046 12402 16098 12414
rect 17950 12402 18002 12414
rect 16594 12350 16606 12402
rect 16658 12350 16670 12402
rect 16046 12338 16098 12350
rect 17950 12338 18002 12350
rect 18734 12402 18786 12414
rect 18734 12338 18786 12350
rect 19854 12402 19906 12414
rect 21422 12402 21474 12414
rect 23662 12402 23714 12414
rect 20626 12350 20638 12402
rect 20690 12350 20702 12402
rect 22866 12350 22878 12402
rect 22930 12350 22942 12402
rect 19854 12338 19906 12350
rect 21422 12338 21474 12350
rect 23662 12338 23714 12350
rect 24222 12402 24274 12414
rect 25566 12402 25618 12414
rect 24546 12350 24558 12402
rect 24610 12350 24622 12402
rect 24222 12338 24274 12350
rect 25566 12338 25618 12350
rect 27582 12402 27634 12414
rect 27582 12338 27634 12350
rect 28590 12402 28642 12414
rect 37550 12402 37602 12414
rect 29810 12350 29822 12402
rect 29874 12350 29886 12402
rect 28590 12338 28642 12350
rect 37550 12338 37602 12350
rect 38334 12402 38386 12414
rect 38334 12338 38386 12350
rect 38670 12402 38722 12414
rect 38670 12338 38722 12350
rect 39230 12402 39282 12414
rect 39230 12338 39282 12350
rect 40014 12402 40066 12414
rect 40014 12338 40066 12350
rect 40574 12402 40626 12414
rect 40574 12338 40626 12350
rect 41470 12402 41522 12414
rect 41470 12338 41522 12350
rect 42254 12402 42306 12414
rect 42254 12338 42306 12350
rect 43374 12402 43426 12414
rect 45726 12402 45778 12414
rect 44818 12350 44830 12402
rect 44882 12350 44894 12402
rect 43374 12338 43426 12350
rect 45726 12338 45778 12350
rect 46174 12402 46226 12414
rect 46174 12338 46226 12350
rect 46734 12402 46786 12414
rect 46734 12338 46786 12350
rect 47294 12402 47346 12414
rect 47294 12338 47346 12350
rect 48750 12402 48802 12414
rect 48750 12338 48802 12350
rect 50878 12402 50930 12414
rect 50878 12338 50930 12350
rect 51662 12402 51714 12414
rect 51662 12338 51714 12350
rect 52558 12402 52610 12414
rect 52558 12338 52610 12350
rect 53118 12402 53170 12414
rect 56590 12402 56642 12414
rect 56018 12350 56030 12402
rect 56082 12350 56094 12402
rect 53118 12338 53170 12350
rect 56590 12338 56642 12350
rect 57374 12402 57426 12414
rect 57374 12338 57426 12350
rect 57822 12402 57874 12414
rect 57822 12338 57874 12350
rect 4062 12290 4114 12302
rect 9662 12290 9714 12302
rect 18958 12290 19010 12302
rect 5058 12238 5070 12290
rect 5122 12238 5134 12290
rect 8082 12238 8094 12290
rect 8146 12238 8158 12290
rect 11106 12238 11118 12290
rect 11170 12238 11182 12290
rect 13458 12238 13470 12290
rect 13522 12238 13534 12290
rect 4062 12226 4114 12238
rect 9662 12226 9714 12238
rect 18958 12226 19010 12238
rect 19518 12290 19570 12302
rect 19518 12226 19570 12238
rect 21870 12290 21922 12302
rect 21870 12226 21922 12238
rect 22094 12290 22146 12302
rect 22094 12226 22146 12238
rect 22206 12290 22258 12302
rect 22206 12226 22258 12238
rect 26462 12290 26514 12302
rect 26462 12226 26514 12238
rect 27470 12290 27522 12302
rect 27470 12226 27522 12238
rect 31166 12290 31218 12302
rect 42702 12290 42754 12302
rect 33954 12238 33966 12290
rect 34018 12238 34030 12290
rect 34402 12238 34414 12290
rect 34466 12238 34478 12290
rect 36306 12238 36318 12290
rect 36370 12238 36382 12290
rect 36866 12238 36878 12290
rect 36930 12238 36942 12290
rect 31166 12226 31218 12238
rect 42702 12226 42754 12238
rect 48638 12290 48690 12302
rect 48638 12226 48690 12238
rect 49870 12290 49922 12302
rect 49870 12226 49922 12238
rect 55134 12290 55186 12302
rect 55134 12226 55186 12238
rect 8990 12178 9042 12190
rect 14366 12178 14418 12190
rect 19854 12178 19906 12190
rect 2818 12126 2830 12178
rect 2882 12126 2894 12178
rect 5170 12126 5182 12178
rect 5234 12126 5246 12178
rect 5842 12126 5854 12178
rect 5906 12126 5918 12178
rect 6962 12126 6974 12178
rect 7026 12126 7038 12178
rect 7634 12126 7646 12178
rect 7698 12126 7710 12178
rect 9874 12126 9886 12178
rect 9938 12126 9950 12178
rect 10434 12126 10446 12178
rect 10498 12126 10510 12178
rect 10994 12126 11006 12178
rect 11058 12126 11070 12178
rect 16818 12126 16830 12178
rect 16882 12126 16894 12178
rect 18498 12126 18510 12178
rect 18562 12126 18574 12178
rect 8990 12114 9042 12126
rect 14366 12114 14418 12126
rect 19854 12114 19906 12126
rect 20078 12178 20130 12190
rect 23214 12178 23266 12190
rect 20850 12126 20862 12178
rect 20914 12126 20926 12178
rect 20078 12114 20130 12126
rect 23214 12114 23266 12126
rect 28926 12178 28978 12190
rect 36094 12178 36146 12190
rect 45390 12178 45442 12190
rect 52222 12178 52274 12190
rect 55694 12178 55746 12190
rect 29586 12126 29598 12178
rect 29650 12126 29662 12178
rect 44594 12126 44606 12178
rect 44658 12126 44670 12178
rect 49634 12126 49646 12178
rect 49698 12126 49710 12178
rect 53330 12126 53342 12178
rect 53394 12126 53406 12178
rect 54226 12126 54238 12178
rect 54290 12126 54302 12178
rect 28926 12114 28978 12126
rect 36094 12114 36146 12126
rect 45390 12114 45442 12126
rect 52222 12114 52274 12126
rect 55694 12114 55746 12126
rect 3614 12066 3666 12078
rect 26014 12066 26066 12078
rect 1922 12014 1934 12066
rect 1986 12014 1998 12066
rect 7970 12014 7982 12066
rect 8034 12014 8046 12066
rect 18834 12014 18846 12066
rect 18898 12014 18910 12066
rect 3614 12002 3666 12014
rect 26014 12002 26066 12014
rect 30270 12066 30322 12078
rect 30270 12002 30322 12014
rect 30718 12066 30770 12078
rect 30718 12002 30770 12014
rect 32846 12066 32898 12078
rect 32846 12002 32898 12014
rect 43710 12066 43762 12078
rect 43710 12002 43762 12014
rect 47742 12066 47794 12078
rect 47742 12002 47794 12014
rect 50318 12066 50370 12078
rect 50318 12002 50370 12014
rect 51214 12066 51266 12078
rect 54338 12014 54350 12066
rect 54402 12014 54414 12066
rect 51214 12002 51266 12014
rect 27694 11954 27746 11966
rect 25442 11902 25454 11954
rect 25506 11951 25518 11954
rect 26002 11951 26014 11954
rect 25506 11905 26014 11951
rect 25506 11902 25518 11905
rect 26002 11902 26014 11905
rect 26066 11902 26078 11954
rect 27694 11890 27746 11902
rect 34638 11954 34690 11966
rect 34638 11890 34690 11902
rect 34974 11954 35026 11966
rect 34974 11890 35026 11902
rect 35758 11954 35810 11966
rect 35758 11890 35810 11902
rect 1344 11786 58576 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 58576 11786
rect 1344 11700 58576 11734
rect 11230 11618 11282 11630
rect 33854 11618 33906 11630
rect 16930 11566 16942 11618
rect 16994 11566 17006 11618
rect 26114 11566 26126 11618
rect 26178 11566 26190 11618
rect 11230 11554 11282 11566
rect 33854 11554 33906 11566
rect 41806 11618 41858 11630
rect 46274 11566 46286 11618
rect 46338 11615 46350 11618
rect 46834 11615 46846 11618
rect 46338 11569 46846 11615
rect 46338 11566 46350 11569
rect 46834 11566 46846 11569
rect 46898 11566 46910 11618
rect 55682 11566 55694 11618
rect 55746 11615 55758 11618
rect 56354 11615 56366 11618
rect 55746 11569 56366 11615
rect 55746 11566 55758 11569
rect 56354 11566 56366 11569
rect 56418 11566 56430 11618
rect 57250 11566 57262 11618
rect 57314 11615 57326 11618
rect 57314 11569 57983 11615
rect 57314 11566 57326 11569
rect 41806 11554 41858 11566
rect 4846 11506 4898 11518
rect 15934 11506 15986 11518
rect 21646 11506 21698 11518
rect 6962 11454 6974 11506
rect 7026 11454 7038 11506
rect 8306 11454 8318 11506
rect 8370 11454 8382 11506
rect 13794 11454 13806 11506
rect 13858 11454 13870 11506
rect 14242 11454 14254 11506
rect 14306 11454 14318 11506
rect 17266 11454 17278 11506
rect 17330 11454 17342 11506
rect 4846 11442 4898 11454
rect 15934 11442 15986 11454
rect 21646 11442 21698 11454
rect 28030 11506 28082 11518
rect 30494 11506 30546 11518
rect 35758 11506 35810 11518
rect 28578 11454 28590 11506
rect 28642 11454 28654 11506
rect 34066 11454 34078 11506
rect 34130 11454 34142 11506
rect 28030 11442 28082 11454
rect 30494 11442 30546 11454
rect 35758 11442 35810 11454
rect 36878 11506 36930 11518
rect 36878 11442 36930 11454
rect 37774 11506 37826 11518
rect 37774 11442 37826 11454
rect 42254 11506 42306 11518
rect 42254 11442 42306 11454
rect 43038 11506 43090 11518
rect 43038 11442 43090 11454
rect 43486 11506 43538 11518
rect 43486 11442 43538 11454
rect 44046 11506 44098 11518
rect 44046 11442 44098 11454
rect 46286 11506 46338 11518
rect 46286 11442 46338 11454
rect 46622 11506 46674 11518
rect 46622 11442 46674 11454
rect 47070 11506 47122 11518
rect 47070 11442 47122 11454
rect 47630 11506 47682 11518
rect 47630 11442 47682 11454
rect 47966 11506 48018 11518
rect 47966 11442 48018 11454
rect 49422 11506 49474 11518
rect 49422 11442 49474 11454
rect 49870 11506 49922 11518
rect 49870 11442 49922 11454
rect 52110 11506 52162 11518
rect 52110 11442 52162 11454
rect 55358 11506 55410 11518
rect 55358 11442 55410 11454
rect 55806 11506 55858 11518
rect 55806 11442 55858 11454
rect 56254 11506 56306 11518
rect 56254 11442 56306 11454
rect 57150 11506 57202 11518
rect 57150 11442 57202 11454
rect 57598 11506 57650 11518
rect 57937 11506 57983 11569
rect 58034 11566 58046 11618
rect 58098 11615 58110 11618
rect 58258 11615 58270 11618
rect 58098 11569 58270 11615
rect 58098 11566 58110 11569
rect 58258 11566 58270 11569
rect 58322 11566 58334 11618
rect 58046 11506 58098 11518
rect 57922 11454 57934 11506
rect 57986 11454 57998 11506
rect 57598 11442 57650 11454
rect 58046 11442 58098 11454
rect 4958 11394 5010 11406
rect 23214 11394 23266 11406
rect 25790 11394 25842 11406
rect 7410 11342 7422 11394
rect 7474 11342 7486 11394
rect 8866 11342 8878 11394
rect 8930 11342 8942 11394
rect 10434 11342 10446 11394
rect 10498 11342 10510 11394
rect 10658 11342 10670 11394
rect 10722 11342 10734 11394
rect 13570 11342 13582 11394
rect 13634 11342 13646 11394
rect 14690 11342 14702 11394
rect 14754 11342 14766 11394
rect 17490 11342 17502 11394
rect 17554 11342 17566 11394
rect 18946 11342 18958 11394
rect 19010 11342 19022 11394
rect 19170 11342 19182 11394
rect 19234 11342 19246 11394
rect 19618 11342 19630 11394
rect 19682 11342 19694 11394
rect 24882 11342 24894 11394
rect 24946 11342 24958 11394
rect 4958 11330 5010 11342
rect 23214 11330 23266 11342
rect 25790 11330 25842 11342
rect 27246 11394 27298 11406
rect 27246 11330 27298 11342
rect 27470 11394 27522 11406
rect 27470 11330 27522 11342
rect 28366 11394 28418 11406
rect 28366 11330 28418 11342
rect 38110 11394 38162 11406
rect 51326 11394 51378 11406
rect 56702 11394 56754 11406
rect 38658 11342 38670 11394
rect 38722 11342 38734 11394
rect 54338 11342 54350 11394
rect 54402 11342 54414 11394
rect 38110 11330 38162 11342
rect 51326 11330 51378 11342
rect 56702 11330 56754 11342
rect 1822 11282 1874 11294
rect 1822 11218 1874 11230
rect 2270 11282 2322 11294
rect 2270 11218 2322 11230
rect 2606 11282 2658 11294
rect 2606 11218 2658 11230
rect 11790 11282 11842 11294
rect 11790 11218 11842 11230
rect 12350 11282 12402 11294
rect 12350 11218 12402 11230
rect 22654 11282 22706 11294
rect 22654 11218 22706 11230
rect 22878 11282 22930 11294
rect 25566 11282 25618 11294
rect 24098 11230 24110 11282
rect 24162 11230 24174 11282
rect 24658 11230 24670 11282
rect 24722 11230 24734 11282
rect 22878 11218 22930 11230
rect 25566 11218 25618 11230
rect 29598 11282 29650 11294
rect 29598 11218 29650 11230
rect 29934 11282 29986 11294
rect 29934 11218 29986 11230
rect 48526 11282 48578 11294
rect 48526 11218 48578 11230
rect 48862 11282 48914 11294
rect 48862 11218 48914 11230
rect 51662 11282 51714 11294
rect 51662 11218 51714 11230
rect 52782 11282 52834 11294
rect 52782 11218 52834 11230
rect 53342 11282 53394 11294
rect 53342 11218 53394 11230
rect 54126 11282 54178 11294
rect 54126 11218 54178 11230
rect 3166 11170 3218 11182
rect 4510 11170 4562 11182
rect 3490 11118 3502 11170
rect 3554 11118 3566 11170
rect 3166 11106 3218 11118
rect 4510 11106 4562 11118
rect 4734 11170 4786 11182
rect 4734 11106 4786 11118
rect 5742 11170 5794 11182
rect 5742 11106 5794 11118
rect 11342 11170 11394 11182
rect 11342 11106 11394 11118
rect 11566 11170 11618 11182
rect 11566 11106 11618 11118
rect 12686 11170 12738 11182
rect 12686 11106 12738 11118
rect 22094 11170 22146 11182
rect 22094 11106 22146 11118
rect 23102 11170 23154 11182
rect 23102 11106 23154 11118
rect 23774 11170 23826 11182
rect 30830 11170 30882 11182
rect 26898 11118 26910 11170
rect 26962 11118 26974 11170
rect 23774 11106 23826 11118
rect 30830 11106 30882 11118
rect 34078 11170 34130 11182
rect 34078 11106 34130 11118
rect 34638 11170 34690 11182
rect 34638 11106 34690 11118
rect 35310 11170 35362 11182
rect 35310 11106 35362 11118
rect 36318 11170 36370 11182
rect 42590 11170 42642 11182
rect 41010 11118 41022 11170
rect 41074 11118 41086 11170
rect 36318 11106 36370 11118
rect 42590 11106 42642 11118
rect 44718 11170 44770 11182
rect 44718 11106 44770 11118
rect 45502 11170 45554 11182
rect 45502 11106 45554 11118
rect 50206 11170 50258 11182
rect 50206 11106 50258 11118
rect 50654 11170 50706 11182
rect 50654 11106 50706 11118
rect 54910 11170 54962 11182
rect 54910 11106 54962 11118
rect 1344 11002 58576 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 58576 11002
rect 1344 10916 58576 10950
rect 2830 10834 2882 10846
rect 2830 10770 2882 10782
rect 3838 10834 3890 10846
rect 3838 10770 3890 10782
rect 4286 10834 4338 10846
rect 4286 10770 4338 10782
rect 4622 10834 4674 10846
rect 12014 10834 12066 10846
rect 6738 10782 6750 10834
rect 6802 10782 6814 10834
rect 4622 10770 4674 10782
rect 12014 10770 12066 10782
rect 12798 10834 12850 10846
rect 12798 10770 12850 10782
rect 14702 10834 14754 10846
rect 14702 10770 14754 10782
rect 15262 10834 15314 10846
rect 15262 10770 15314 10782
rect 17950 10834 18002 10846
rect 24222 10834 24274 10846
rect 18274 10782 18286 10834
rect 18338 10782 18350 10834
rect 17950 10770 18002 10782
rect 24222 10770 24274 10782
rect 25790 10834 25842 10846
rect 29822 10834 29874 10846
rect 26114 10782 26126 10834
rect 26178 10782 26190 10834
rect 27010 10782 27022 10834
rect 27074 10782 27086 10834
rect 25790 10770 25842 10782
rect 29822 10770 29874 10782
rect 37326 10834 37378 10846
rect 37326 10770 37378 10782
rect 38670 10834 38722 10846
rect 38670 10770 38722 10782
rect 39118 10834 39170 10846
rect 39118 10770 39170 10782
rect 40126 10834 40178 10846
rect 40126 10770 40178 10782
rect 40574 10834 40626 10846
rect 40574 10770 40626 10782
rect 41582 10834 41634 10846
rect 41582 10770 41634 10782
rect 42590 10834 42642 10846
rect 42590 10770 42642 10782
rect 43150 10834 43202 10846
rect 49422 10834 49474 10846
rect 47954 10782 47966 10834
rect 48018 10782 48030 10834
rect 43150 10770 43202 10782
rect 49422 10770 49474 10782
rect 49870 10834 49922 10846
rect 49870 10770 49922 10782
rect 50766 10834 50818 10846
rect 50766 10770 50818 10782
rect 51774 10834 51826 10846
rect 51774 10770 51826 10782
rect 52670 10834 52722 10846
rect 52670 10770 52722 10782
rect 53566 10834 53618 10846
rect 53566 10770 53618 10782
rect 53902 10834 53954 10846
rect 53902 10770 53954 10782
rect 54350 10834 54402 10846
rect 54350 10770 54402 10782
rect 54798 10834 54850 10846
rect 54798 10770 54850 10782
rect 55358 10834 55410 10846
rect 55358 10770 55410 10782
rect 55694 10834 55746 10846
rect 55694 10770 55746 10782
rect 57374 10834 57426 10846
rect 57374 10770 57426 10782
rect 57934 10834 57986 10846
rect 57934 10770 57986 10782
rect 2158 10722 2210 10734
rect 2158 10658 2210 10670
rect 2270 10722 2322 10734
rect 8878 10722 8930 10734
rect 3154 10670 3166 10722
rect 3218 10670 3230 10722
rect 5170 10670 5182 10722
rect 5234 10670 5246 10722
rect 6290 10670 6302 10722
rect 6354 10670 6366 10722
rect 7858 10670 7870 10722
rect 7922 10670 7934 10722
rect 8306 10670 8318 10722
rect 8370 10670 8382 10722
rect 2270 10658 2322 10670
rect 8878 10658 8930 10670
rect 14590 10722 14642 10734
rect 14590 10658 14642 10670
rect 14814 10722 14866 10734
rect 27582 10722 27634 10734
rect 15810 10670 15822 10722
rect 15874 10670 15886 10722
rect 18834 10670 18846 10722
rect 18898 10670 18910 10722
rect 20402 10670 20414 10722
rect 20466 10670 20478 10722
rect 22194 10670 22206 10722
rect 22258 10670 22270 10722
rect 14814 10658 14866 10670
rect 27582 10658 27634 10670
rect 28478 10722 28530 10734
rect 28478 10658 28530 10670
rect 30158 10722 30210 10734
rect 30158 10658 30210 10670
rect 34974 10722 35026 10734
rect 34974 10658 35026 10670
rect 36094 10722 36146 10734
rect 36094 10658 36146 10670
rect 5518 10610 5570 10622
rect 12350 10610 12402 10622
rect 6402 10558 6414 10610
rect 6466 10558 6478 10610
rect 7746 10558 7758 10610
rect 7810 10558 7822 10610
rect 10098 10558 10110 10610
rect 10162 10558 10174 10610
rect 10770 10558 10782 10610
rect 10834 10558 10846 10610
rect 11330 10558 11342 10610
rect 11394 10558 11406 10610
rect 5518 10546 5570 10558
rect 12350 10546 12402 10558
rect 13358 10610 13410 10622
rect 19182 10610 19234 10622
rect 23886 10610 23938 10622
rect 16034 10558 16046 10610
rect 16098 10558 16110 10610
rect 16930 10558 16942 10610
rect 16994 10558 17006 10610
rect 19954 10558 19966 10610
rect 20018 10558 20030 10610
rect 20290 10558 20302 10610
rect 20354 10558 20366 10610
rect 22082 10558 22094 10610
rect 22146 10558 22158 10610
rect 23090 10558 23102 10610
rect 23154 10558 23166 10610
rect 13358 10546 13410 10558
rect 19182 10546 19234 10558
rect 23886 10546 23938 10558
rect 23998 10610 24050 10622
rect 23998 10546 24050 10558
rect 24334 10610 24386 10622
rect 24334 10546 24386 10558
rect 27358 10610 27410 10622
rect 27358 10546 27410 10558
rect 28142 10610 28194 10622
rect 45054 10610 45106 10622
rect 51214 10610 51266 10622
rect 34738 10558 34750 10610
rect 34802 10558 34814 10610
rect 35858 10558 35870 10610
rect 35922 10558 35934 10610
rect 45378 10558 45390 10610
rect 45442 10558 45454 10610
rect 28142 10546 28194 10558
rect 45054 10546 45106 10558
rect 51214 10546 51266 10558
rect 13918 10498 13970 10510
rect 21534 10498 21586 10510
rect 24782 10498 24834 10510
rect 10434 10446 10446 10498
rect 10498 10446 10510 10498
rect 16258 10446 16270 10498
rect 16322 10446 16334 10498
rect 20178 10446 20190 10498
rect 20242 10446 20254 10498
rect 22530 10446 22542 10498
rect 22594 10446 22606 10498
rect 13918 10434 13970 10446
rect 21534 10434 21586 10446
rect 24782 10434 24834 10446
rect 29262 10498 29314 10510
rect 29262 10434 29314 10446
rect 37662 10498 37714 10510
rect 37662 10434 37714 10446
rect 38222 10498 38274 10510
rect 38222 10434 38274 10446
rect 39454 10498 39506 10510
rect 39454 10434 39506 10446
rect 41918 10498 41970 10510
rect 41918 10434 41970 10446
rect 43598 10498 43650 10510
rect 43598 10434 43650 10446
rect 44046 10498 44098 10510
rect 44046 10434 44098 10446
rect 44382 10498 44434 10510
rect 44382 10434 44434 10446
rect 50430 10498 50482 10510
rect 50430 10434 50482 10446
rect 52110 10498 52162 10510
rect 52110 10434 52162 10446
rect 53006 10498 53058 10510
rect 53006 10434 53058 10446
rect 56478 10498 56530 10510
rect 56478 10434 56530 10446
rect 48526 10386 48578 10398
rect 43922 10334 43934 10386
rect 43986 10383 43998 10386
rect 44370 10383 44382 10386
rect 43986 10337 44382 10383
rect 43986 10334 43998 10337
rect 44370 10334 44382 10337
rect 44434 10383 44446 10386
rect 44706 10383 44718 10386
rect 44434 10337 44718 10383
rect 44434 10334 44446 10337
rect 44706 10334 44718 10337
rect 44770 10334 44782 10386
rect 50418 10334 50430 10386
rect 50482 10383 50494 10386
rect 51650 10383 51662 10386
rect 50482 10337 51662 10383
rect 50482 10334 50494 10337
rect 51650 10334 51662 10337
rect 51714 10334 51726 10386
rect 53890 10334 53902 10386
rect 53954 10383 53966 10386
rect 54450 10383 54462 10386
rect 53954 10337 54462 10383
rect 53954 10334 53966 10337
rect 54450 10334 54462 10337
rect 54514 10334 54526 10386
rect 48526 10322 48578 10334
rect 1344 10218 58576 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 58576 10218
rect 1344 10132 58576 10166
rect 25678 10050 25730 10062
rect 1922 9998 1934 10050
rect 1986 10047 1998 10050
rect 3154 10047 3166 10050
rect 1986 10001 3166 10047
rect 1986 9998 1998 10001
rect 3154 9998 3166 10001
rect 3218 9998 3230 10050
rect 5954 9998 5966 10050
rect 6018 9998 6030 10050
rect 25678 9986 25730 9998
rect 26574 10050 26626 10062
rect 26574 9986 26626 9998
rect 41694 10050 41746 10062
rect 41694 9986 41746 9998
rect 49086 10050 49138 10062
rect 49086 9986 49138 9998
rect 1934 9938 1986 9950
rect 1934 9874 1986 9886
rect 2382 9938 2434 9950
rect 2382 9874 2434 9886
rect 4062 9938 4114 9950
rect 8094 9938 8146 9950
rect 11342 9938 11394 9950
rect 6402 9886 6414 9938
rect 6466 9886 6478 9938
rect 8866 9886 8878 9938
rect 8930 9886 8942 9938
rect 9986 9886 9998 9938
rect 10050 9886 10062 9938
rect 4062 9874 4114 9886
rect 8094 9874 8146 9886
rect 11342 9874 11394 9886
rect 14142 9938 14194 9950
rect 14142 9874 14194 9886
rect 19854 9938 19906 9950
rect 28254 9938 28306 9950
rect 20402 9886 20414 9938
rect 20466 9886 20478 9938
rect 22194 9886 22206 9938
rect 22258 9886 22270 9938
rect 19854 9874 19906 9886
rect 28254 9874 28306 9886
rect 29486 9938 29538 9950
rect 29486 9874 29538 9886
rect 43038 9938 43090 9950
rect 43038 9874 43090 9886
rect 43374 9938 43426 9950
rect 43374 9874 43426 9886
rect 44382 9938 44434 9950
rect 44382 9874 44434 9886
rect 49422 9938 49474 9950
rect 49422 9874 49474 9886
rect 52446 9938 52498 9950
rect 52446 9874 52498 9886
rect 53342 9938 53394 9950
rect 53342 9874 53394 9886
rect 53790 9938 53842 9950
rect 53790 9874 53842 9886
rect 55134 9938 55186 9950
rect 55134 9874 55186 9886
rect 55582 9938 55634 9950
rect 55582 9874 55634 9886
rect 56254 9938 56306 9950
rect 56254 9874 56306 9886
rect 56702 9938 56754 9950
rect 56702 9874 56754 9886
rect 57262 9938 57314 9950
rect 57262 9874 57314 9886
rect 57598 9938 57650 9950
rect 57598 9874 57650 9886
rect 58046 9938 58098 9950
rect 58046 9874 58098 9886
rect 4958 9826 5010 9838
rect 4958 9762 5010 9774
rect 6190 9826 6242 9838
rect 6190 9762 6242 9774
rect 7086 9826 7138 9838
rect 13806 9826 13858 9838
rect 8978 9774 8990 9826
rect 9042 9774 9054 9826
rect 9650 9774 9662 9826
rect 9714 9774 9726 9826
rect 7086 9762 7138 9774
rect 13806 9762 13858 9774
rect 14366 9826 14418 9838
rect 14366 9762 14418 9774
rect 14926 9826 14978 9838
rect 15934 9826 15986 9838
rect 17502 9826 17554 9838
rect 18958 9826 19010 9838
rect 25902 9826 25954 9838
rect 15250 9774 15262 9826
rect 15314 9774 15326 9826
rect 16146 9774 16158 9826
rect 16210 9774 16222 9826
rect 17826 9774 17838 9826
rect 17890 9774 17902 9826
rect 22306 9774 22318 9826
rect 22370 9774 22382 9826
rect 22530 9774 22542 9826
rect 22594 9774 22606 9826
rect 14926 9762 14978 9774
rect 15934 9762 15986 9774
rect 17502 9762 17554 9774
rect 18958 9762 19010 9774
rect 25902 9762 25954 9774
rect 26126 9826 26178 9838
rect 26126 9762 26178 9774
rect 27022 9826 27074 9838
rect 27022 9762 27074 9774
rect 38222 9826 38274 9838
rect 38658 9774 38670 9826
rect 38722 9774 38734 9826
rect 45490 9774 45502 9826
rect 45554 9774 45566 9826
rect 45938 9774 45950 9826
rect 46002 9774 46014 9826
rect 38222 9762 38274 9774
rect 4622 9714 4674 9726
rect 4622 9650 4674 9662
rect 7310 9714 7362 9726
rect 7310 9650 7362 9662
rect 7422 9714 7474 9726
rect 7422 9650 7474 9662
rect 8542 9714 8594 9726
rect 13918 9714 13970 9726
rect 18622 9714 18674 9726
rect 25454 9714 25506 9726
rect 48302 9714 48354 9726
rect 12898 9662 12910 9714
rect 12962 9662 12974 9714
rect 15362 9662 15374 9714
rect 15426 9662 15438 9714
rect 24098 9662 24110 9714
rect 24162 9662 24174 9714
rect 27346 9662 27358 9714
rect 27410 9662 27422 9714
rect 51874 9662 51886 9714
rect 51938 9662 51950 9714
rect 8542 9650 8594 9662
rect 13918 9650 13970 9662
rect 18622 9650 18674 9662
rect 25454 9650 25506 9662
rect 48302 9650 48354 9662
rect 2830 9602 2882 9614
rect 2830 9538 2882 9550
rect 3166 9602 3218 9614
rect 3166 9538 3218 9550
rect 3726 9602 3778 9614
rect 3726 9538 3778 9550
rect 10782 9602 10834 9614
rect 10782 9538 10834 9550
rect 12014 9602 12066 9614
rect 12014 9538 12066 9550
rect 12574 9602 12626 9614
rect 12574 9538 12626 9550
rect 17950 9602 18002 9614
rect 17950 9538 18002 9550
rect 20862 9602 20914 9614
rect 23774 9602 23826 9614
rect 23202 9550 23214 9602
rect 23266 9550 23278 9602
rect 20862 9538 20914 9550
rect 23774 9538 23826 9550
rect 24558 9602 24610 9614
rect 24558 9538 24610 9550
rect 27806 9602 27858 9614
rect 27806 9538 27858 9550
rect 28702 9602 28754 9614
rect 28702 9538 28754 9550
rect 37550 9602 37602 9614
rect 42478 9602 42530 9614
rect 41010 9550 41022 9602
rect 41074 9550 41086 9602
rect 42130 9550 42142 9602
rect 42194 9550 42206 9602
rect 37550 9538 37602 9550
rect 42478 9538 42530 9550
rect 43934 9602 43986 9614
rect 43934 9538 43986 9550
rect 44718 9602 44770 9614
rect 44718 9538 44770 9550
rect 54238 9602 54290 9614
rect 54238 9538 54290 9550
rect 54686 9602 54738 9614
rect 54686 9538 54738 9550
rect 1344 9434 58576 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 58576 9434
rect 1344 9348 58576 9382
rect 3726 9266 3778 9278
rect 3726 9202 3778 9214
rect 4062 9266 4114 9278
rect 4062 9202 4114 9214
rect 5070 9266 5122 9278
rect 7198 9266 7250 9278
rect 6290 9214 6302 9266
rect 6354 9214 6366 9266
rect 5070 9202 5122 9214
rect 7198 9202 7250 9214
rect 8206 9266 8258 9278
rect 8206 9202 8258 9214
rect 9102 9266 9154 9278
rect 9102 9202 9154 9214
rect 11678 9266 11730 9278
rect 11678 9202 11730 9214
rect 13246 9266 13298 9278
rect 13246 9202 13298 9214
rect 13694 9266 13746 9278
rect 13694 9202 13746 9214
rect 14702 9266 14754 9278
rect 14702 9202 14754 9214
rect 14814 9266 14866 9278
rect 14814 9202 14866 9214
rect 15934 9266 15986 9278
rect 15934 9202 15986 9214
rect 16158 9266 16210 9278
rect 16158 9202 16210 9214
rect 17054 9266 17106 9278
rect 21310 9266 21362 9278
rect 22542 9266 22594 9278
rect 19954 9214 19966 9266
rect 20018 9214 20030 9266
rect 21746 9214 21758 9266
rect 21810 9214 21822 9266
rect 17054 9202 17106 9214
rect 21310 9202 21362 9214
rect 22542 9202 22594 9214
rect 23998 9266 24050 9278
rect 23998 9202 24050 9214
rect 28366 9266 28418 9278
rect 40910 9266 40962 9278
rect 40338 9214 40350 9266
rect 40402 9214 40414 9266
rect 28366 9202 28418 9214
rect 40910 9202 40962 9214
rect 41806 9266 41858 9278
rect 41806 9202 41858 9214
rect 46062 9266 46114 9278
rect 46062 9202 46114 9214
rect 46846 9266 46898 9278
rect 46846 9202 46898 9214
rect 47406 9266 47458 9278
rect 47406 9202 47458 9214
rect 47854 9266 47906 9278
rect 47854 9202 47906 9214
rect 48302 9266 48354 9278
rect 48302 9202 48354 9214
rect 48638 9266 48690 9278
rect 48638 9202 48690 9214
rect 49534 9266 49586 9278
rect 49534 9202 49586 9214
rect 49982 9266 50034 9278
rect 49982 9202 50034 9214
rect 51102 9266 51154 9278
rect 51102 9202 51154 9214
rect 51550 9266 51602 9278
rect 51550 9202 51602 9214
rect 52894 9266 52946 9278
rect 52894 9202 52946 9214
rect 53678 9266 53730 9278
rect 53678 9202 53730 9214
rect 54350 9266 54402 9278
rect 54350 9202 54402 9214
rect 54686 9266 54738 9278
rect 54686 9202 54738 9214
rect 55134 9266 55186 9278
rect 55134 9202 55186 9214
rect 55694 9266 55746 9278
rect 55694 9202 55746 9214
rect 56142 9266 56194 9278
rect 56142 9202 56194 9214
rect 1934 9154 1986 9166
rect 9774 9154 9826 9166
rect 6514 9102 6526 9154
rect 6578 9102 6590 9154
rect 1934 9090 1986 9102
rect 9774 9090 9826 9102
rect 12574 9154 12626 9166
rect 12574 9090 12626 9102
rect 14030 9154 14082 9166
rect 14030 9090 14082 9102
rect 14926 9154 14978 9166
rect 14926 9090 14978 9102
rect 15822 9154 15874 9166
rect 42590 9154 42642 9166
rect 18162 9102 18174 9154
rect 18226 9102 18238 9154
rect 15822 9090 15874 9102
rect 42590 9090 42642 9102
rect 57486 9154 57538 9166
rect 57486 9090 57538 9102
rect 2830 9042 2882 9054
rect 10334 9042 10386 9054
rect 6402 8990 6414 9042
rect 6466 8990 6478 9042
rect 2830 8978 2882 8990
rect 10334 8978 10386 8990
rect 10894 9042 10946 9054
rect 10894 8978 10946 8990
rect 12238 9042 12290 9054
rect 19630 9042 19682 9054
rect 15250 8990 15262 9042
rect 15314 8990 15326 9042
rect 18050 8990 18062 9042
rect 18114 8990 18126 9042
rect 19170 8990 19182 9042
rect 19234 8990 19246 9042
rect 12238 8978 12290 8990
rect 19630 8978 19682 8990
rect 22094 9042 22146 9054
rect 22094 8978 22146 8990
rect 25790 9042 25842 9054
rect 25790 8978 25842 8990
rect 26014 9042 26066 9054
rect 26910 9042 26962 9054
rect 26338 8990 26350 9042
rect 26402 8990 26414 9042
rect 26014 8978 26066 8990
rect 26910 8978 26962 8990
rect 27134 9042 27186 9054
rect 27134 8978 27186 8990
rect 37438 9042 37490 9054
rect 45502 9042 45554 9054
rect 37762 8990 37774 9042
rect 37826 8990 37838 9042
rect 44818 8990 44830 9042
rect 44882 8990 44894 9042
rect 57698 8990 57710 9042
rect 57762 8990 57774 9042
rect 37438 8978 37490 8990
rect 45502 8978 45554 8990
rect 2382 8930 2434 8942
rect 2382 8866 2434 8878
rect 3278 8930 3330 8942
rect 3278 8866 3330 8878
rect 4510 8930 4562 8942
rect 4510 8866 4562 8878
rect 5518 8930 5570 8942
rect 5518 8866 5570 8878
rect 7758 8930 7810 8942
rect 7758 8866 7810 8878
rect 8542 8930 8594 8942
rect 8542 8866 8594 8878
rect 16494 8930 16546 8942
rect 20750 8930 20802 8942
rect 18274 8878 18286 8930
rect 18338 8878 18350 8930
rect 16494 8866 16546 8878
rect 20750 8866 20802 8878
rect 22990 8930 23042 8942
rect 22990 8866 23042 8878
rect 23438 8930 23490 8942
rect 24558 8930 24610 8942
rect 23650 8878 23662 8930
rect 23714 8878 23726 8930
rect 23438 8866 23490 8878
rect 2930 8766 2942 8818
rect 2994 8815 3006 8818
rect 3266 8815 3278 8818
rect 2994 8769 3278 8815
rect 2994 8766 3006 8769
rect 3266 8766 3278 8769
rect 3330 8766 3342 8818
rect 23665 8815 23711 8878
rect 24558 8866 24610 8878
rect 25902 8930 25954 8942
rect 25902 8866 25954 8878
rect 27918 8930 27970 8942
rect 27918 8866 27970 8878
rect 36878 8930 36930 8942
rect 36878 8866 36930 8878
rect 46398 8930 46450 8942
rect 46398 8866 46450 8878
rect 50430 8930 50482 8942
rect 50430 8866 50482 8878
rect 51886 8930 51938 8942
rect 51886 8866 51938 8878
rect 52334 8930 52386 8942
rect 52334 8866 52386 8878
rect 53230 8930 53282 8942
rect 53230 8866 53282 8878
rect 56702 8930 56754 8942
rect 56702 8866 56754 8878
rect 24546 8815 24558 8818
rect 23665 8769 24558 8815
rect 24546 8766 24558 8769
rect 24610 8766 24622 8818
rect 27458 8766 27470 8818
rect 27522 8766 27534 8818
rect 27906 8766 27918 8818
rect 27970 8815 27982 8818
rect 28242 8815 28254 8818
rect 27970 8769 28254 8815
rect 27970 8766 27982 8769
rect 28242 8766 28254 8769
rect 28306 8766 28318 8818
rect 1344 8650 58576 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 58576 8650
rect 1344 8564 58576 8598
rect 57810 8430 57822 8482
rect 57874 8479 57886 8482
rect 58034 8479 58046 8482
rect 57874 8433 58046 8479
rect 57874 8430 57886 8433
rect 58034 8430 58046 8433
rect 58098 8430 58110 8482
rect 1822 8370 1874 8382
rect 1822 8306 1874 8318
rect 2830 8370 2882 8382
rect 2830 8306 2882 8318
rect 3614 8370 3666 8382
rect 3614 8306 3666 8318
rect 4062 8370 4114 8382
rect 4062 8306 4114 8318
rect 4510 8370 4562 8382
rect 4510 8306 4562 8318
rect 5070 8370 5122 8382
rect 5070 8306 5122 8318
rect 6862 8370 6914 8382
rect 12798 8370 12850 8382
rect 11666 8318 11678 8370
rect 11730 8318 11742 8370
rect 6862 8306 6914 8318
rect 12798 8306 12850 8318
rect 15822 8370 15874 8382
rect 15822 8306 15874 8318
rect 16158 8370 16210 8382
rect 16158 8306 16210 8318
rect 16718 8370 16770 8382
rect 20638 8370 20690 8382
rect 17938 8318 17950 8370
rect 18002 8318 18014 8370
rect 18386 8318 18398 8370
rect 18450 8318 18462 8370
rect 16718 8306 16770 8318
rect 20638 8306 20690 8318
rect 21758 8370 21810 8382
rect 21758 8306 21810 8318
rect 24670 8370 24722 8382
rect 24670 8306 24722 8318
rect 42254 8370 42306 8382
rect 42254 8306 42306 8318
rect 42814 8370 42866 8382
rect 42814 8306 42866 8318
rect 43262 8370 43314 8382
rect 43262 8306 43314 8318
rect 43598 8370 43650 8382
rect 43598 8306 43650 8318
rect 44158 8370 44210 8382
rect 44158 8306 44210 8318
rect 44830 8370 44882 8382
rect 44830 8306 44882 8318
rect 50430 8370 50482 8382
rect 50430 8306 50482 8318
rect 50878 8370 50930 8382
rect 50878 8306 50930 8318
rect 51662 8370 51714 8382
rect 51662 8306 51714 8318
rect 52558 8370 52610 8382
rect 52558 8306 52610 8318
rect 53342 8370 53394 8382
rect 53342 8306 53394 8318
rect 53790 8370 53842 8382
rect 56590 8370 56642 8382
rect 55346 8318 55358 8370
rect 55410 8318 55422 8370
rect 53790 8306 53842 8318
rect 56590 8306 56642 8318
rect 57150 8370 57202 8382
rect 57150 8306 57202 8318
rect 6750 8258 6802 8270
rect 49982 8258 50034 8270
rect 6402 8206 6414 8258
rect 6466 8206 6478 8258
rect 7634 8206 7646 8258
rect 7698 8206 7710 8258
rect 8754 8206 8766 8258
rect 8818 8206 8830 8258
rect 10210 8206 10222 8258
rect 10274 8206 10286 8258
rect 10770 8206 10782 8258
rect 10834 8206 10846 8258
rect 17490 8206 17502 8258
rect 17554 8206 17566 8258
rect 18610 8206 18622 8258
rect 18674 8206 18686 8258
rect 19282 8206 19294 8258
rect 19346 8206 19358 8258
rect 26674 8206 26686 8258
rect 26738 8206 26750 8258
rect 38210 8206 38222 8258
rect 38274 8206 38286 8258
rect 38658 8206 38670 8258
rect 38722 8206 38734 8258
rect 45490 8206 45502 8258
rect 45554 8206 45566 8258
rect 45938 8206 45950 8258
rect 46002 8206 46014 8258
rect 6750 8194 6802 8206
rect 49982 8194 50034 8206
rect 51214 8258 51266 8270
rect 56130 8206 56142 8258
rect 56194 8206 56206 8258
rect 51214 8194 51266 8206
rect 23102 8146 23154 8158
rect 7410 8094 7422 8146
rect 7474 8094 7486 8146
rect 11778 8094 11790 8146
rect 11842 8094 11854 8146
rect 14018 8094 14030 8146
rect 14082 8094 14094 8146
rect 14690 8094 14702 8146
rect 14754 8094 14766 8146
rect 23102 8082 23154 8094
rect 23438 8146 23490 8158
rect 23438 8082 23490 8094
rect 25566 8146 25618 8158
rect 25566 8082 25618 8094
rect 26462 8146 26514 8158
rect 26462 8082 26514 8094
rect 41022 8146 41074 8158
rect 41022 8082 41074 8094
rect 41806 8146 41858 8158
rect 41806 8082 41858 8094
rect 52110 8146 52162 8158
rect 52110 8082 52162 8094
rect 2382 8034 2434 8046
rect 2382 7970 2434 7982
rect 3166 8034 3218 8046
rect 3166 7970 3218 7982
rect 13694 8034 13746 8046
rect 13694 7970 13746 7982
rect 15038 8034 15090 8046
rect 20078 8034 20130 8046
rect 19506 7982 19518 8034
rect 19570 7982 19582 8034
rect 15038 7970 15090 7982
rect 20078 7970 20130 7982
rect 22206 8034 22258 8046
rect 23886 8034 23938 8046
rect 22530 7982 22542 8034
rect 22594 7982 22606 8034
rect 22206 7970 22258 7982
rect 23886 7970 23938 7982
rect 25230 8034 25282 8046
rect 25230 7970 25282 7982
rect 27246 8034 27298 8046
rect 27246 7970 27298 7982
rect 27694 8034 27746 8046
rect 27694 7970 27746 7982
rect 37662 8034 37714 8046
rect 49086 8034 49138 8046
rect 48290 7982 48302 8034
rect 48354 7982 48366 8034
rect 37662 7970 37714 7982
rect 49086 7970 49138 7982
rect 49422 8034 49474 8046
rect 49422 7970 49474 7982
rect 54238 8034 54290 8046
rect 54238 7970 54290 7982
rect 57598 8034 57650 8046
rect 57598 7970 57650 7982
rect 58046 8034 58098 8046
rect 58046 7970 58098 7982
rect 1344 7866 58576 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 58576 7866
rect 1344 7780 58576 7814
rect 2494 7698 2546 7710
rect 2494 7634 2546 7646
rect 2942 7698 2994 7710
rect 2942 7634 2994 7646
rect 4286 7698 4338 7710
rect 4286 7634 4338 7646
rect 4622 7698 4674 7710
rect 6526 7698 6578 7710
rect 5170 7646 5182 7698
rect 5234 7646 5246 7698
rect 4622 7634 4674 7646
rect 6526 7634 6578 7646
rect 7310 7698 7362 7710
rect 7310 7634 7362 7646
rect 8990 7698 9042 7710
rect 8990 7634 9042 7646
rect 13582 7698 13634 7710
rect 15150 7698 15202 7710
rect 19854 7698 19906 7710
rect 14242 7646 14254 7698
rect 14306 7646 14318 7698
rect 17826 7646 17838 7698
rect 17890 7646 17902 7698
rect 13582 7634 13634 7646
rect 15150 7634 15202 7646
rect 19854 7634 19906 7646
rect 20862 7698 20914 7710
rect 20862 7634 20914 7646
rect 23886 7698 23938 7710
rect 23886 7634 23938 7646
rect 24894 7698 24946 7710
rect 24894 7634 24946 7646
rect 25678 7698 25730 7710
rect 25678 7634 25730 7646
rect 26910 7698 26962 7710
rect 26910 7634 26962 7646
rect 37998 7698 38050 7710
rect 37998 7634 38050 7646
rect 38334 7698 38386 7710
rect 38334 7634 38386 7646
rect 39118 7698 39170 7710
rect 39118 7634 39170 7646
rect 39566 7698 39618 7710
rect 39566 7634 39618 7646
rect 40462 7698 40514 7710
rect 40462 7634 40514 7646
rect 40910 7698 40962 7710
rect 40910 7634 40962 7646
rect 47294 7698 47346 7710
rect 47294 7634 47346 7646
rect 47854 7698 47906 7710
rect 47854 7634 47906 7646
rect 48526 7698 48578 7710
rect 48526 7634 48578 7646
rect 49534 7698 49586 7710
rect 49534 7634 49586 7646
rect 49870 7698 49922 7710
rect 49870 7634 49922 7646
rect 50318 7698 50370 7710
rect 50318 7634 50370 7646
rect 51662 7698 51714 7710
rect 51662 7634 51714 7646
rect 52334 7698 52386 7710
rect 52334 7634 52386 7646
rect 52782 7698 52834 7710
rect 52782 7634 52834 7646
rect 53230 7698 53282 7710
rect 53230 7634 53282 7646
rect 54014 7698 54066 7710
rect 54014 7634 54066 7646
rect 54350 7698 54402 7710
rect 54350 7634 54402 7646
rect 54798 7698 54850 7710
rect 54798 7634 54850 7646
rect 56590 7698 56642 7710
rect 56590 7634 56642 7646
rect 57374 7698 57426 7710
rect 57374 7634 57426 7646
rect 2046 7586 2098 7598
rect 2046 7522 2098 7534
rect 6638 7586 6690 7598
rect 6638 7522 6690 7534
rect 7534 7586 7586 7598
rect 7534 7522 7586 7534
rect 7758 7586 7810 7598
rect 21870 7586 21922 7598
rect 8642 7534 8654 7586
rect 8706 7534 8718 7586
rect 12114 7534 12126 7586
rect 12178 7534 12190 7586
rect 7758 7522 7810 7534
rect 21870 7522 21922 7534
rect 26126 7586 26178 7598
rect 26126 7522 26178 7534
rect 26462 7586 26514 7598
rect 26462 7522 26514 7534
rect 55246 7586 55298 7598
rect 55246 7522 55298 7534
rect 5518 7474 5570 7486
rect 6414 7474 6466 7486
rect 6066 7422 6078 7474
rect 6130 7422 6142 7474
rect 5518 7410 5570 7422
rect 6414 7410 6466 7422
rect 7086 7474 7138 7486
rect 13694 7474 13746 7486
rect 10322 7422 10334 7474
rect 10386 7422 10398 7474
rect 11442 7422 11454 7474
rect 11506 7422 11518 7474
rect 7086 7410 7138 7422
rect 13694 7410 13746 7422
rect 14590 7474 14642 7486
rect 14590 7410 14642 7422
rect 16382 7474 16434 7486
rect 16382 7410 16434 7422
rect 16942 7474 16994 7486
rect 16942 7410 16994 7422
rect 18174 7474 18226 7486
rect 18174 7410 18226 7422
rect 19070 7474 19122 7486
rect 19070 7410 19122 7422
rect 19294 7474 19346 7486
rect 24558 7474 24610 7486
rect 21634 7422 21646 7474
rect 21698 7422 21710 7474
rect 22754 7422 22766 7474
rect 22818 7422 22830 7474
rect 45714 7422 45726 7474
rect 45778 7422 45790 7474
rect 19294 7410 19346 7422
rect 24558 7410 24610 7422
rect 3390 7362 3442 7374
rect 3390 7298 3442 7310
rect 3838 7362 3890 7374
rect 13022 7362 13074 7374
rect 10546 7310 10558 7362
rect 10610 7310 10622 7362
rect 12674 7310 12686 7362
rect 12738 7310 12750 7362
rect 3838 7298 3890 7310
rect 13022 7298 13074 7310
rect 15710 7362 15762 7374
rect 15710 7298 15762 7310
rect 20302 7362 20354 7374
rect 23438 7362 23490 7374
rect 22530 7310 22542 7362
rect 22594 7310 22606 7362
rect 20302 7298 20354 7310
rect 23438 7298 23490 7310
rect 40014 7362 40066 7374
rect 50878 7362 50930 7374
rect 42130 7310 42142 7362
rect 42194 7310 42206 7362
rect 40014 7298 40066 7310
rect 50878 7298 50930 7310
rect 55694 7362 55746 7374
rect 55694 7298 55746 7310
rect 57822 7362 57874 7374
rect 57822 7298 57874 7310
rect 3378 7198 3390 7250
rect 3442 7247 3454 7250
rect 4498 7247 4510 7250
rect 3442 7201 4510 7247
rect 3442 7198 3454 7201
rect 4498 7198 4510 7201
rect 4562 7198 4574 7250
rect 18722 7198 18734 7250
rect 18786 7198 18798 7250
rect 1344 7082 58576 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 58576 7082
rect 1344 6996 58576 7030
rect 9550 6914 9602 6926
rect 6738 6862 6750 6914
rect 6802 6862 6814 6914
rect 9550 6850 9602 6862
rect 9886 6914 9938 6926
rect 9886 6850 9938 6862
rect 15038 6914 15090 6926
rect 15038 6850 15090 6862
rect 19294 6914 19346 6926
rect 19294 6850 19346 6862
rect 5742 6802 5794 6814
rect 5742 6738 5794 6750
rect 8430 6802 8482 6814
rect 8430 6738 8482 6750
rect 11566 6802 11618 6814
rect 20974 6802 21026 6814
rect 51774 6802 51826 6814
rect 12226 6750 12238 6802
rect 12290 6750 12302 6802
rect 17266 6750 17278 6802
rect 17330 6750 17342 6802
rect 24322 6750 24334 6802
rect 24386 6750 24398 6802
rect 43698 6750 43710 6802
rect 43762 6750 43774 6802
rect 11566 6738 11618 6750
rect 20974 6738 21026 6750
rect 51774 6738 51826 6750
rect 52558 6802 52610 6814
rect 52558 6738 52610 6750
rect 56254 6802 56306 6814
rect 56254 6738 56306 6750
rect 1934 6690 1986 6702
rect 3278 6690 3330 6702
rect 2594 6638 2606 6690
rect 2658 6638 2670 6690
rect 1934 6626 1986 6638
rect 3278 6626 3330 6638
rect 4174 6690 4226 6702
rect 4174 6626 4226 6638
rect 6414 6690 6466 6702
rect 12910 6690 12962 6702
rect 7074 6638 7086 6690
rect 7138 6638 7150 6690
rect 12114 6638 12126 6690
rect 12178 6638 12190 6690
rect 6414 6626 6466 6638
rect 12910 6626 12962 6638
rect 13582 6690 13634 6702
rect 19518 6690 19570 6702
rect 16594 6638 16606 6690
rect 16658 6638 16670 6690
rect 17826 6638 17838 6690
rect 17890 6638 17902 6690
rect 13582 6626 13634 6638
rect 19518 6626 19570 6638
rect 22990 6690 23042 6702
rect 23774 6690 23826 6702
rect 23538 6638 23550 6690
rect 23602 6638 23614 6690
rect 22990 6626 23042 6638
rect 23774 6626 23826 6638
rect 38222 6690 38274 6702
rect 50318 6690 50370 6702
rect 38770 6638 38782 6690
rect 38834 6638 38846 6690
rect 45490 6638 45502 6690
rect 45554 6638 45566 6690
rect 45938 6638 45950 6690
rect 46002 6638 46014 6690
rect 38222 6626 38274 6638
rect 50318 6626 50370 6638
rect 50766 6690 50818 6702
rect 50766 6626 50818 6638
rect 51214 6690 51266 6702
rect 51214 6626 51266 6638
rect 53454 6690 53506 6702
rect 53454 6626 53506 6638
rect 54014 6690 54066 6702
rect 54014 6626 54066 6638
rect 54910 6690 54962 6702
rect 54910 6626 54962 6638
rect 55806 6690 55858 6702
rect 55806 6626 55858 6638
rect 56702 6690 56754 6702
rect 56702 6626 56754 6638
rect 57262 6690 57314 6702
rect 57262 6626 57314 6638
rect 58046 6690 58098 6702
rect 58046 6626 58098 6638
rect 4510 6578 4562 6590
rect 4510 6514 4562 6526
rect 10110 6578 10162 6590
rect 10110 6514 10162 6526
rect 10670 6578 10722 6590
rect 10670 6514 10722 6526
rect 11006 6578 11058 6590
rect 11006 6514 11058 6526
rect 14030 6578 14082 6590
rect 14030 6514 14082 6526
rect 14254 6578 14306 6590
rect 14254 6514 14306 6526
rect 15150 6578 15202 6590
rect 15150 6514 15202 6526
rect 16382 6578 16434 6590
rect 16382 6514 16434 6526
rect 18062 6578 18114 6590
rect 18062 6514 18114 6526
rect 20078 6578 20130 6590
rect 21758 6578 21810 6590
rect 20402 6526 20414 6578
rect 20466 6526 20478 6578
rect 20078 6514 20130 6526
rect 21758 6514 21810 6526
rect 22094 6578 22146 6590
rect 22094 6514 22146 6526
rect 23886 6578 23938 6590
rect 23886 6514 23938 6526
rect 24894 6578 24946 6590
rect 24894 6514 24946 6526
rect 25230 6578 25282 6590
rect 25230 6514 25282 6526
rect 25678 6578 25730 6590
rect 25678 6514 25730 6526
rect 26126 6578 26178 6590
rect 44494 6578 44546 6590
rect 42578 6526 42590 6578
rect 42642 6526 42654 6578
rect 26126 6514 26178 6526
rect 44494 6514 44546 6526
rect 48302 6578 48354 6590
rect 48302 6514 48354 6526
rect 49422 6578 49474 6590
rect 49422 6514 49474 6526
rect 49870 6578 49922 6590
rect 49870 6514 49922 6526
rect 54462 6578 54514 6590
rect 54462 6514 54514 6526
rect 55358 6578 55410 6590
rect 55358 6514 55410 6526
rect 2382 6466 2434 6478
rect 2382 6402 2434 6414
rect 3726 6466 3778 6478
rect 3726 6402 3778 6414
rect 5070 6466 5122 6478
rect 5070 6402 5122 6414
rect 7870 6466 7922 6478
rect 7870 6402 7922 6414
rect 8990 6466 9042 6478
rect 8990 6402 9042 6414
rect 13918 6466 13970 6478
rect 13918 6402 13970 6414
rect 15710 6466 15762 6478
rect 22542 6466 22594 6478
rect 18946 6414 18958 6466
rect 19010 6414 19022 6466
rect 15710 6402 15762 6414
rect 22542 6402 22594 6414
rect 26574 6466 26626 6478
rect 26574 6402 26626 6414
rect 37774 6466 37826 6478
rect 41918 6466 41970 6478
rect 41346 6414 41358 6466
rect 41410 6414 41422 6466
rect 37774 6402 37826 6414
rect 41918 6402 41970 6414
rect 49086 6466 49138 6478
rect 49086 6402 49138 6414
rect 52222 6466 52274 6478
rect 52222 6402 52274 6414
rect 57598 6466 57650 6478
rect 57598 6402 57650 6414
rect 1344 6298 58576 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 58576 6298
rect 1344 6212 58576 6246
rect 3950 6130 4002 6142
rect 3950 6066 4002 6078
rect 4510 6130 4562 6142
rect 4510 6066 4562 6078
rect 4958 6130 5010 6142
rect 4958 6066 5010 6078
rect 5294 6130 5346 6142
rect 5294 6066 5346 6078
rect 5742 6130 5794 6142
rect 5742 6066 5794 6078
rect 6302 6130 6354 6142
rect 6302 6066 6354 6078
rect 6750 6130 6802 6142
rect 6750 6066 6802 6078
rect 7310 6130 7362 6142
rect 7310 6066 7362 6078
rect 8542 6130 8594 6142
rect 8542 6066 8594 6078
rect 10334 6130 10386 6142
rect 10334 6066 10386 6078
rect 11342 6130 11394 6142
rect 13694 6130 13746 6142
rect 12226 6078 12238 6130
rect 12290 6078 12302 6130
rect 12786 6078 12798 6130
rect 12850 6078 12862 6130
rect 11342 6066 11394 6078
rect 13694 6066 13746 6078
rect 14142 6130 14194 6142
rect 14142 6066 14194 6078
rect 15150 6130 15202 6142
rect 15150 6066 15202 6078
rect 15710 6130 15762 6142
rect 15710 6066 15762 6078
rect 16270 6130 16322 6142
rect 16270 6066 16322 6078
rect 18398 6130 18450 6142
rect 18398 6066 18450 6078
rect 19406 6130 19458 6142
rect 19406 6066 19458 6078
rect 20638 6130 20690 6142
rect 20638 6066 20690 6078
rect 21086 6130 21138 6142
rect 21086 6066 21138 6078
rect 22318 6130 22370 6142
rect 22318 6066 22370 6078
rect 22766 6130 22818 6142
rect 22766 6066 22818 6078
rect 23438 6130 23490 6142
rect 23438 6066 23490 6078
rect 25566 6130 25618 6142
rect 25566 6066 25618 6078
rect 36318 6130 36370 6142
rect 45166 6130 45218 6142
rect 40338 6078 40350 6130
rect 40402 6078 40414 6130
rect 44594 6078 44606 6130
rect 44658 6078 44670 6130
rect 36318 6066 36370 6078
rect 45166 6066 45218 6078
rect 46510 6130 46562 6142
rect 46510 6066 46562 6078
rect 46958 6130 47010 6142
rect 46958 6066 47010 6078
rect 48190 6130 48242 6142
rect 48190 6066 48242 6078
rect 48526 6130 48578 6142
rect 48526 6066 48578 6078
rect 53118 6130 53170 6142
rect 53118 6066 53170 6078
rect 53566 6130 53618 6142
rect 53566 6066 53618 6078
rect 54238 6130 54290 6142
rect 54238 6066 54290 6078
rect 54686 6130 54738 6142
rect 54686 6066 54738 6078
rect 55134 6130 55186 6142
rect 55134 6066 55186 6078
rect 55582 6130 55634 6142
rect 55582 6066 55634 6078
rect 56478 6130 56530 6142
rect 56478 6066 56530 6078
rect 57486 6130 57538 6142
rect 57486 6066 57538 6078
rect 57822 6130 57874 6142
rect 57822 6066 57874 6078
rect 10782 6018 10834 6030
rect 10782 5954 10834 5966
rect 13134 6018 13186 6030
rect 13134 5954 13186 5966
rect 24334 6018 24386 6030
rect 24334 5954 24386 5966
rect 45950 6018 46002 6030
rect 45950 5954 46002 5966
rect 52334 6018 52386 6030
rect 52334 5954 52386 5966
rect 23774 5906 23826 5918
rect 2818 5854 2830 5906
rect 2882 5854 2894 5906
rect 12002 5854 12014 5906
rect 12066 5854 12078 5906
rect 19618 5854 19630 5906
rect 19682 5854 19694 5906
rect 23774 5842 23826 5854
rect 24670 5906 24722 5918
rect 24670 5842 24722 5854
rect 37438 5906 37490 5918
rect 41470 5906 41522 5918
rect 45614 5906 45666 5918
rect 37762 5854 37774 5906
rect 37826 5854 37838 5906
rect 42018 5854 42030 5906
rect 42082 5854 42094 5906
rect 37438 5842 37490 5854
rect 41470 5842 41522 5854
rect 45614 5842 45666 5854
rect 49422 5906 49474 5918
rect 49970 5854 49982 5906
rect 50034 5854 50046 5906
rect 49422 5842 49474 5854
rect 3502 5794 3554 5806
rect 1922 5742 1934 5794
rect 1986 5742 1998 5794
rect 3502 5730 3554 5742
rect 7646 5794 7698 5806
rect 7646 5730 7698 5742
rect 8206 5794 8258 5806
rect 8206 5730 8258 5742
rect 9102 5794 9154 5806
rect 14590 5794 14642 5806
rect 9874 5742 9886 5794
rect 9938 5742 9950 5794
rect 9102 5730 9154 5742
rect 14590 5730 14642 5742
rect 16942 5794 16994 5806
rect 16942 5730 16994 5742
rect 17950 5794 18002 5806
rect 17950 5730 18002 5742
rect 18846 5794 18898 5806
rect 18846 5730 18898 5742
rect 21646 5794 21698 5806
rect 21646 5730 21698 5742
rect 36878 5794 36930 5806
rect 36878 5730 36930 5742
rect 47294 5794 47346 5806
rect 47294 5730 47346 5742
rect 55918 5794 55970 5806
rect 55918 5730 55970 5742
rect 40910 5682 40962 5694
rect 13458 5630 13470 5682
rect 13522 5679 13534 5682
rect 14578 5679 14590 5682
rect 13522 5633 14590 5679
rect 13522 5630 13534 5633
rect 14578 5630 14590 5633
rect 14642 5630 14654 5682
rect 40910 5618 40962 5630
rect 1344 5514 58576 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 58576 5514
rect 1344 5428 58576 5462
rect 41134 5346 41186 5358
rect 11106 5294 11118 5346
rect 11170 5343 11182 5346
rect 11330 5343 11342 5346
rect 11170 5297 11342 5343
rect 11170 5294 11182 5297
rect 11330 5294 11342 5297
rect 11394 5294 11406 5346
rect 41134 5282 41186 5294
rect 49086 5346 49138 5358
rect 50754 5294 50766 5346
rect 50818 5343 50830 5346
rect 51202 5343 51214 5346
rect 50818 5297 51214 5343
rect 50818 5294 50830 5297
rect 51202 5294 51214 5297
rect 51266 5294 51278 5346
rect 49086 5282 49138 5294
rect 2158 5234 2210 5246
rect 2158 5170 2210 5182
rect 3390 5234 3442 5246
rect 3390 5170 3442 5182
rect 3726 5234 3778 5246
rect 3726 5170 3778 5182
rect 4510 5234 4562 5246
rect 4510 5170 4562 5182
rect 4958 5234 5010 5246
rect 4958 5170 5010 5182
rect 5854 5234 5906 5246
rect 5854 5170 5906 5182
rect 6302 5234 6354 5246
rect 6302 5170 6354 5182
rect 7310 5234 7362 5246
rect 7310 5170 7362 5182
rect 8206 5234 8258 5246
rect 8206 5170 8258 5182
rect 8766 5234 8818 5246
rect 8766 5170 8818 5182
rect 9214 5234 9266 5246
rect 9214 5170 9266 5182
rect 9662 5234 9714 5246
rect 9662 5170 9714 5182
rect 10110 5234 10162 5246
rect 10110 5170 10162 5182
rect 10558 5234 10610 5246
rect 10558 5170 10610 5182
rect 11118 5234 11170 5246
rect 11118 5170 11170 5182
rect 11566 5234 11618 5246
rect 11566 5170 11618 5182
rect 12910 5234 12962 5246
rect 12910 5170 12962 5182
rect 14030 5234 14082 5246
rect 14030 5170 14082 5182
rect 14814 5234 14866 5246
rect 14814 5170 14866 5182
rect 15374 5234 15426 5246
rect 15374 5170 15426 5182
rect 15822 5234 15874 5246
rect 15822 5170 15874 5182
rect 16270 5234 16322 5246
rect 16270 5170 16322 5182
rect 17838 5234 17890 5246
rect 17838 5170 17890 5182
rect 18286 5234 18338 5246
rect 18286 5170 18338 5182
rect 19070 5234 19122 5246
rect 19070 5170 19122 5182
rect 19518 5234 19570 5246
rect 19518 5170 19570 5182
rect 19966 5234 20018 5246
rect 19966 5170 20018 5182
rect 20862 5234 20914 5246
rect 20862 5170 20914 5182
rect 21534 5234 21586 5246
rect 21534 5170 21586 5182
rect 22094 5234 22146 5246
rect 22094 5170 22146 5182
rect 22990 5234 23042 5246
rect 22990 5170 23042 5182
rect 23662 5234 23714 5246
rect 23662 5170 23714 5182
rect 28814 5234 28866 5246
rect 28814 5170 28866 5182
rect 36430 5234 36482 5246
rect 36430 5170 36482 5182
rect 43934 5234 43986 5246
rect 43934 5170 43986 5182
rect 44718 5234 44770 5246
rect 44718 5170 44770 5182
rect 49870 5234 49922 5246
rect 49870 5170 49922 5182
rect 50318 5234 50370 5246
rect 50318 5170 50370 5182
rect 50766 5234 50818 5246
rect 50766 5170 50818 5182
rect 51102 5234 51154 5246
rect 51102 5170 51154 5182
rect 51662 5234 51714 5246
rect 51662 5170 51714 5182
rect 52110 5234 52162 5246
rect 52110 5170 52162 5182
rect 53342 5234 53394 5246
rect 53342 5170 53394 5182
rect 54238 5234 54290 5246
rect 54238 5170 54290 5182
rect 54574 5234 54626 5246
rect 54574 5170 54626 5182
rect 56702 5234 56754 5246
rect 56702 5170 56754 5182
rect 57150 5234 57202 5246
rect 57150 5170 57202 5182
rect 57598 5234 57650 5246
rect 57598 5170 57650 5182
rect 2606 5122 2658 5134
rect 2606 5058 2658 5070
rect 6862 5122 6914 5134
rect 6862 5058 6914 5070
rect 7870 5122 7922 5134
rect 7870 5058 7922 5070
rect 12238 5122 12290 5134
rect 12238 5058 12290 5070
rect 17278 5122 17330 5134
rect 17278 5058 17330 5070
rect 22430 5122 22482 5134
rect 22430 5058 22482 5070
rect 24110 5122 24162 5134
rect 24110 5058 24162 5070
rect 24894 5122 24946 5134
rect 24894 5058 24946 5070
rect 33854 5122 33906 5134
rect 33854 5058 33906 5070
rect 34638 5122 34690 5134
rect 34638 5058 34690 5070
rect 37438 5122 37490 5134
rect 45614 5122 45666 5134
rect 52446 5122 52498 5134
rect 37986 5070 37998 5122
rect 38050 5070 38062 5122
rect 45938 5070 45950 5122
rect 46002 5070 46014 5122
rect 37438 5058 37490 5070
rect 45614 5058 45666 5070
rect 52446 5058 52498 5070
rect 28366 5010 28418 5022
rect 56254 5010 56306 5022
rect 41906 4958 41918 5010
rect 41970 4958 41982 5010
rect 28366 4946 28418 4958
rect 56254 4946 56306 4958
rect 16830 4898 16882 4910
rect 16830 4834 16882 4846
rect 20302 4898 20354 4910
rect 20302 4834 20354 4846
rect 28030 4898 28082 4910
rect 28030 4834 28082 4846
rect 34190 4898 34242 4910
rect 34190 4834 34242 4846
rect 36878 4898 36930 4910
rect 55022 4898 55074 4910
rect 40562 4846 40574 4898
rect 40626 4846 40638 4898
rect 48514 4846 48526 4898
rect 48578 4846 48590 4898
rect 36878 4834 36930 4846
rect 55022 4834 55074 4846
rect 55918 4898 55970 4910
rect 55918 4834 55970 4846
rect 58046 4898 58098 4910
rect 58046 4834 58098 4846
rect 1344 4730 58576 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 58576 4730
rect 1344 4644 58576 4678
rect 3278 4562 3330 4574
rect 3278 4498 3330 4510
rect 4062 4562 4114 4574
rect 4062 4498 4114 4510
rect 4622 4562 4674 4574
rect 4622 4498 4674 4510
rect 4958 4562 5010 4574
rect 4958 4498 5010 4510
rect 5518 4562 5570 4574
rect 5518 4498 5570 4510
rect 5966 4562 6018 4574
rect 5966 4498 6018 4510
rect 6414 4562 6466 4574
rect 6414 4498 6466 4510
rect 6862 4562 6914 4574
rect 6862 4498 6914 4510
rect 7310 4562 7362 4574
rect 7310 4498 7362 4510
rect 8654 4562 8706 4574
rect 8654 4498 8706 4510
rect 9998 4562 10050 4574
rect 9998 4498 10050 4510
rect 10446 4562 10498 4574
rect 10446 4498 10498 4510
rect 10894 4562 10946 4574
rect 10894 4498 10946 4510
rect 12350 4562 12402 4574
rect 12350 4498 12402 4510
rect 13022 4562 13074 4574
rect 13022 4498 13074 4510
rect 14142 4562 14194 4574
rect 14142 4498 14194 4510
rect 14590 4562 14642 4574
rect 14590 4498 14642 4510
rect 15822 4562 15874 4574
rect 15822 4498 15874 4510
rect 16494 4562 16546 4574
rect 16494 4498 16546 4510
rect 16942 4562 16994 4574
rect 16942 4498 16994 4510
rect 18398 4562 18450 4574
rect 18398 4498 18450 4510
rect 18846 4562 18898 4574
rect 18846 4498 18898 4510
rect 19294 4562 19346 4574
rect 19294 4498 19346 4510
rect 19966 4562 20018 4574
rect 19966 4498 20018 4510
rect 20414 4562 20466 4574
rect 20414 4498 20466 4510
rect 21310 4562 21362 4574
rect 21310 4498 21362 4510
rect 22430 4562 22482 4574
rect 22430 4498 22482 4510
rect 40462 4562 40514 4574
rect 40462 4498 40514 4510
rect 40798 4562 40850 4574
rect 40798 4498 40850 4510
rect 47742 4562 47794 4574
rect 53790 4562 53842 4574
rect 48066 4510 48078 4562
rect 48130 4510 48142 4562
rect 49970 4510 49982 4562
rect 50034 4510 50046 4562
rect 47742 4498 47794 4510
rect 53790 4498 53842 4510
rect 2382 4450 2434 4462
rect 2382 4386 2434 4398
rect 2718 4450 2770 4462
rect 2718 4386 2770 4398
rect 3614 4450 3666 4462
rect 3614 4386 3666 4398
rect 13806 4450 13858 4462
rect 13806 4386 13858 4398
rect 17726 4450 17778 4462
rect 57486 4450 57538 4462
rect 36866 4398 36878 4450
rect 36930 4398 36942 4450
rect 17726 4386 17778 4398
rect 57486 4386 57538 4398
rect 11230 4338 11282 4350
rect 52894 4338 52946 4350
rect 39554 4286 39566 4338
rect 39618 4286 39630 4338
rect 42130 4286 42142 4338
rect 42194 4286 42206 4338
rect 52546 4286 52558 4338
rect 52610 4286 52622 4338
rect 56130 4286 56142 4338
rect 56194 4286 56206 4338
rect 57698 4286 57710 4338
rect 57762 4286 57774 4338
rect 11230 4274 11282 4286
rect 52894 4274 52946 4286
rect 7758 4226 7810 4238
rect 7758 4162 7810 4174
rect 8094 4226 8146 4238
rect 8094 4162 8146 4174
rect 8990 4226 9042 4238
rect 8990 4162 9042 4174
rect 11678 4226 11730 4238
rect 11678 4162 11730 4174
rect 15374 4226 15426 4238
rect 48750 4226 48802 4238
rect 46722 4174 46734 4226
rect 46786 4174 46798 4226
rect 15374 4162 15426 4174
rect 48750 4162 48802 4174
rect 54126 4226 54178 4238
rect 56590 4226 56642 4238
rect 55346 4174 55358 4226
rect 55410 4174 55422 4226
rect 54126 4162 54178 4174
rect 56590 4162 56642 4174
rect 49422 4114 49474 4126
rect 7746 4062 7758 4114
rect 7810 4111 7822 4114
rect 8082 4111 8094 4114
rect 7810 4065 8094 4111
rect 7810 4062 7822 4065
rect 8082 4062 8094 4065
rect 8146 4062 8158 4114
rect 10546 4062 10558 4114
rect 10610 4111 10622 4114
rect 11666 4111 11678 4114
rect 10610 4065 11678 4111
rect 10610 4062 10622 4065
rect 11666 4062 11678 4065
rect 11730 4062 11742 4114
rect 49422 4050 49474 4062
rect 1344 3946 58576 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 58576 3946
rect 1344 3860 58576 3894
rect 18946 3726 18958 3778
rect 19010 3775 19022 3778
rect 19730 3775 19742 3778
rect 19010 3729 19742 3775
rect 19010 3726 19022 3729
rect 19730 3726 19742 3729
rect 19794 3726 19806 3778
rect 5070 3666 5122 3678
rect 7758 3666 7810 3678
rect 7186 3614 7198 3666
rect 7250 3614 7262 3666
rect 5070 3602 5122 3614
rect 7758 3602 7810 3614
rect 8206 3666 8258 3678
rect 8206 3602 8258 3614
rect 8654 3666 8706 3678
rect 8654 3602 8706 3614
rect 9774 3666 9826 3678
rect 9774 3602 9826 3614
rect 10110 3666 10162 3678
rect 10110 3602 10162 3614
rect 10670 3666 10722 3678
rect 10670 3602 10722 3614
rect 11118 3666 11170 3678
rect 11118 3602 11170 3614
rect 13582 3666 13634 3678
rect 13582 3602 13634 3614
rect 14254 3666 14306 3678
rect 14254 3602 14306 3614
rect 14702 3666 14754 3678
rect 14702 3602 14754 3614
rect 15150 3666 15202 3678
rect 15150 3602 15202 3614
rect 15598 3666 15650 3678
rect 15598 3602 15650 3614
rect 16158 3666 16210 3678
rect 16158 3602 16210 3614
rect 16830 3666 16882 3678
rect 16830 3602 16882 3614
rect 19294 3666 19346 3678
rect 19294 3602 19346 3614
rect 19742 3666 19794 3678
rect 19742 3602 19794 3614
rect 20190 3666 20242 3678
rect 20190 3602 20242 3614
rect 25342 3666 25394 3678
rect 25342 3602 25394 3614
rect 31054 3666 31106 3678
rect 38446 3666 38498 3678
rect 35186 3614 35198 3666
rect 35250 3614 35262 3666
rect 31054 3602 31106 3614
rect 38446 3602 38498 3614
rect 41358 3666 41410 3678
rect 41358 3602 41410 3614
rect 41694 3666 41746 3678
rect 45838 3666 45890 3678
rect 43810 3614 43822 3666
rect 43874 3614 43886 3666
rect 41694 3602 41746 3614
rect 45838 3602 45890 3614
rect 46174 3666 46226 3678
rect 46174 3602 46226 3614
rect 46734 3666 46786 3678
rect 46734 3602 46786 3614
rect 47070 3666 47122 3678
rect 47070 3602 47122 3614
rect 47518 3666 47570 3678
rect 47518 3602 47570 3614
rect 48078 3666 48130 3678
rect 48078 3602 48130 3614
rect 48862 3666 48914 3678
rect 48862 3602 48914 3614
rect 49310 3666 49362 3678
rect 49310 3602 49362 3614
rect 51102 3666 51154 3678
rect 51102 3602 51154 3614
rect 51438 3666 51490 3678
rect 51438 3602 51490 3614
rect 51998 3666 52050 3678
rect 56702 3666 56754 3678
rect 53442 3614 53454 3666
rect 53506 3614 53518 3666
rect 55234 3614 55246 3666
rect 55298 3614 55310 3666
rect 51998 3602 52050 3614
rect 56702 3602 56754 3614
rect 57038 3666 57090 3678
rect 57038 3602 57090 3614
rect 57486 3666 57538 3678
rect 57486 3602 57538 3614
rect 57934 3666 57986 3678
rect 57934 3602 57986 3614
rect 45278 3554 45330 3566
rect 2818 3502 2830 3554
rect 2882 3502 2894 3554
rect 12786 3502 12798 3554
rect 12850 3502 12862 3554
rect 18722 3502 18734 3554
rect 18786 3502 18798 3554
rect 24322 3502 24334 3554
rect 24386 3502 24398 3554
rect 30482 3502 30494 3554
rect 30546 3502 30558 3554
rect 34514 3502 34526 3554
rect 34578 3502 34590 3554
rect 39218 3502 39230 3554
rect 39282 3502 39294 3554
rect 45278 3490 45330 3502
rect 49758 3554 49810 3566
rect 49758 3490 49810 3502
rect 50206 3554 50258 3566
rect 52770 3502 52782 3554
rect 52834 3502 52846 3554
rect 55906 3502 55918 3554
rect 55970 3502 55982 3554
rect 50206 3490 50258 3502
rect 4622 3442 4674 3454
rect 1922 3390 1934 3442
rect 1986 3390 1998 3442
rect 5842 3390 5854 3442
rect 5906 3390 5918 3442
rect 11666 3390 11678 3442
rect 11730 3390 11742 3442
rect 17602 3390 17614 3442
rect 17666 3390 17678 3442
rect 23202 3390 23214 3442
rect 23266 3390 23278 3442
rect 29362 3390 29374 3442
rect 29426 3390 29438 3442
rect 40114 3390 40126 3442
rect 40178 3390 40190 3442
rect 42466 3390 42478 3442
rect 42530 3390 42542 3442
rect 44930 3390 44942 3442
rect 44994 3390 45006 3442
rect 4622 3378 4674 3390
rect 37662 3330 37714 3342
rect 37662 3266 37714 3278
rect 38110 3330 38162 3342
rect 38110 3266 38162 3278
rect 50542 3330 50594 3342
rect 50542 3266 50594 3278
rect 1344 3162 58576 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 58576 3162
rect 1344 3076 58576 3110
<< via1 >>
rect 36990 56590 37042 56642
rect 37886 56590 37938 56642
rect 19838 56422 19890 56474
rect 19942 56422 19994 56474
rect 20046 56422 20098 56474
rect 50558 56422 50610 56474
rect 50662 56422 50714 56474
rect 50766 56422 50818 56474
rect 4734 56254 4786 56306
rect 3054 56142 3106 56194
rect 19518 56142 19570 56194
rect 25902 56142 25954 56194
rect 54238 56142 54290 56194
rect 57822 56142 57874 56194
rect 4174 56030 4226 56082
rect 8878 56030 8930 56082
rect 14366 56030 14418 56082
rect 20638 56030 20690 56082
rect 21422 56030 21474 56082
rect 27022 56030 27074 56082
rect 37214 56030 37266 56082
rect 40910 56030 40962 56082
rect 41246 56030 41298 56082
rect 41582 56030 41634 56082
rect 42926 56030 42978 56082
rect 48862 56030 48914 56082
rect 54686 56030 54738 56082
rect 56702 56030 56754 56082
rect 8094 55918 8146 55970
rect 13918 55918 13970 55970
rect 15150 55918 15202 55970
rect 27582 55918 27634 55970
rect 36430 55918 36482 55970
rect 37886 55918 37938 55970
rect 41134 55918 41186 55970
rect 42478 55918 42530 55970
rect 43710 55918 43762 55970
rect 49534 55918 49586 55970
rect 55470 55918 55522 55970
rect 4478 55638 4530 55690
rect 4582 55638 4634 55690
rect 4686 55638 4738 55690
rect 35198 55638 35250 55690
rect 35302 55638 35354 55690
rect 35406 55638 35458 55690
rect 1934 55358 1986 55410
rect 31390 55358 31442 55410
rect 3054 55246 3106 55298
rect 37774 55246 37826 55298
rect 39790 55246 39842 55298
rect 40238 55246 40290 55298
rect 42590 55246 42642 55298
rect 43710 55246 43762 55298
rect 54350 55246 54402 55298
rect 55134 55246 55186 55298
rect 23326 55134 23378 55186
rect 23662 55134 23714 55186
rect 26798 55134 26850 55186
rect 27134 55134 27186 55186
rect 29598 55134 29650 55186
rect 29934 55134 29986 55186
rect 31950 55134 32002 55186
rect 37550 55134 37602 55186
rect 39342 55134 39394 55186
rect 42254 55134 42306 55186
rect 44158 55134 44210 55186
rect 46622 55134 46674 55186
rect 46958 55134 47010 55186
rect 56030 55134 56082 55186
rect 3502 55022 3554 55074
rect 22878 55022 22930 55074
rect 34414 55022 34466 55074
rect 56590 55022 56642 55074
rect 19838 54854 19890 54906
rect 19942 54854 19994 54906
rect 20046 54854 20098 54906
rect 50558 54854 50610 54906
rect 50662 54854 50714 54906
rect 50766 54854 50818 54906
rect 39678 54686 39730 54738
rect 40574 54686 40626 54738
rect 37550 54574 37602 54626
rect 42142 54574 42194 54626
rect 38222 54462 38274 54514
rect 40798 54462 40850 54514
rect 42478 54462 42530 54514
rect 42702 54462 42754 54514
rect 43262 54462 43314 54514
rect 43710 54462 43762 54514
rect 43822 54462 43874 54514
rect 43934 54462 43986 54514
rect 38446 54350 38498 54402
rect 39118 54350 39170 54402
rect 39342 54350 39394 54402
rect 40462 54350 40514 54402
rect 42254 54350 42306 54402
rect 4478 54070 4530 54122
rect 4582 54070 4634 54122
rect 4686 54070 4738 54122
rect 35198 54070 35250 54122
rect 35302 54070 35354 54122
rect 35406 54070 35458 54122
rect 40462 53790 40514 53842
rect 42814 53790 42866 53842
rect 39006 53678 39058 53730
rect 39342 53678 39394 53730
rect 40350 53678 40402 53730
rect 41582 53678 41634 53730
rect 43150 53678 43202 53730
rect 43486 53678 43538 53730
rect 2718 53566 2770 53618
rect 3166 53566 3218 53618
rect 40462 53566 40514 53618
rect 41694 53566 41746 53618
rect 2382 53454 2434 53506
rect 39118 53454 39170 53506
rect 42478 53454 42530 53506
rect 42926 53454 42978 53506
rect 43934 53454 43986 53506
rect 44382 53454 44434 53506
rect 19838 53286 19890 53338
rect 19942 53286 19994 53338
rect 20046 53286 20098 53338
rect 50558 53286 50610 53338
rect 50662 53286 50714 53338
rect 50766 53286 50818 53338
rect 35086 53118 35138 53170
rect 35982 53118 36034 53170
rect 40910 53118 40962 53170
rect 42030 53118 42082 53170
rect 42814 53118 42866 53170
rect 47070 53118 47122 53170
rect 38894 53006 38946 53058
rect 40686 53006 40738 53058
rect 42590 53006 42642 53058
rect 43038 53006 43090 53058
rect 43598 53006 43650 53058
rect 43822 53006 43874 53058
rect 33630 52894 33682 52946
rect 33966 52894 34018 52946
rect 34190 52894 34242 52946
rect 39230 52894 39282 52946
rect 40574 52894 40626 52946
rect 41470 52894 41522 52946
rect 41806 52894 41858 52946
rect 44382 52894 44434 52946
rect 46846 52894 46898 52946
rect 47182 52894 47234 52946
rect 47406 52894 47458 52946
rect 33742 52782 33794 52834
rect 34750 52782 34802 52834
rect 35646 52782 35698 52834
rect 36542 52782 36594 52834
rect 38334 52782 38386 52834
rect 39790 52782 39842 52834
rect 41694 52782 41746 52834
rect 42702 52782 42754 52834
rect 45054 52782 45106 52834
rect 46398 52782 46450 52834
rect 47966 52782 48018 52834
rect 43710 52670 43762 52722
rect 44158 52670 44210 52722
rect 4478 52502 4530 52554
rect 4582 52502 4634 52554
rect 4686 52502 4738 52554
rect 35198 52502 35250 52554
rect 35302 52502 35354 52554
rect 35406 52502 35458 52554
rect 34862 52334 34914 52386
rect 39006 52334 39058 52386
rect 40798 52334 40850 52386
rect 41806 52334 41858 52386
rect 42030 52334 42082 52386
rect 42814 52334 42866 52386
rect 43262 52334 43314 52386
rect 43934 52334 43986 52386
rect 45950 52334 46002 52386
rect 35086 52222 35138 52274
rect 36654 52222 36706 52274
rect 38334 52222 38386 52274
rect 40462 52222 40514 52274
rect 40910 52222 40962 52274
rect 42478 52222 42530 52274
rect 43710 52222 43762 52274
rect 44158 52222 44210 52274
rect 45390 52222 45442 52274
rect 47070 52222 47122 52274
rect 49310 52222 49362 52274
rect 2830 52110 2882 52162
rect 32510 52110 32562 52162
rect 33182 52110 33234 52162
rect 33854 52110 33906 52162
rect 36430 52110 36482 52162
rect 37438 52110 37490 52162
rect 39118 52110 39170 52162
rect 39790 52110 39842 52162
rect 41358 52110 41410 52162
rect 42254 52110 42306 52162
rect 47630 52110 47682 52162
rect 48750 52110 48802 52162
rect 1934 51998 1986 52050
rect 32734 51998 32786 52050
rect 34526 51998 34578 52050
rect 35870 51998 35922 52050
rect 36094 51998 36146 52050
rect 36206 51998 36258 52050
rect 42590 51998 42642 52050
rect 44382 51998 44434 52050
rect 46510 51998 46562 52050
rect 47518 51998 47570 52050
rect 47742 51998 47794 52050
rect 26798 51886 26850 51938
rect 32622 51886 32674 51938
rect 37886 51886 37938 51938
rect 46062 51886 46114 51938
rect 46286 51886 46338 51938
rect 48414 51886 48466 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 23550 51550 23602 51602
rect 24670 51550 24722 51602
rect 38334 51550 38386 51602
rect 43150 51550 43202 51602
rect 49870 51550 49922 51602
rect 26238 51438 26290 51490
rect 28030 51438 28082 51490
rect 40350 51438 40402 51490
rect 41470 51438 41522 51490
rect 43822 51438 43874 51490
rect 23438 51326 23490 51378
rect 23662 51326 23714 51378
rect 24110 51326 24162 51378
rect 24558 51326 24610 51378
rect 24894 51326 24946 51378
rect 27358 51326 27410 51378
rect 32398 51326 32450 51378
rect 33742 51326 33794 51378
rect 34190 51326 34242 51378
rect 35310 51326 35362 51378
rect 36094 51326 36146 51378
rect 37438 51326 37490 51378
rect 38334 51326 38386 51378
rect 40126 51326 40178 51378
rect 40462 51326 40514 51378
rect 43262 51326 43314 51378
rect 47294 51326 47346 51378
rect 47966 51326 48018 51378
rect 49534 51326 49586 51378
rect 49758 51326 49810 51378
rect 50206 51326 50258 51378
rect 21870 51214 21922 51266
rect 27694 51214 27746 51266
rect 32286 51214 32338 51266
rect 34638 51214 34690 51266
rect 37550 51214 37602 51266
rect 39342 51214 39394 51266
rect 39678 51214 39730 51266
rect 42030 51214 42082 51266
rect 42702 51214 42754 51266
rect 44830 51214 44882 51266
rect 45166 51214 45218 51266
rect 45726 51214 45778 51266
rect 46174 51214 46226 51266
rect 46510 51214 46562 51266
rect 48750 51214 48802 51266
rect 50766 51214 50818 51266
rect 26126 51102 26178 51154
rect 26462 51102 26514 51154
rect 32734 51102 32786 51154
rect 38446 51102 38498 51154
rect 38670 51102 38722 51154
rect 43486 51102 43538 51154
rect 44046 51102 44098 51154
rect 47518 51102 47570 51154
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 36318 50766 36370 50818
rect 37438 50766 37490 50818
rect 37886 50766 37938 50818
rect 38446 50766 38498 50818
rect 40126 50766 40178 50818
rect 47406 50766 47458 50818
rect 48302 50766 48354 50818
rect 49198 50766 49250 50818
rect 49534 50766 49586 50818
rect 50318 50766 50370 50818
rect 50766 50766 50818 50818
rect 51326 50766 51378 50818
rect 24670 50654 24722 50706
rect 27470 50654 27522 50706
rect 37438 50654 37490 50706
rect 38334 50654 38386 50706
rect 39790 50654 39842 50706
rect 42478 50654 42530 50706
rect 48302 50654 48354 50706
rect 50430 50654 50482 50706
rect 50878 50654 50930 50706
rect 51326 50654 51378 50706
rect 22206 50542 22258 50594
rect 22542 50542 22594 50594
rect 22766 50542 22818 50594
rect 24110 50542 24162 50594
rect 26126 50542 26178 50594
rect 26350 50542 26402 50594
rect 36094 50542 36146 50594
rect 36542 50542 36594 50594
rect 36766 50542 36818 50594
rect 37886 50542 37938 50594
rect 39006 50542 39058 50594
rect 41022 50542 41074 50594
rect 42702 50542 42754 50594
rect 43486 50542 43538 50594
rect 44718 50542 44770 50594
rect 45390 50542 45442 50594
rect 9214 50430 9266 50482
rect 25006 50430 25058 50482
rect 27022 50430 27074 50482
rect 34750 50430 34802 50482
rect 35198 50430 35250 50482
rect 39230 50430 39282 50482
rect 39902 50430 39954 50482
rect 42030 50430 42082 50482
rect 42590 50430 42642 50482
rect 43374 50430 43426 50482
rect 45726 50430 45778 50482
rect 49758 50430 49810 50482
rect 52110 50430 52162 50482
rect 8878 50318 8930 50370
rect 23214 50318 23266 50370
rect 31838 50318 31890 50370
rect 33070 50318 33122 50370
rect 33518 50318 33570 50370
rect 35646 50318 35698 50370
rect 40686 50318 40738 50370
rect 41582 50318 41634 50370
rect 45614 50318 45666 50370
rect 46174 50318 46226 50370
rect 46846 50318 46898 50370
rect 47182 50318 47234 50370
rect 47854 50318 47906 50370
rect 48638 50318 48690 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 40910 49982 40962 50034
rect 42366 49982 42418 50034
rect 43598 49982 43650 50034
rect 47518 49982 47570 50034
rect 9774 49870 9826 49922
rect 24222 49870 24274 49922
rect 26798 49870 26850 49922
rect 28142 49870 28194 49922
rect 30046 49870 30098 49922
rect 31614 49870 31666 49922
rect 36094 49870 36146 49922
rect 42254 49870 42306 49922
rect 10446 49758 10498 49810
rect 13246 49758 13298 49810
rect 13470 49758 13522 49810
rect 13918 49758 13970 49810
rect 20638 49758 20690 49810
rect 21534 49758 21586 49810
rect 22206 49758 22258 49810
rect 22430 49758 22482 49810
rect 23662 49758 23714 49810
rect 23998 49758 24050 49810
rect 26574 49758 26626 49810
rect 26686 49758 26738 49810
rect 27694 49758 27746 49810
rect 28254 49758 28306 49810
rect 30270 49758 30322 49810
rect 31166 49758 31218 49810
rect 36206 49758 36258 49810
rect 36430 49758 36482 49810
rect 46846 49758 46898 49810
rect 9998 49646 10050 49698
rect 13358 49646 13410 49698
rect 19966 49646 20018 49698
rect 21198 49646 21250 49698
rect 27918 49646 27970 49698
rect 32062 49646 32114 49698
rect 32510 49646 32562 49698
rect 34190 49646 34242 49698
rect 36990 49646 37042 49698
rect 37438 49646 37490 49698
rect 38894 49646 38946 49698
rect 39342 49646 39394 49698
rect 39790 49646 39842 49698
rect 40462 49646 40514 49698
rect 41470 49646 41522 49698
rect 42926 49646 42978 49698
rect 44158 49646 44210 49698
rect 44606 49646 44658 49698
rect 45166 49646 45218 49698
rect 45502 49646 45554 49698
rect 46286 49646 46338 49698
rect 47406 49646 47458 49698
rect 47966 49646 48018 49698
rect 48638 49646 48690 49698
rect 49534 49646 49586 49698
rect 49982 49646 50034 49698
rect 50318 49646 50370 49698
rect 50766 49646 50818 49698
rect 51326 49646 51378 49698
rect 51998 49646 52050 49698
rect 52446 49646 52498 49698
rect 52894 49646 52946 49698
rect 53230 49646 53282 49698
rect 53790 49646 53842 49698
rect 54238 49646 54290 49698
rect 54574 49646 54626 49698
rect 55134 49646 55186 49698
rect 55470 49646 55522 49698
rect 22542 49534 22594 49586
rect 23438 49534 23490 49586
rect 24110 49534 24162 49586
rect 27246 49534 27298 49586
rect 33630 49534 33682 49586
rect 33966 49534 34018 49586
rect 35646 49534 35698 49586
rect 39006 49534 39058 49586
rect 39566 49534 39618 49586
rect 40014 49534 40066 49586
rect 40238 49534 40290 49586
rect 43934 49534 43986 49586
rect 49422 49534 49474 49586
rect 50318 49534 50370 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 13918 49198 13970 49250
rect 23438 49198 23490 49250
rect 23774 49198 23826 49250
rect 26126 49198 26178 49250
rect 32734 49198 32786 49250
rect 33294 49198 33346 49250
rect 39902 49198 39954 49250
rect 46174 49198 46226 49250
rect 48078 49198 48130 49250
rect 48190 49198 48242 49250
rect 15822 49086 15874 49138
rect 20862 49086 20914 49138
rect 21758 49086 21810 49138
rect 26798 49086 26850 49138
rect 31278 49086 31330 49138
rect 33742 49086 33794 49138
rect 40126 49086 40178 49138
rect 43710 49086 43762 49138
rect 46398 49086 46450 49138
rect 46958 49086 47010 49138
rect 47742 49086 47794 49138
rect 49982 49086 50034 49138
rect 51102 49086 51154 49138
rect 51998 49086 52050 49138
rect 9662 48974 9714 49026
rect 12798 48974 12850 49026
rect 13694 48974 13746 49026
rect 14142 48974 14194 49026
rect 16046 48974 16098 49026
rect 16942 48974 16994 49026
rect 21646 48974 21698 49026
rect 26910 48974 26962 49026
rect 30270 48974 30322 49026
rect 30606 48974 30658 49026
rect 32398 48974 32450 49026
rect 33518 48974 33570 49026
rect 34190 48974 34242 49026
rect 35086 48974 35138 49026
rect 35534 48974 35586 49026
rect 37886 48974 37938 49026
rect 39230 48974 39282 49026
rect 40014 48974 40066 49026
rect 40462 48974 40514 49026
rect 40686 48974 40738 49026
rect 43934 48974 43986 49026
rect 46734 48974 46786 49026
rect 47854 48974 47906 49026
rect 49534 48974 49586 49026
rect 50430 48974 50482 49026
rect 55134 48974 55186 49026
rect 10110 48862 10162 48914
rect 10334 48862 10386 48914
rect 12462 48862 12514 48914
rect 12686 48862 12738 48914
rect 17054 48862 17106 48914
rect 18958 48862 19010 48914
rect 21982 48862 22034 48914
rect 23662 48862 23714 48914
rect 29598 48862 29650 48914
rect 30046 48862 30098 48914
rect 31614 48862 31666 48914
rect 32174 48862 32226 48914
rect 34862 48862 34914 48914
rect 41694 48862 41746 48914
rect 42478 48862 42530 48914
rect 43374 48862 43426 48914
rect 45390 48862 45442 48914
rect 46398 48862 46450 48914
rect 48638 48862 48690 48914
rect 56030 48862 56082 48914
rect 9998 48750 10050 48802
rect 12910 48750 12962 48802
rect 13806 48750 13858 48802
rect 16382 48750 16434 48802
rect 17278 48750 17330 48802
rect 18734 48750 18786 48802
rect 18846 48750 18898 48802
rect 22430 48750 22482 48802
rect 22878 48750 22930 48802
rect 30270 48750 30322 48802
rect 31390 48750 31442 48802
rect 33966 48750 34018 48802
rect 34078 48750 34130 48802
rect 35198 48750 35250 48802
rect 35310 48750 35362 48802
rect 35982 48750 36034 48802
rect 36654 48750 36706 48802
rect 37550 48750 37602 48802
rect 38334 48750 38386 48802
rect 39342 48750 39394 48802
rect 41246 48750 41298 48802
rect 42814 48750 42866 48802
rect 43598 48750 43650 48802
rect 43822 48750 43874 48802
rect 44494 48750 44546 48802
rect 51550 48750 51602 48802
rect 52782 48750 52834 48802
rect 53454 48750 53506 48802
rect 53902 48750 53954 48802
rect 54350 48750 54402 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 3278 48414 3330 48466
rect 9774 48414 9826 48466
rect 17726 48414 17778 48466
rect 17950 48414 18002 48466
rect 21198 48414 21250 48466
rect 21870 48414 21922 48466
rect 31390 48414 31442 48466
rect 32734 48414 32786 48466
rect 34526 48414 34578 48466
rect 37326 48414 37378 48466
rect 39566 48414 39618 48466
rect 40798 48414 40850 48466
rect 43150 48414 43202 48466
rect 47070 48414 47122 48466
rect 47182 48414 47234 48466
rect 48078 48414 48130 48466
rect 51662 48414 51714 48466
rect 52334 48414 52386 48466
rect 54238 48414 54290 48466
rect 2382 48302 2434 48354
rect 2718 48302 2770 48354
rect 10446 48302 10498 48354
rect 11790 48302 11842 48354
rect 12462 48302 12514 48354
rect 14142 48302 14194 48354
rect 18174 48302 18226 48354
rect 18958 48302 19010 48354
rect 21982 48302 22034 48354
rect 24334 48302 24386 48354
rect 27134 48302 27186 48354
rect 27246 48302 27298 48354
rect 30830 48302 30882 48354
rect 35870 48302 35922 48354
rect 48638 48302 48690 48354
rect 51326 48302 51378 48354
rect 52782 48302 52834 48354
rect 9774 48190 9826 48242
rect 9998 48190 10050 48242
rect 10222 48190 10274 48242
rect 11678 48190 11730 48242
rect 12014 48190 12066 48242
rect 13134 48190 13186 48242
rect 13806 48190 13858 48242
rect 16606 48190 16658 48242
rect 18846 48190 18898 48242
rect 19742 48190 19794 48242
rect 23214 48190 23266 48242
rect 23438 48190 23490 48242
rect 24110 48190 24162 48242
rect 24446 48190 24498 48242
rect 26910 48190 26962 48242
rect 29710 48190 29762 48242
rect 30494 48190 30546 48242
rect 31726 48190 31778 48242
rect 35758 48190 35810 48242
rect 36990 48190 37042 48242
rect 39342 48190 39394 48242
rect 40126 48190 40178 48242
rect 40350 48190 40402 48242
rect 40574 48190 40626 48242
rect 40798 48190 40850 48242
rect 46734 48190 46786 48242
rect 46958 48190 47010 48242
rect 47406 48190 47458 48242
rect 47854 48190 47906 48242
rect 48190 48190 48242 48242
rect 50318 48190 50370 48242
rect 51550 48190 51602 48242
rect 51774 48190 51826 48242
rect 53454 48190 53506 48242
rect 15150 48078 15202 48130
rect 15934 48078 15986 48130
rect 16270 48078 16322 48130
rect 17838 48078 17890 48130
rect 19518 48078 19570 48130
rect 23550 48078 23602 48130
rect 24894 48078 24946 48130
rect 26126 48078 26178 48130
rect 29934 48078 29986 48130
rect 32846 48078 32898 48130
rect 33630 48078 33682 48130
rect 34862 48078 34914 48130
rect 38222 48078 38274 48130
rect 38670 48078 38722 48130
rect 41582 48078 41634 48130
rect 41918 48078 41970 48130
rect 42366 48078 42418 48130
rect 43710 48078 43762 48130
rect 44158 48078 44210 48130
rect 44606 48078 44658 48130
rect 45054 48078 45106 48130
rect 45502 48078 45554 48130
rect 46062 48078 46114 48130
rect 49646 48078 49698 48130
rect 49982 48078 50034 48130
rect 53678 48078 53730 48130
rect 54798 48078 54850 48130
rect 55246 48078 55298 48130
rect 55582 48078 55634 48130
rect 56030 48078 56082 48130
rect 56478 48078 56530 48130
rect 57486 48078 57538 48130
rect 21870 47966 21922 48018
rect 26686 47966 26738 48018
rect 27470 47966 27522 48018
rect 29374 47966 29426 48018
rect 32510 47966 32562 48018
rect 33854 47966 33906 48018
rect 34078 47966 34130 48018
rect 35534 47966 35586 48018
rect 36094 47966 36146 48018
rect 36318 47966 36370 48018
rect 43486 47966 43538 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 8990 47630 9042 47682
rect 11454 47630 11506 47682
rect 14478 47630 14530 47682
rect 16606 47630 16658 47682
rect 19630 47630 19682 47682
rect 22318 47630 22370 47682
rect 34750 47630 34802 47682
rect 35086 47630 35138 47682
rect 39118 47630 39170 47682
rect 40238 47630 40290 47682
rect 54238 47630 54290 47682
rect 8766 47518 8818 47570
rect 10334 47518 10386 47570
rect 16718 47518 16770 47570
rect 18286 47518 18338 47570
rect 19518 47518 19570 47570
rect 22878 47518 22930 47570
rect 25566 47518 25618 47570
rect 26462 47518 26514 47570
rect 33742 47518 33794 47570
rect 34750 47518 34802 47570
rect 35198 47518 35250 47570
rect 36766 47518 36818 47570
rect 41694 47518 41746 47570
rect 51662 47518 51714 47570
rect 57038 47518 57090 47570
rect 57486 47518 57538 47570
rect 57934 47518 57986 47570
rect 10446 47406 10498 47458
rect 11454 47406 11506 47458
rect 12238 47406 12290 47458
rect 12686 47406 12738 47458
rect 12910 47406 12962 47458
rect 13806 47406 13858 47458
rect 14030 47406 14082 47458
rect 16270 47406 16322 47458
rect 19294 47406 19346 47458
rect 22654 47406 22706 47458
rect 23438 47406 23490 47458
rect 23774 47406 23826 47458
rect 26014 47406 26066 47458
rect 30046 47406 30098 47458
rect 31166 47406 31218 47458
rect 33294 47406 33346 47458
rect 37550 47406 37602 47458
rect 37774 47406 37826 47458
rect 37998 47406 38050 47458
rect 39454 47406 39506 47458
rect 39678 47406 39730 47458
rect 40686 47406 40738 47458
rect 40910 47406 40962 47458
rect 41134 47406 41186 47458
rect 43038 47406 43090 47458
rect 43486 47406 43538 47458
rect 44046 47406 44098 47458
rect 46510 47406 46562 47458
rect 47854 47406 47906 47458
rect 48862 47406 48914 47458
rect 49646 47406 49698 47458
rect 51550 47406 51602 47458
rect 51886 47406 51938 47458
rect 53566 47406 53618 47458
rect 54014 47406 54066 47458
rect 9886 47294 9938 47346
rect 11790 47294 11842 47346
rect 13918 47294 13970 47346
rect 23550 47294 23602 47346
rect 30942 47294 30994 47346
rect 33630 47294 33682 47346
rect 33854 47294 33906 47346
rect 34302 47294 34354 47346
rect 41022 47294 41074 47346
rect 43710 47294 43762 47346
rect 44382 47294 44434 47346
rect 46846 47294 46898 47346
rect 53454 47294 53506 47346
rect 53790 47294 53842 47346
rect 54910 47294 54962 47346
rect 55246 47294 55298 47346
rect 9326 47182 9378 47234
rect 12574 47182 12626 47234
rect 14926 47182 14978 47234
rect 17950 47182 18002 47234
rect 18174 47182 18226 47234
rect 18398 47182 18450 47234
rect 24110 47182 24162 47234
rect 30158 47182 30210 47234
rect 35646 47182 35698 47234
rect 36318 47182 36370 47234
rect 42254 47182 42306 47234
rect 45390 47182 45442 47234
rect 46062 47182 46114 47234
rect 51326 47182 51378 47234
rect 52558 47182 52610 47234
rect 55694 47182 55746 47234
rect 56142 47182 56194 47234
rect 56590 47182 56642 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 12798 46846 12850 46898
rect 14366 46846 14418 46898
rect 16830 46846 16882 46898
rect 17054 46846 17106 46898
rect 18286 46846 18338 46898
rect 22654 46846 22706 46898
rect 22878 46846 22930 46898
rect 23214 46846 23266 46898
rect 24894 46846 24946 46898
rect 34862 46846 34914 46898
rect 40462 46846 40514 46898
rect 40686 46846 40738 46898
rect 43262 46846 43314 46898
rect 44270 46846 44322 46898
rect 48302 46846 48354 46898
rect 49870 46846 49922 46898
rect 53566 46846 53618 46898
rect 54462 46846 54514 46898
rect 55694 46846 55746 46898
rect 56142 46846 56194 46898
rect 16718 46734 16770 46786
rect 18510 46734 18562 46786
rect 26910 46734 26962 46786
rect 33742 46734 33794 46786
rect 33966 46734 34018 46786
rect 36878 46734 36930 46786
rect 39566 46734 39618 46786
rect 42926 46734 42978 46786
rect 45054 46734 45106 46786
rect 46734 46734 46786 46786
rect 51998 46734 52050 46786
rect 57822 46734 57874 46786
rect 10110 46622 10162 46674
rect 14030 46622 14082 46674
rect 18622 46622 18674 46674
rect 19630 46622 19682 46674
rect 22542 46622 22594 46674
rect 24222 46622 24274 46674
rect 24670 46622 24722 46674
rect 25902 46622 25954 46674
rect 26126 46622 26178 46674
rect 27246 46622 27298 46674
rect 30270 46622 30322 46674
rect 32398 46622 32450 46674
rect 34414 46622 34466 46674
rect 37550 46622 37602 46674
rect 37774 46622 37826 46674
rect 39342 46622 39394 46674
rect 40238 46622 40290 46674
rect 40350 46622 40402 46674
rect 40574 46622 40626 46674
rect 43038 46622 43090 46674
rect 43486 46622 43538 46674
rect 44046 46622 44098 46674
rect 44606 46622 44658 46674
rect 47294 46622 47346 46674
rect 48078 46622 48130 46674
rect 48414 46622 48466 46674
rect 49646 46622 49698 46674
rect 52446 46622 52498 46674
rect 52894 46622 52946 46674
rect 53902 46622 53954 46674
rect 54686 46622 54738 46674
rect 9102 46510 9154 46562
rect 10334 46510 10386 46562
rect 10782 46510 10834 46562
rect 13246 46510 13298 46562
rect 13806 46510 13858 46562
rect 19742 46510 19794 46562
rect 24782 46510 24834 46562
rect 26462 46510 26514 46562
rect 27358 46510 27410 46562
rect 30046 46510 30098 46562
rect 32510 46510 32562 46562
rect 33630 46510 33682 46562
rect 38334 46510 38386 46562
rect 41470 46510 41522 46562
rect 42254 46510 42306 46562
rect 42702 46510 42754 46562
rect 44158 46510 44210 46562
rect 45614 46510 45666 46562
rect 45950 46510 46002 46562
rect 47406 46510 47458 46562
rect 50318 46510 50370 46562
rect 50878 46510 50930 46562
rect 51214 46510 51266 46562
rect 55358 46510 55410 46562
rect 56590 46510 56642 46562
rect 57374 46510 57426 46562
rect 20190 46398 20242 46450
rect 29934 46398 29986 46450
rect 31838 46398 31890 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 12350 46062 12402 46114
rect 13694 46062 13746 46114
rect 19182 46062 19234 46114
rect 23326 46062 23378 46114
rect 25454 46062 25506 46114
rect 52670 46062 52722 46114
rect 57262 46062 57314 46114
rect 58046 46062 58098 46114
rect 6414 45950 6466 46002
rect 10110 45950 10162 46002
rect 22878 45950 22930 46002
rect 26126 45950 26178 46002
rect 27022 45950 27074 46002
rect 29822 45950 29874 46002
rect 35310 45950 35362 46002
rect 41694 45950 41746 46002
rect 42926 45950 42978 46002
rect 43710 45950 43762 46002
rect 46958 45950 47010 46002
rect 47182 45950 47234 46002
rect 48862 45950 48914 46002
rect 50318 45950 50370 46002
rect 50766 45950 50818 46002
rect 51214 45950 51266 46002
rect 57262 45950 57314 46002
rect 2830 45838 2882 45890
rect 12686 45838 12738 45890
rect 14030 45838 14082 45890
rect 14254 45838 14306 45890
rect 22990 45838 23042 45890
rect 24894 45838 24946 45890
rect 25118 45838 25170 45890
rect 26574 45838 26626 45890
rect 28254 45838 28306 45890
rect 28478 45838 28530 45890
rect 28926 45838 28978 45890
rect 29934 45838 29986 45890
rect 37774 45838 37826 45890
rect 39118 45838 39170 45890
rect 43486 45838 43538 45890
rect 46622 45838 46674 45890
rect 47518 45838 47570 45890
rect 48414 45838 48466 45890
rect 49758 45838 49810 45890
rect 1934 45726 1986 45778
rect 5854 45726 5906 45778
rect 5966 45726 6018 45778
rect 9102 45726 9154 45778
rect 12910 45726 12962 45778
rect 19518 45726 19570 45778
rect 19966 45726 20018 45778
rect 30606 45726 30658 45778
rect 36654 45726 36706 45778
rect 40014 45726 40066 45778
rect 40350 45726 40402 45778
rect 45726 45726 45778 45778
rect 47966 45726 48018 45778
rect 49534 45726 49586 45778
rect 52558 45726 52610 45778
rect 53454 45726 53506 45778
rect 5630 45614 5682 45666
rect 7310 45614 7362 45666
rect 8206 45614 8258 45666
rect 10558 45614 10610 45666
rect 11118 45614 11170 45666
rect 11790 45614 11842 45666
rect 14702 45614 14754 45666
rect 19294 45614 19346 45666
rect 28366 45614 28418 45666
rect 33070 45614 33122 45666
rect 33630 45614 33682 45666
rect 37438 45614 37490 45666
rect 37662 45614 37714 45666
rect 38222 45614 38274 45666
rect 38782 45614 38834 45666
rect 40798 45614 40850 45666
rect 41246 45614 41298 45666
rect 42254 45614 42306 45666
rect 44382 45614 44434 45666
rect 45614 45614 45666 45666
rect 52110 45614 52162 45666
rect 53790 45614 53842 45666
rect 54238 45614 54290 45666
rect 54798 45614 54850 45666
rect 55246 45614 55298 45666
rect 55806 45614 55858 45666
rect 56254 45614 56306 45666
rect 56590 45614 56642 45666
rect 57598 45614 57650 45666
rect 58046 45614 58098 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 2382 45278 2434 45330
rect 3278 45278 3330 45330
rect 8430 45278 8482 45330
rect 13022 45278 13074 45330
rect 13582 45278 13634 45330
rect 19182 45278 19234 45330
rect 19406 45278 19458 45330
rect 20302 45278 20354 45330
rect 23214 45278 23266 45330
rect 26574 45278 26626 45330
rect 30270 45278 30322 45330
rect 37214 45278 37266 45330
rect 42366 45278 42418 45330
rect 47518 45278 47570 45330
rect 52446 45278 52498 45330
rect 53230 45278 53282 45330
rect 2718 45166 2770 45218
rect 9774 45166 9826 45218
rect 12014 45166 12066 45218
rect 12574 45166 12626 45218
rect 13134 45166 13186 45218
rect 16718 45166 16770 45218
rect 22878 45166 22930 45218
rect 22990 45166 23042 45218
rect 25902 45166 25954 45218
rect 29710 45166 29762 45218
rect 36430 45166 36482 45218
rect 40686 45166 40738 45218
rect 43934 45166 43986 45218
rect 44606 45166 44658 45218
rect 45502 45166 45554 45218
rect 48078 45166 48130 45218
rect 54014 45166 54066 45218
rect 57486 45166 57538 45218
rect 57822 45166 57874 45218
rect 5406 45054 5458 45106
rect 5854 45054 5906 45106
rect 10110 45054 10162 45106
rect 12798 45054 12850 45106
rect 16270 45054 16322 45106
rect 18510 45054 18562 45106
rect 19070 45054 19122 45106
rect 19966 45054 20018 45106
rect 29934 45054 29986 45106
rect 30830 45054 30882 45106
rect 31726 45054 31778 45106
rect 32622 45054 32674 45106
rect 33742 45054 33794 45106
rect 34190 45054 34242 45106
rect 39566 45054 39618 45106
rect 40462 45054 40514 45106
rect 42702 45054 42754 45106
rect 43822 45054 43874 45106
rect 44494 45054 44546 45106
rect 45614 45054 45666 45106
rect 46286 45054 46338 45106
rect 46510 45054 46562 45106
rect 47966 45054 48018 45106
rect 48190 45054 48242 45106
rect 49534 45054 49586 45106
rect 50094 45054 50146 45106
rect 53790 45054 53842 45106
rect 54462 45054 54514 45106
rect 10894 44942 10946 44994
rect 11566 44942 11618 44994
rect 14030 44942 14082 44994
rect 15262 44942 15314 44994
rect 15934 44942 15986 44994
rect 17726 44942 17778 44994
rect 18062 44942 18114 44994
rect 20302 44942 20354 44994
rect 20862 44942 20914 44994
rect 26686 44942 26738 44994
rect 31054 44942 31106 44994
rect 32174 44942 32226 44994
rect 37662 44942 37714 44994
rect 38334 44942 38386 44994
rect 38894 44942 38946 44994
rect 41470 44942 41522 44994
rect 41918 44942 41970 44994
rect 45390 44942 45442 44994
rect 48750 44942 48802 44994
rect 55022 44942 55074 44994
rect 55582 44942 55634 44994
rect 55918 44942 55970 44994
rect 56366 44942 56418 44994
rect 8990 44830 9042 44882
rect 20190 44830 20242 44882
rect 25678 44830 25730 44882
rect 26014 44830 26066 44882
rect 31166 44830 31218 44882
rect 53678 44830 53730 44882
rect 54238 44830 54290 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 5966 44494 6018 44546
rect 24222 44494 24274 44546
rect 36318 44494 36370 44546
rect 42702 44494 42754 44546
rect 46174 44494 46226 44546
rect 47406 44494 47458 44546
rect 49646 44494 49698 44546
rect 49982 44494 50034 44546
rect 10446 44382 10498 44434
rect 20638 44382 20690 44434
rect 23214 44382 23266 44434
rect 25566 44382 25618 44434
rect 40238 44382 40290 44434
rect 41134 44382 41186 44434
rect 43934 44382 43986 44434
rect 47854 44382 47906 44434
rect 7870 44270 7922 44322
rect 8542 44270 8594 44322
rect 14254 44270 14306 44322
rect 14814 44270 14866 44322
rect 15038 44270 15090 44322
rect 15822 44270 15874 44322
rect 16046 44270 16098 44322
rect 16494 44270 16546 44322
rect 16942 44270 16994 44322
rect 17838 44270 17890 44322
rect 18174 44270 18226 44322
rect 19742 44270 19794 44322
rect 20414 44270 20466 44322
rect 22766 44270 22818 44322
rect 23102 44270 23154 44322
rect 23662 44270 23714 44322
rect 24334 44270 24386 44322
rect 24558 44270 24610 44322
rect 24670 44270 24722 44322
rect 26014 44270 26066 44322
rect 26462 44270 26514 44322
rect 29934 44270 29986 44322
rect 30382 44270 30434 44322
rect 35422 44270 35474 44322
rect 36430 44270 36482 44322
rect 42926 44270 42978 44322
rect 46062 44270 46114 44322
rect 46398 44270 46450 44322
rect 47182 44270 47234 44322
rect 47630 44270 47682 44322
rect 48638 44270 48690 44322
rect 48862 44270 48914 44322
rect 49086 44270 49138 44322
rect 50206 44270 50258 44322
rect 51326 44270 51378 44322
rect 6078 44158 6130 44210
rect 6638 44158 6690 44210
rect 7534 44158 7586 44210
rect 8766 44158 8818 44210
rect 9326 44158 9378 44210
rect 9662 44158 9714 44210
rect 10558 44158 10610 44210
rect 11118 44158 11170 44210
rect 15150 44158 15202 44210
rect 18398 44158 18450 44210
rect 29598 44158 29650 44210
rect 30942 44158 30994 44210
rect 31278 44158 31330 44210
rect 31502 44158 31554 44210
rect 32174 44158 32226 44210
rect 35086 44158 35138 44210
rect 36318 44158 36370 44210
rect 38894 44158 38946 44210
rect 39342 44158 39394 44210
rect 45838 44158 45890 44210
rect 48414 44158 48466 44210
rect 50878 44158 50930 44210
rect 5070 44046 5122 44098
rect 5966 44046 6018 44098
rect 6750 44046 6802 44098
rect 6862 44046 6914 44098
rect 10334 44046 10386 44098
rect 11454 44046 11506 44098
rect 12014 44046 12066 44098
rect 12910 44046 12962 44098
rect 15598 44046 15650 44098
rect 16270 44046 16322 44098
rect 16382 44046 16434 44098
rect 17278 44046 17330 44098
rect 18062 44046 18114 44098
rect 31166 44046 31218 44098
rect 32734 44046 32786 44098
rect 32846 44046 32898 44098
rect 32958 44046 33010 44098
rect 33182 44046 33234 44098
rect 37438 44046 37490 44098
rect 37998 44046 38050 44098
rect 38334 44046 38386 44098
rect 38782 44046 38834 44098
rect 39118 44046 39170 44098
rect 39902 44046 39954 44098
rect 40686 44046 40738 44098
rect 41694 44046 41746 44098
rect 42366 44046 42418 44098
rect 42590 44046 42642 44098
rect 43598 44046 43650 44098
rect 44494 44046 44546 44098
rect 46734 44046 46786 44098
rect 51998 44494 52050 44546
rect 54350 44494 54402 44546
rect 52222 44382 52274 44434
rect 55470 44382 55522 44434
rect 53454 44270 53506 44322
rect 53678 44270 53730 44322
rect 53902 44270 53954 44322
rect 55582 44270 55634 44322
rect 57486 44270 57538 44322
rect 55134 44158 55186 44210
rect 49646 44046 49698 44098
rect 50430 44046 50482 44098
rect 51550 44046 51602 44098
rect 51886 44046 51938 44098
rect 52670 44046 52722 44098
rect 56590 44046 56642 44098
rect 57150 44046 57202 44098
rect 57934 44046 57986 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 5742 43710 5794 43762
rect 6302 43710 6354 43762
rect 8206 43710 8258 43762
rect 8990 43710 9042 43762
rect 15934 43710 15986 43762
rect 16942 43710 16994 43762
rect 18062 43710 18114 43762
rect 19406 43710 19458 43762
rect 20974 43710 21026 43762
rect 25902 43710 25954 43762
rect 26126 43710 26178 43762
rect 34526 43710 34578 43762
rect 38782 43710 38834 43762
rect 39566 43710 39618 43762
rect 41918 43710 41970 43762
rect 46286 43710 46338 43762
rect 7086 43598 7138 43650
rect 7310 43598 7362 43650
rect 11790 43598 11842 43650
rect 13134 43598 13186 43650
rect 13582 43598 13634 43650
rect 14254 43598 14306 43650
rect 16830 43598 16882 43650
rect 18398 43598 18450 43650
rect 18510 43598 18562 43650
rect 22990 43598 23042 43650
rect 23214 43598 23266 43650
rect 25790 43598 25842 43650
rect 28478 43598 28530 43650
rect 32286 43598 32338 43650
rect 40238 43598 40290 43650
rect 40350 43598 40402 43650
rect 44718 43598 44770 43650
rect 45054 43598 45106 43650
rect 47294 43598 47346 43650
rect 47518 43598 47570 43650
rect 48078 43598 48130 43650
rect 49758 43598 49810 43650
rect 50318 43598 50370 43650
rect 51662 43598 51714 43650
rect 51998 43598 52050 43650
rect 54350 43598 54402 43650
rect 2830 43486 2882 43538
rect 3166 43486 3218 43538
rect 6974 43486 7026 43538
rect 8430 43486 8482 43538
rect 10222 43486 10274 43538
rect 10894 43486 10946 43538
rect 11118 43486 11170 43538
rect 11902 43486 11954 43538
rect 12574 43486 12626 43538
rect 15038 43486 15090 43538
rect 15486 43486 15538 43538
rect 16270 43486 16322 43538
rect 16606 43486 16658 43538
rect 18286 43486 18338 43538
rect 19070 43486 19122 43538
rect 20302 43486 20354 43538
rect 21422 43486 21474 43538
rect 23102 43486 23154 43538
rect 25678 43486 25730 43538
rect 29598 43486 29650 43538
rect 31278 43486 31330 43538
rect 31726 43486 31778 43538
rect 35870 43486 35922 43538
rect 36430 43486 36482 43538
rect 40014 43486 40066 43538
rect 40798 43486 40850 43538
rect 41694 43486 41746 43538
rect 42478 43486 42530 43538
rect 42814 43486 42866 43538
rect 44830 43486 44882 43538
rect 45278 43486 45330 43538
rect 45838 43486 45890 43538
rect 46174 43486 46226 43538
rect 46622 43486 46674 43538
rect 48526 43486 48578 43538
rect 49646 43486 49698 43538
rect 51326 43486 51378 43538
rect 53902 43486 53954 43538
rect 54126 43486 54178 43538
rect 56142 43486 56194 43538
rect 57374 43486 57426 43538
rect 7646 43374 7698 43426
rect 9662 43374 9714 43426
rect 22318 43374 22370 43426
rect 29038 43374 29090 43426
rect 32846 43374 32898 43426
rect 35086 43374 35138 43426
rect 35422 43374 35474 43426
rect 40238 43374 40290 43426
rect 43710 43374 43762 43426
rect 44942 43374 44994 43426
rect 47630 43374 47682 43426
rect 49422 43374 49474 43426
rect 52110 43374 52162 43426
rect 52782 43374 52834 43426
rect 53230 43374 53282 43426
rect 55358 43374 55410 43426
rect 56590 43374 56642 43426
rect 57934 43374 57986 43426
rect 12126 43262 12178 43314
rect 12350 43262 12402 43314
rect 14142 43262 14194 43314
rect 15262 43262 15314 43314
rect 20078 43262 20130 43314
rect 20638 43262 20690 43314
rect 20862 43262 20914 43314
rect 43150 43262 43202 43314
rect 46286 43262 46338 43314
rect 51102 43262 51154 43314
rect 52446 43262 52498 43314
rect 52670 43262 52722 43314
rect 54462 43262 54514 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 4958 42926 5010 42978
rect 6414 42926 6466 42978
rect 11342 42926 11394 42978
rect 11902 42926 11954 42978
rect 12462 42926 12514 42978
rect 20302 42926 20354 42978
rect 22990 42926 23042 42978
rect 29822 42926 29874 42978
rect 31054 42926 31106 42978
rect 38446 42926 38498 42978
rect 39454 42926 39506 42978
rect 40238 42926 40290 42978
rect 43486 42926 43538 42978
rect 45726 42926 45778 42978
rect 46286 42926 46338 42978
rect 47070 42926 47122 42978
rect 3054 42814 3106 42866
rect 5742 42814 5794 42866
rect 7198 42814 7250 42866
rect 12014 42814 12066 42866
rect 12462 42814 12514 42866
rect 13806 42814 13858 42866
rect 15374 42814 15426 42866
rect 18846 42814 18898 42866
rect 23326 42814 23378 42866
rect 24334 42814 24386 42866
rect 26350 42814 26402 42866
rect 28366 42814 28418 42866
rect 31950 42814 32002 42866
rect 33966 42814 34018 42866
rect 36094 42814 36146 42866
rect 36654 42814 36706 42866
rect 40014 42814 40066 42866
rect 41806 42814 41858 42866
rect 47070 42814 47122 42866
rect 47742 42926 47794 42978
rect 49310 42926 49362 42978
rect 54014 42926 54066 42978
rect 57150 42926 57202 42978
rect 57710 42926 57762 42978
rect 47854 42814 47906 42866
rect 48414 42814 48466 42866
rect 49310 42814 49362 42866
rect 50094 42814 50146 42866
rect 53342 42814 53394 42866
rect 57710 42814 57762 42866
rect 6302 42702 6354 42754
rect 7310 42702 7362 42754
rect 11006 42702 11058 42754
rect 11118 42702 11170 42754
rect 13582 42702 13634 42754
rect 15822 42702 15874 42754
rect 19518 42702 19570 42754
rect 20526 42702 20578 42754
rect 20750 42702 20802 42754
rect 22878 42702 22930 42754
rect 26910 42702 26962 42754
rect 28142 42702 28194 42754
rect 30382 42702 30434 42754
rect 30606 42702 30658 42754
rect 31502 42702 31554 42754
rect 31726 42702 31778 42754
rect 32510 42702 32562 42754
rect 32734 42702 32786 42754
rect 37662 42702 37714 42754
rect 37886 42702 37938 42754
rect 39678 42702 39730 42754
rect 40686 42702 40738 42754
rect 42814 42702 42866 42754
rect 43038 42702 43090 42754
rect 44270 42702 44322 42754
rect 45950 42702 46002 42754
rect 46510 42702 46562 42754
rect 50318 42702 50370 42754
rect 50878 42702 50930 42754
rect 51550 42702 51602 42754
rect 52558 42702 52610 42754
rect 54574 42702 54626 42754
rect 55022 42702 55074 42754
rect 55918 42702 55970 42754
rect 56254 42702 56306 42754
rect 2942 42590 2994 42642
rect 3278 42590 3330 42642
rect 3502 42590 3554 42642
rect 4846 42590 4898 42642
rect 6974 42590 7026 42642
rect 14142 42590 14194 42642
rect 15262 42590 15314 42642
rect 15598 42590 15650 42642
rect 20414 42590 20466 42642
rect 20862 42590 20914 42642
rect 24110 42590 24162 42642
rect 28814 42590 28866 42642
rect 30270 42590 30322 42642
rect 32622 42590 32674 42642
rect 35646 42590 35698 42642
rect 38222 42590 38274 42642
rect 40014 42590 40066 42642
rect 42926 42590 42978 42642
rect 44046 42590 44098 42642
rect 46062 42590 46114 42642
rect 50430 42590 50482 42642
rect 52222 42590 52274 42642
rect 54014 42590 54066 42642
rect 54126 42590 54178 42642
rect 55806 42590 55858 42642
rect 6750 42478 6802 42530
rect 7758 42478 7810 42530
rect 11006 42478 11058 42530
rect 13022 42478 13074 42530
rect 13918 42478 13970 42530
rect 14702 42478 14754 42530
rect 16270 42478 16322 42530
rect 17054 42478 17106 42530
rect 17614 42478 17666 42530
rect 18062 42478 18114 42530
rect 19742 42478 19794 42530
rect 24334 42478 24386 42530
rect 27246 42478 27298 42530
rect 32958 42478 33010 42530
rect 33518 42478 33570 42530
rect 34750 42478 34802 42530
rect 35422 42478 35474 42530
rect 35534 42478 35586 42530
rect 37550 42478 37602 42530
rect 41134 42478 41186 42530
rect 41246 42478 41298 42530
rect 41358 42478 41410 42530
rect 47518 42478 47570 42530
rect 48078 42478 48130 42530
rect 48974 42478 49026 42530
rect 55134 42478 55186 42530
rect 55246 42478 55298 42530
rect 57374 42478 57426 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 14030 42142 14082 42194
rect 15710 42142 15762 42194
rect 19966 42142 20018 42194
rect 20190 42142 20242 42194
rect 20750 42142 20802 42194
rect 21310 42142 21362 42194
rect 26014 42142 26066 42194
rect 35870 42142 35922 42194
rect 36094 42142 36146 42194
rect 36990 42142 37042 42194
rect 37998 42142 38050 42194
rect 38894 42142 38946 42194
rect 40238 42142 40290 42194
rect 45278 42142 45330 42194
rect 52110 42142 52162 42194
rect 52446 42142 52498 42194
rect 53118 42142 53170 42194
rect 56366 42142 56418 42194
rect 1822 42030 1874 42082
rect 3726 42030 3778 42082
rect 5518 42030 5570 42082
rect 6750 42030 6802 42082
rect 6974 42030 7026 42082
rect 12350 42030 12402 42082
rect 13918 42030 13970 42082
rect 16606 42030 16658 42082
rect 32398 42030 32450 42082
rect 34078 42030 34130 42082
rect 36766 42030 36818 42082
rect 37326 42030 37378 42082
rect 38110 42030 38162 42082
rect 39342 42030 39394 42082
rect 40462 42030 40514 42082
rect 44830 42030 44882 42082
rect 47630 42030 47682 42082
rect 55470 42030 55522 42082
rect 56142 42030 56194 42082
rect 2494 41918 2546 41970
rect 5406 41918 5458 41970
rect 5742 41918 5794 41970
rect 5966 41918 6018 41970
rect 6414 41918 6466 41970
rect 9774 41918 9826 41970
rect 9998 41918 10050 41970
rect 12910 41918 12962 41970
rect 14254 41918 14306 41970
rect 14478 41918 14530 41970
rect 16718 41918 16770 41970
rect 18062 41918 18114 41970
rect 18958 41918 19010 41970
rect 19854 41918 19906 41970
rect 20638 41918 20690 41970
rect 25790 41918 25842 41970
rect 26014 41918 26066 41970
rect 26350 41918 26402 41970
rect 26686 41918 26738 41970
rect 31838 41918 31890 41970
rect 33630 41918 33682 41970
rect 34750 41918 34802 41970
rect 35646 41918 35698 41970
rect 37102 41918 37154 41970
rect 37774 41918 37826 41970
rect 38670 41918 38722 41970
rect 39118 41918 39170 41970
rect 39902 41918 39954 41970
rect 40126 41918 40178 41970
rect 41806 41918 41858 41970
rect 42030 41918 42082 41970
rect 43822 41918 43874 41970
rect 45950 41918 46002 41970
rect 46622 41918 46674 41970
rect 46846 41918 46898 41970
rect 48190 41918 48242 41970
rect 48526 41918 48578 41970
rect 50206 41918 50258 41970
rect 50430 41918 50482 41970
rect 51102 41918 51154 41970
rect 55246 41918 55298 41970
rect 56702 41918 56754 41970
rect 3838 41806 3890 41858
rect 6862 41806 6914 41858
rect 8766 41806 8818 41858
rect 10782 41806 10834 41858
rect 11342 41806 11394 41858
rect 13134 41806 13186 41858
rect 14926 41806 14978 41858
rect 17726 41806 17778 41858
rect 18622 41806 18674 41858
rect 31614 41806 31666 41858
rect 34974 41806 35026 41858
rect 35758 41806 35810 41858
rect 47742 41806 47794 41858
rect 49870 41806 49922 41858
rect 51550 41806 51602 41858
rect 53678 41806 53730 41858
rect 54126 41806 54178 41858
rect 54574 41806 54626 41858
rect 55582 41806 55634 41858
rect 56254 41806 56306 41858
rect 57374 41806 57426 41858
rect 57822 41806 57874 41858
rect 10110 41694 10162 41746
rect 16046 41694 16098 41746
rect 17726 41694 17778 41746
rect 18622 41694 18674 41746
rect 20750 41694 20802 41746
rect 39230 41694 39282 41746
rect 46398 41694 46450 41746
rect 54126 41694 54178 41746
rect 55022 41694 55074 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 3950 41358 4002 41410
rect 7870 41358 7922 41410
rect 8990 41358 9042 41410
rect 13918 41358 13970 41410
rect 14254 41358 14306 41410
rect 16158 41358 16210 41410
rect 23102 41358 23154 41410
rect 27246 41358 27298 41410
rect 49310 41358 49362 41410
rect 51326 41358 51378 41410
rect 51550 41358 51602 41410
rect 3726 41246 3778 41298
rect 10446 41246 10498 41298
rect 13694 41246 13746 41298
rect 17838 41246 17890 41298
rect 18286 41246 18338 41298
rect 26350 41246 26402 41298
rect 35646 41246 35698 41298
rect 37886 41246 37938 41298
rect 39118 41246 39170 41298
rect 40574 41246 40626 41298
rect 41022 41246 41074 41298
rect 42142 41246 42194 41298
rect 51326 41246 51378 41298
rect 2606 41134 2658 41186
rect 2942 41134 2994 41186
rect 6526 41134 6578 41186
rect 8542 41134 8594 41186
rect 9438 41134 9490 41186
rect 10222 41134 10274 41186
rect 10782 41134 10834 41186
rect 15822 41134 15874 41186
rect 16494 41134 16546 41186
rect 17614 41134 17666 41186
rect 19294 41134 19346 41186
rect 21870 41134 21922 41186
rect 25006 41134 25058 41186
rect 27806 41134 27858 41186
rect 28590 41134 28642 41186
rect 29598 41134 29650 41186
rect 34190 41134 34242 41186
rect 34302 41134 34354 41186
rect 35422 41134 35474 41186
rect 36318 41134 36370 41186
rect 38670 41134 38722 41186
rect 38894 41134 38946 41186
rect 42254 41134 42306 41186
rect 42702 41134 42754 41186
rect 43598 41134 43650 41186
rect 46510 41134 46562 41186
rect 54126 41134 54178 41186
rect 55246 41134 55298 41186
rect 56590 41134 56642 41186
rect 3054 41022 3106 41074
rect 3726 41022 3778 41074
rect 5742 41022 5794 41074
rect 6190 41022 6242 41074
rect 6302 41022 6354 41074
rect 8206 41022 8258 41074
rect 9550 41022 9602 41074
rect 9662 41022 9714 41074
rect 10670 41022 10722 41074
rect 21646 41022 21698 41074
rect 22766 41022 22818 41074
rect 25902 41022 25954 41074
rect 27358 41022 27410 41074
rect 28702 41022 28754 41074
rect 29934 41022 29986 41074
rect 30158 41022 30210 41074
rect 31502 41022 31554 41074
rect 31726 41022 31778 41074
rect 31838 41022 31890 41074
rect 33854 41022 33906 41074
rect 35646 41022 35698 41074
rect 36094 41022 36146 41074
rect 39118 41022 39170 41074
rect 39678 41022 39730 41074
rect 40014 41022 40066 41074
rect 44382 41022 44434 41074
rect 45390 41022 45442 41074
rect 46286 41022 46338 41074
rect 46846 41022 46898 41074
rect 47742 41022 47794 41074
rect 48974 41022 49026 41074
rect 49198 41022 49250 41074
rect 53790 41022 53842 41074
rect 56254 41022 56306 41074
rect 7310 40910 7362 40962
rect 7982 40910 8034 40962
rect 11678 40910 11730 40962
rect 12574 40910 12626 40962
rect 13022 40910 13074 40962
rect 15150 40910 15202 40962
rect 18846 40910 18898 40962
rect 19630 40910 19682 40962
rect 20190 40910 20242 40962
rect 20862 40910 20914 40962
rect 22206 40910 22258 40962
rect 22990 40910 23042 40962
rect 24670 40910 24722 40962
rect 27246 40910 27298 40962
rect 28926 40910 28978 40962
rect 29822 40910 29874 40962
rect 34078 40910 34130 40962
rect 37550 40910 37602 40962
rect 41582 40910 41634 40962
rect 43822 40910 43874 40962
rect 44718 40910 44770 40962
rect 46398 40910 46450 40962
rect 48078 40910 48130 40962
rect 49758 40910 49810 40962
rect 50206 40910 50258 40962
rect 50654 40910 50706 40962
rect 51774 40910 51826 40962
rect 52222 40910 52274 40962
rect 52782 40910 52834 40962
rect 55358 40910 55410 40962
rect 56366 40910 56418 40962
rect 57038 40910 57090 40962
rect 57374 40910 57426 40962
rect 57822 40910 57874 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 4958 40574 5010 40626
rect 6302 40574 6354 40626
rect 6750 40574 6802 40626
rect 9886 40574 9938 40626
rect 9998 40574 10050 40626
rect 13246 40574 13298 40626
rect 19518 40574 19570 40626
rect 20638 40574 20690 40626
rect 25790 40574 25842 40626
rect 34750 40574 34802 40626
rect 36206 40574 36258 40626
rect 36318 40574 36370 40626
rect 36430 40574 36482 40626
rect 36878 40574 36930 40626
rect 39118 40574 39170 40626
rect 39566 40574 39618 40626
rect 40462 40574 40514 40626
rect 41694 40574 41746 40626
rect 43038 40574 43090 40626
rect 43262 40574 43314 40626
rect 44606 40574 44658 40626
rect 44718 40574 44770 40626
rect 45166 40574 45218 40626
rect 45614 40574 45666 40626
rect 48526 40574 48578 40626
rect 48638 40574 48690 40626
rect 48750 40574 48802 40626
rect 51214 40574 51266 40626
rect 51886 40574 51938 40626
rect 54350 40574 54402 40626
rect 7534 40462 7586 40514
rect 7646 40462 7698 40514
rect 10222 40462 10274 40514
rect 14478 40462 14530 40514
rect 16382 40462 16434 40514
rect 19406 40462 19458 40514
rect 20526 40462 20578 40514
rect 21646 40462 21698 40514
rect 23886 40462 23938 40514
rect 26798 40462 26850 40514
rect 33742 40462 33794 40514
rect 33854 40462 33906 40514
rect 38222 40462 38274 40514
rect 41918 40462 41970 40514
rect 42142 40462 42194 40514
rect 44494 40462 44546 40514
rect 46958 40462 47010 40514
rect 48302 40462 48354 40514
rect 49534 40462 49586 40514
rect 49870 40462 49922 40514
rect 52334 40462 52386 40514
rect 52558 40462 52610 40514
rect 55134 40462 55186 40514
rect 2830 40350 2882 40402
rect 8094 40350 8146 40402
rect 9774 40350 9826 40402
rect 11566 40350 11618 40402
rect 12126 40350 12178 40402
rect 15374 40350 15426 40402
rect 16046 40350 16098 40402
rect 16942 40350 16994 40402
rect 17726 40350 17778 40402
rect 18734 40350 18786 40402
rect 19294 40350 19346 40402
rect 19742 40350 19794 40402
rect 20302 40350 20354 40402
rect 20974 40350 21026 40402
rect 21534 40350 21586 40402
rect 23326 40350 23378 40402
rect 24334 40350 24386 40402
rect 27470 40350 27522 40402
rect 28366 40350 28418 40402
rect 28926 40350 28978 40402
rect 30046 40350 30098 40402
rect 30494 40350 30546 40402
rect 31390 40350 31442 40402
rect 33518 40350 33570 40402
rect 35310 40350 35362 40402
rect 35758 40350 35810 40402
rect 37998 40350 38050 40402
rect 38334 40350 38386 40402
rect 38670 40350 38722 40402
rect 41582 40350 41634 40402
rect 42702 40350 42754 40402
rect 44046 40350 44098 40402
rect 44270 40350 44322 40402
rect 46622 40350 46674 40402
rect 47406 40350 47458 40402
rect 50766 40350 50818 40402
rect 1934 40238 1986 40290
rect 5406 40238 5458 40290
rect 5854 40238 5906 40290
rect 7870 40238 7922 40290
rect 9102 40238 9154 40290
rect 11118 40238 11170 40290
rect 14142 40238 14194 40290
rect 18286 40238 18338 40290
rect 22206 40238 22258 40290
rect 22654 40238 22706 40290
rect 24670 40238 24722 40290
rect 25678 40238 25730 40290
rect 27694 40238 27746 40290
rect 29150 40238 29202 40290
rect 31166 40238 31218 40290
rect 37326 40238 37378 40290
rect 40014 40238 40066 40290
rect 42926 40238 42978 40290
rect 46846 40238 46898 40290
rect 50430 40238 50482 40290
rect 52446 40294 52498 40346
rect 53230 40350 53282 40402
rect 54126 40350 54178 40402
rect 55022 40350 55074 40402
rect 55806 40350 55858 40402
rect 56142 40350 56194 40402
rect 56702 40238 56754 40290
rect 57374 40238 57426 40290
rect 57934 40238 57986 40290
rect 5518 40126 5570 40178
rect 6190 40126 6242 40178
rect 7310 40126 7362 40178
rect 12350 40126 12402 40178
rect 12574 40126 12626 40178
rect 12798 40126 12850 40178
rect 13806 40126 13858 40178
rect 13918 40126 13970 40178
rect 14366 40126 14418 40178
rect 17614 40126 17666 40178
rect 18286 40126 18338 40178
rect 21646 40126 21698 40178
rect 26014 40126 26066 40178
rect 35086 40126 35138 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 6862 39790 6914 39842
rect 8430 39790 8482 39842
rect 8654 39790 8706 39842
rect 9102 39790 9154 39842
rect 19630 39790 19682 39842
rect 29598 39790 29650 39842
rect 35646 39790 35698 39842
rect 44046 39790 44098 39842
rect 44606 39790 44658 39842
rect 52782 39790 52834 39842
rect 56814 39790 56866 39842
rect 3166 39678 3218 39730
rect 5742 39678 5794 39730
rect 7310 39678 7362 39730
rect 7758 39678 7810 39730
rect 8206 39678 8258 39730
rect 13918 39678 13970 39730
rect 22094 39678 22146 39730
rect 22766 39678 22818 39730
rect 31726 39678 31778 39730
rect 33518 39678 33570 39730
rect 36206 39678 36258 39730
rect 38670 39678 38722 39730
rect 39342 39678 39394 39730
rect 41694 39678 41746 39730
rect 43262 39678 43314 39730
rect 46174 39678 46226 39730
rect 54238 39678 54290 39730
rect 2718 39566 2770 39618
rect 4174 39566 4226 39618
rect 4398 39566 4450 39618
rect 4734 39566 4786 39618
rect 5966 39566 6018 39618
rect 6190 39566 6242 39618
rect 6414 39566 6466 39618
rect 13806 39566 13858 39618
rect 14142 39566 14194 39618
rect 14478 39566 14530 39618
rect 17838 39566 17890 39618
rect 19966 39566 20018 39618
rect 21646 39566 21698 39618
rect 31166 39566 31218 39618
rect 32286 39566 32338 39618
rect 33630 39566 33682 39618
rect 35758 39566 35810 39618
rect 38110 39566 38162 39618
rect 39006 39566 39058 39618
rect 42590 39566 42642 39618
rect 43374 39566 43426 39618
rect 46062 39566 46114 39618
rect 46398 39566 46450 39618
rect 46510 39566 46562 39618
rect 46734 39566 46786 39618
rect 47742 39566 47794 39618
rect 49086 39566 49138 39618
rect 49646 39566 49698 39618
rect 55246 39566 55298 39618
rect 55694 39566 55746 39618
rect 55918 39566 55970 39618
rect 56366 39566 56418 39618
rect 57038 39566 57090 39618
rect 57262 39566 57314 39618
rect 57710 39566 57762 39618
rect 2382 39454 2434 39506
rect 4958 39454 5010 39506
rect 10334 39454 10386 39506
rect 10670 39454 10722 39506
rect 20190 39454 20242 39506
rect 20526 39454 20578 39506
rect 29822 39454 29874 39506
rect 31614 39454 31666 39506
rect 32846 39454 32898 39506
rect 36654 39454 36706 39506
rect 37774 39454 37826 39506
rect 43038 39454 43090 39506
rect 43150 39454 43202 39506
rect 44046 39454 44098 39506
rect 48078 39454 48130 39506
rect 54910 39454 54962 39506
rect 55806 39454 55858 39506
rect 4062 39342 4114 39394
rect 9886 39342 9938 39394
rect 11118 39342 11170 39394
rect 11678 39342 11730 39394
rect 12126 39342 12178 39394
rect 12574 39342 12626 39394
rect 13022 39342 13074 39394
rect 14030 39342 14082 39394
rect 15038 39342 15090 39394
rect 15598 39342 15650 39394
rect 16046 39342 16098 39394
rect 16830 39342 16882 39394
rect 17278 39342 17330 39394
rect 18062 39342 18114 39394
rect 18622 39342 18674 39394
rect 19070 39342 19122 39394
rect 21982 39342 22034 39394
rect 22206 39342 22258 39394
rect 23214 39342 23266 39394
rect 24782 39342 24834 39394
rect 25342 39342 25394 39394
rect 25790 39342 25842 39394
rect 29710 39342 29762 39394
rect 30606 39342 30658 39394
rect 35646 39342 35698 39394
rect 37886 39342 37938 39394
rect 39902 39342 39954 39394
rect 40350 39342 40402 39394
rect 40798 39342 40850 39394
rect 41246 39342 41298 39394
rect 42142 39342 42194 39394
rect 44494 39342 44546 39394
rect 45502 39342 45554 39394
rect 48526 39342 48578 39394
rect 52110 39342 52162 39394
rect 53454 39342 53506 39394
rect 53790 39342 53842 39394
rect 55022 39342 55074 39394
rect 57486 39342 57538 39394
rect 57598 39342 57650 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 3726 39006 3778 39058
rect 5518 39006 5570 39058
rect 6190 39006 6242 39058
rect 7646 39006 7698 39058
rect 8206 39006 8258 39058
rect 11566 39006 11618 39058
rect 14478 39006 14530 39058
rect 21086 39006 21138 39058
rect 22542 39006 22594 39058
rect 33630 39006 33682 39058
rect 37102 39006 37154 39058
rect 39566 39006 39618 39058
rect 40574 39006 40626 39058
rect 41806 39006 41858 39058
rect 46062 39006 46114 39058
rect 47518 39006 47570 39058
rect 48302 39006 48354 39058
rect 48526 39006 48578 39058
rect 50990 39006 51042 39058
rect 51438 39006 51490 39058
rect 52334 39006 52386 39058
rect 54574 39006 54626 39058
rect 56590 39006 56642 39058
rect 57374 39006 57426 39058
rect 8990 38894 9042 38946
rect 12462 38894 12514 38946
rect 15598 38894 15650 38946
rect 16830 38894 16882 38946
rect 16942 38894 16994 38946
rect 18062 38894 18114 38946
rect 20414 38894 20466 38946
rect 20862 38894 20914 38946
rect 21758 38894 21810 38946
rect 22990 38894 23042 38946
rect 24334 38894 24386 38946
rect 25790 38894 25842 38946
rect 28814 38894 28866 38946
rect 30270 38894 30322 38946
rect 34078 38894 34130 38946
rect 34302 38894 34354 38946
rect 38446 38894 38498 38946
rect 42030 38894 42082 38946
rect 43150 38894 43202 38946
rect 44606 38894 44658 38946
rect 46510 38894 46562 38946
rect 47630 38894 47682 38946
rect 51998 38894 52050 38946
rect 54350 38894 54402 38946
rect 4174 38782 4226 38834
rect 4622 38782 4674 38834
rect 4734 38782 4786 38834
rect 5406 38782 5458 38834
rect 7086 38782 7138 38834
rect 7422 38782 7474 38834
rect 8654 38782 8706 38834
rect 10782 38782 10834 38834
rect 10894 38782 10946 38834
rect 11342 38782 11394 38834
rect 13022 38782 13074 38834
rect 14030 38782 14082 38834
rect 14254 38782 14306 38834
rect 14926 38782 14978 38834
rect 15486 38782 15538 38834
rect 15822 38782 15874 38834
rect 16606 38782 16658 38834
rect 17726 38782 17778 38834
rect 17950 38782 18002 38834
rect 19182 38782 19234 38834
rect 21982 38782 22034 38834
rect 22542 38782 22594 38834
rect 24446 38782 24498 38834
rect 25902 38782 25954 38834
rect 26910 38782 26962 38834
rect 29822 38782 29874 38834
rect 30382 38782 30434 38834
rect 34190 38782 34242 38834
rect 35534 38782 35586 38834
rect 36094 38782 36146 38834
rect 36318 38782 36370 38834
rect 36766 38782 36818 38834
rect 37998 38782 38050 38834
rect 38222 38782 38274 38834
rect 39006 38782 39058 38834
rect 41582 38782 41634 38834
rect 42478 38782 42530 38834
rect 44158 38782 44210 38834
rect 44942 38782 44994 38834
rect 48190 38782 48242 38834
rect 49870 38782 49922 38834
rect 50542 38782 50594 38834
rect 53678 38782 53730 38834
rect 54126 38782 54178 38834
rect 6750 38670 6802 38722
rect 9998 38670 10050 38722
rect 10558 38670 10610 38722
rect 12126 38670 12178 38722
rect 13470 38670 13522 38722
rect 13918 38670 13970 38722
rect 16158 38670 16210 38722
rect 19854 38670 19906 38722
rect 22206 38670 22258 38722
rect 23662 38670 23714 38722
rect 25006 38670 25058 38722
rect 26014 38670 26066 38722
rect 27022 38670 27074 38722
rect 27806 38670 27858 38722
rect 28254 38670 28306 38722
rect 36206 38670 36258 38722
rect 38334 38670 38386 38722
rect 39230 38670 39282 38722
rect 40126 38670 40178 38722
rect 41918 38670 41970 38722
rect 45502 38670 45554 38722
rect 47070 38670 47122 38722
rect 50094 38670 50146 38722
rect 5182 38558 5234 38610
rect 6190 38558 6242 38610
rect 6638 38558 6690 38610
rect 7758 38558 7810 38610
rect 12574 38558 12626 38610
rect 12798 38558 12850 38610
rect 14814 38558 14866 38610
rect 18286 38558 18338 38610
rect 18510 38558 18562 38610
rect 21198 38558 21250 38610
rect 24334 38558 24386 38610
rect 29038 38558 29090 38610
rect 43598 38558 43650 38610
rect 45726 38558 45778 38610
rect 57598 39006 57650 39058
rect 55246 38894 55298 38946
rect 57710 38894 57762 38946
rect 56030 38782 56082 38834
rect 54910 38670 54962 38722
rect 55022 38558 55074 38610
rect 56254 38558 56306 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 5070 38222 5122 38274
rect 18510 38222 18562 38274
rect 25230 38222 25282 38274
rect 36766 38222 36818 38274
rect 40798 38222 40850 38274
rect 42030 38222 42082 38274
rect 52782 38222 52834 38274
rect 56142 38222 56194 38274
rect 57262 38222 57314 38274
rect 5630 38110 5682 38162
rect 7422 38110 7474 38162
rect 8206 38110 8258 38162
rect 8766 38110 8818 38162
rect 10222 38110 10274 38162
rect 11006 38110 11058 38162
rect 14478 38110 14530 38162
rect 14590 38110 14642 38162
rect 17390 38110 17442 38162
rect 20862 38110 20914 38162
rect 23214 38110 23266 38162
rect 30046 38110 30098 38162
rect 30718 38110 30770 38162
rect 33966 38110 34018 38162
rect 34862 38110 34914 38162
rect 36542 38110 36594 38162
rect 40574 38110 40626 38162
rect 43374 38110 43426 38162
rect 50206 38110 50258 38162
rect 53342 38110 53394 38162
rect 55806 38110 55858 38162
rect 57822 38110 57874 38162
rect 3614 37998 3666 38050
rect 4174 37998 4226 38050
rect 4622 37998 4674 38050
rect 5742 37998 5794 38050
rect 6302 37998 6354 38050
rect 7758 37998 7810 38050
rect 9662 37998 9714 38050
rect 11454 37998 11506 38050
rect 12238 37998 12290 38050
rect 12686 37998 12738 38050
rect 12910 37998 12962 38050
rect 14030 37998 14082 38050
rect 14814 37998 14866 38050
rect 17614 37998 17666 38050
rect 19518 37998 19570 38050
rect 19742 37998 19794 38050
rect 22206 37998 22258 38050
rect 23998 37998 24050 38050
rect 25454 37998 25506 38050
rect 25902 37998 25954 38050
rect 27806 37998 27858 38050
rect 28366 37998 28418 38050
rect 30158 37998 30210 38050
rect 33518 37998 33570 38050
rect 34078 37998 34130 38050
rect 35982 37998 36034 38050
rect 36206 37998 36258 38050
rect 37438 37998 37490 38050
rect 37774 37998 37826 38050
rect 39342 37998 39394 38050
rect 40462 37998 40514 38050
rect 41694 37998 41746 38050
rect 45838 37998 45890 38050
rect 51886 37998 51938 38050
rect 52110 37998 52162 38050
rect 52334 37998 52386 38050
rect 54910 37998 54962 38050
rect 56030 37998 56082 38050
rect 57598 37998 57650 38050
rect 4286 37886 4338 37938
rect 4398 37886 4450 37938
rect 5966 37886 6018 37938
rect 11006 37886 11058 37938
rect 11230 37886 11282 37938
rect 15038 37886 15090 37938
rect 16046 37886 16098 37938
rect 16158 37886 16210 37938
rect 16270 37886 16322 37938
rect 18846 37886 18898 37938
rect 20078 37886 20130 37938
rect 22430 37886 22482 37938
rect 24334 37886 24386 37938
rect 27694 37886 27746 37938
rect 31054 37886 31106 37938
rect 31838 37886 31890 37938
rect 34862 37886 34914 37938
rect 35310 37886 35362 37938
rect 36542 37886 36594 37938
rect 37662 37886 37714 37938
rect 39006 37886 39058 37938
rect 41470 37886 41522 37938
rect 43150 37886 43202 37938
rect 43262 37886 43314 37938
rect 44046 37886 44098 37938
rect 45502 37886 45554 37938
rect 48750 37886 48802 37938
rect 55022 37886 55074 37938
rect 6190 37774 6242 37826
rect 9102 37774 9154 37826
rect 10894 37774 10946 37826
rect 12350 37774 12402 37826
rect 12462 37774 12514 37826
rect 15822 37774 15874 37826
rect 15934 37774 15986 37826
rect 17950 37774 18002 37826
rect 18622 37774 18674 37826
rect 19630 37774 19682 37826
rect 21534 37774 21586 37826
rect 29710 37774 29762 37826
rect 29934 37774 29986 37826
rect 30830 37774 30882 37826
rect 31502 37774 31554 37826
rect 31726 37774 31778 37826
rect 32398 37774 32450 37826
rect 32734 37774 32786 37826
rect 33854 37774 33906 37826
rect 35086 37774 35138 37826
rect 38446 37774 38498 37826
rect 43374 37774 43426 37826
rect 43598 37774 43650 37826
rect 44494 37774 44546 37826
rect 45614 37774 45666 37826
rect 46174 37774 46226 37826
rect 46622 37774 46674 37826
rect 47182 37774 47234 37826
rect 47966 37774 48018 37826
rect 48302 37774 48354 37826
rect 49422 37774 49474 37826
rect 49758 37774 49810 37826
rect 50654 37774 50706 37826
rect 51214 37774 51266 37826
rect 53790 37774 53842 37826
rect 54798 37774 54850 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 4062 37438 4114 37490
rect 4734 37438 4786 37490
rect 4846 37438 4898 37490
rect 4958 37438 5010 37490
rect 6862 37438 6914 37490
rect 7086 37438 7138 37490
rect 8094 37438 8146 37490
rect 10558 37438 10610 37490
rect 12238 37438 12290 37490
rect 13918 37438 13970 37490
rect 20638 37438 20690 37490
rect 25566 37438 25618 37490
rect 26350 37438 26402 37490
rect 27358 37438 27410 37490
rect 27470 37438 27522 37490
rect 32958 37438 33010 37490
rect 35310 37438 35362 37490
rect 36878 37438 36930 37490
rect 36990 37438 37042 37490
rect 38334 37438 38386 37490
rect 39566 37438 39618 37490
rect 44158 37438 44210 37490
rect 47406 37438 47458 37490
rect 52670 37438 52722 37490
rect 11454 37326 11506 37378
rect 13806 37326 13858 37378
rect 14590 37326 14642 37378
rect 16718 37326 16770 37378
rect 19854 37326 19906 37378
rect 20862 37326 20914 37378
rect 22654 37326 22706 37378
rect 24110 37326 24162 37378
rect 25790 37326 25842 37378
rect 25902 37326 25954 37378
rect 27582 37326 27634 37378
rect 28030 37326 28082 37378
rect 28814 37326 28866 37378
rect 32622 37326 32674 37378
rect 32734 37326 32786 37378
rect 39902 37326 39954 37378
rect 41694 37326 41746 37378
rect 46398 37326 46450 37378
rect 48302 37326 48354 37378
rect 50206 37326 50258 37378
rect 53566 37326 53618 37378
rect 57374 37326 57426 37378
rect 4510 37214 4562 37266
rect 5182 37214 5234 37266
rect 6862 37214 6914 37266
rect 7310 37214 7362 37266
rect 7422 37214 7474 37266
rect 11902 37214 11954 37266
rect 13358 37214 13410 37266
rect 13582 37214 13634 37266
rect 14366 37214 14418 37266
rect 14926 37214 14978 37266
rect 15598 37214 15650 37266
rect 18398 37214 18450 37266
rect 19070 37214 19122 37266
rect 19966 37214 20018 37266
rect 20638 37214 20690 37266
rect 21534 37214 21586 37266
rect 23438 37214 23490 37266
rect 23886 37214 23938 37266
rect 24670 37214 24722 37266
rect 29710 37214 29762 37266
rect 31838 37214 31890 37266
rect 33630 37214 33682 37266
rect 33742 37214 33794 37266
rect 34078 37214 34130 37266
rect 36206 37214 36258 37266
rect 36766 37214 36818 37266
rect 37438 37214 37490 37266
rect 41806 37214 41858 37266
rect 41918 37214 41970 37266
rect 42814 37214 42866 37266
rect 43934 37214 43986 37266
rect 44158 37214 44210 37266
rect 44494 37214 44546 37266
rect 46734 37214 46786 37266
rect 48414 37214 48466 37266
rect 50430 37214 50482 37266
rect 50766 37214 50818 37266
rect 52782 37214 52834 37266
rect 53006 37214 53058 37266
rect 56366 37214 56418 37266
rect 5630 37102 5682 37154
rect 6302 37102 6354 37154
rect 11006 37102 11058 37154
rect 12910 37102 12962 37154
rect 14254 37102 14306 37154
rect 16606 37102 16658 37154
rect 17726 37102 17778 37154
rect 18174 37102 18226 37154
rect 24558 37102 24610 37154
rect 29486 37102 29538 37154
rect 31054 37102 31106 37154
rect 31166 37102 31218 37154
rect 37998 37102 38050 37154
rect 38782 37102 38834 37154
rect 40350 37102 40402 37154
rect 40798 37102 40850 37154
rect 43262 37102 43314 37154
rect 44942 37102 44994 37154
rect 45502 37102 45554 37154
rect 45950 37102 46002 37154
rect 49534 37102 49586 37154
rect 50318 37102 50370 37154
rect 51214 37102 51266 37154
rect 55694 37102 55746 37154
rect 57822 37102 57874 37154
rect 16942 36990 16994 37042
rect 18622 36990 18674 37042
rect 35758 36990 35810 37042
rect 35982 36990 36034 37042
rect 37662 36990 37714 37042
rect 38446 36990 38498 37042
rect 42366 36990 42418 37042
rect 42590 36990 42642 37042
rect 43598 36990 43650 37042
rect 47742 36990 47794 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 7422 36654 7474 36706
rect 7646 36654 7698 36706
rect 38670 36654 38722 36706
rect 45502 36654 45554 36706
rect 54350 36654 54402 36706
rect 55246 36654 55298 36706
rect 7870 36542 7922 36594
rect 8766 36542 8818 36594
rect 9550 36542 9602 36594
rect 13918 36542 13970 36594
rect 15598 36542 15650 36594
rect 16270 36542 16322 36594
rect 18734 36542 18786 36594
rect 24334 36542 24386 36594
rect 33182 36542 33234 36594
rect 37438 36542 37490 36594
rect 47966 36542 48018 36594
rect 52222 36542 52274 36594
rect 56142 36542 56194 36594
rect 8318 36430 8370 36482
rect 9774 36430 9826 36482
rect 14814 36430 14866 36482
rect 15150 36430 15202 36482
rect 16718 36430 16770 36482
rect 19854 36430 19906 36482
rect 20190 36430 20242 36482
rect 27134 36430 27186 36482
rect 32286 36430 32338 36482
rect 32734 36430 32786 36482
rect 33630 36430 33682 36482
rect 39678 36430 39730 36482
rect 45838 36430 45890 36482
rect 48078 36430 48130 36482
rect 49646 36430 49698 36482
rect 51214 36430 51266 36482
rect 52110 36430 52162 36482
rect 52670 36430 52722 36482
rect 53902 36430 53954 36482
rect 54238 36430 54290 36482
rect 57262 36430 57314 36482
rect 57710 36430 57762 36482
rect 9438 36318 9490 36370
rect 14366 36318 14418 36370
rect 14590 36318 14642 36370
rect 17278 36318 17330 36370
rect 20414 36318 20466 36370
rect 21646 36318 21698 36370
rect 21982 36318 22034 36370
rect 24558 36318 24610 36370
rect 24782 36318 24834 36370
rect 24894 36318 24946 36370
rect 37998 36318 38050 36370
rect 38782 36318 38834 36370
rect 40574 36318 40626 36370
rect 43038 36318 43090 36370
rect 43262 36318 43314 36370
rect 43822 36318 43874 36370
rect 44158 36318 44210 36370
rect 46062 36318 46114 36370
rect 47294 36318 47346 36370
rect 48190 36318 48242 36370
rect 52446 36318 52498 36370
rect 53454 36318 53506 36370
rect 53678 36318 53730 36370
rect 56814 36318 56866 36370
rect 5070 36206 5122 36258
rect 6078 36206 6130 36258
rect 6526 36206 6578 36258
rect 6974 36206 7026 36258
rect 7310 36206 7362 36258
rect 10222 36206 10274 36258
rect 11006 36206 11058 36258
rect 12014 36206 12066 36258
rect 12462 36206 12514 36258
rect 12910 36206 12962 36258
rect 14702 36206 14754 36258
rect 17166 36206 17218 36258
rect 17726 36206 17778 36258
rect 18174 36206 18226 36258
rect 19182 36206 19234 36258
rect 20078 36206 20130 36258
rect 23774 36206 23826 36258
rect 25118 36206 25170 36258
rect 25678 36206 25730 36258
rect 26014 36206 26066 36258
rect 26798 36206 26850 36258
rect 31278 36206 31330 36258
rect 36430 36206 36482 36258
rect 38670 36206 38722 36258
rect 39342 36206 39394 36258
rect 40238 36206 40290 36258
rect 41022 36206 41074 36258
rect 41582 36206 41634 36258
rect 41918 36206 41970 36258
rect 42478 36206 42530 36258
rect 43150 36206 43202 36258
rect 44606 36206 44658 36258
rect 46734 36206 46786 36258
rect 53790 36206 53842 36258
rect 54798 36206 54850 36258
rect 55134 36206 55186 36258
rect 55582 36206 55634 36258
rect 56254 36206 56306 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 7086 35870 7138 35922
rect 7198 35870 7250 35922
rect 8318 35870 8370 35922
rect 8654 35870 8706 35922
rect 9998 35870 10050 35922
rect 13134 35870 13186 35922
rect 14142 35870 14194 35922
rect 16606 35870 16658 35922
rect 16942 35870 16994 35922
rect 17726 35870 17778 35922
rect 30494 35870 30546 35922
rect 31838 35870 31890 35922
rect 32398 35870 32450 35922
rect 35646 35870 35698 35922
rect 36990 35870 37042 35922
rect 38558 35870 38610 35922
rect 45726 35870 45778 35922
rect 46286 35870 46338 35922
rect 48302 35870 48354 35922
rect 51102 35870 51154 35922
rect 51662 35870 51714 35922
rect 52670 35870 52722 35922
rect 57822 35870 57874 35922
rect 4398 35758 4450 35810
rect 8878 35758 8930 35810
rect 11230 35758 11282 35810
rect 11790 35758 11842 35810
rect 12462 35758 12514 35810
rect 12910 35758 12962 35810
rect 14030 35758 14082 35810
rect 18062 35758 18114 35810
rect 20414 35758 20466 35810
rect 36318 35758 36370 35810
rect 36430 35758 36482 35810
rect 37438 35758 37490 35810
rect 38222 35758 38274 35810
rect 42926 35758 42978 35810
rect 43710 35758 43762 35810
rect 44606 35758 44658 35810
rect 50542 35758 50594 35810
rect 51550 35758 51602 35810
rect 51886 35758 51938 35810
rect 54014 35758 54066 35810
rect 56590 35758 56642 35810
rect 57486 35758 57538 35810
rect 58046 35758 58098 35810
rect 4958 35646 5010 35698
rect 6526 35646 6578 35698
rect 6974 35646 7026 35698
rect 8990 35646 9042 35698
rect 10222 35646 10274 35698
rect 10334 35646 10386 35698
rect 10670 35646 10722 35698
rect 14254 35646 14306 35698
rect 14814 35646 14866 35698
rect 15374 35646 15426 35698
rect 19854 35646 19906 35698
rect 20078 35646 20130 35698
rect 24110 35646 24162 35698
rect 24670 35646 24722 35698
rect 30046 35646 30098 35698
rect 30718 35646 30770 35698
rect 31502 35646 31554 35698
rect 35310 35646 35362 35698
rect 38446 35646 38498 35698
rect 38670 35646 38722 35698
rect 38894 35646 38946 35698
rect 39566 35646 39618 35698
rect 39902 35646 39954 35698
rect 40910 35646 40962 35698
rect 43150 35646 43202 35698
rect 43598 35646 43650 35698
rect 45166 35646 45218 35698
rect 46846 35646 46898 35698
rect 48190 35646 48242 35698
rect 48526 35646 48578 35698
rect 48750 35646 48802 35698
rect 50430 35646 50482 35698
rect 50654 35646 50706 35698
rect 52222 35646 52274 35698
rect 52894 35646 52946 35698
rect 57710 35646 57762 35698
rect 5294 35534 5346 35586
rect 6078 35534 6130 35586
rect 6414 35534 6466 35586
rect 7758 35534 7810 35586
rect 6078 35422 6130 35474
rect 10110 35534 10162 35586
rect 13246 35534 13298 35586
rect 16046 35534 16098 35586
rect 18846 35534 18898 35586
rect 19294 35534 19346 35586
rect 20862 35534 20914 35586
rect 21422 35534 21474 35586
rect 21870 35534 21922 35586
rect 25566 35534 25618 35586
rect 26126 35534 26178 35586
rect 30606 35534 30658 35586
rect 32734 35534 32786 35586
rect 34750 35534 34802 35586
rect 41470 35534 41522 35586
rect 41918 35534 41970 35586
rect 43486 35534 43538 35586
rect 47742 35534 47794 35586
rect 49534 35534 49586 35586
rect 11342 35422 11394 35474
rect 20302 35422 20354 35474
rect 36430 35422 36482 35474
rect 40686 35422 40738 35474
rect 45390 35422 45442 35474
rect 46622 35422 46674 35474
rect 56254 35422 56306 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 4062 35086 4114 35138
rect 4286 35086 4338 35138
rect 4846 35086 4898 35138
rect 8654 35086 8706 35138
rect 10334 35086 10386 35138
rect 15374 35086 15426 35138
rect 18286 35086 18338 35138
rect 32398 35086 32450 35138
rect 36094 35086 36146 35138
rect 36430 35086 36482 35138
rect 41022 35086 41074 35138
rect 6190 34974 6242 35026
rect 7198 34974 7250 35026
rect 9102 34974 9154 35026
rect 9550 34974 9602 35026
rect 12238 34974 12290 35026
rect 14366 34974 14418 35026
rect 17390 34974 17442 35026
rect 18398 34974 18450 35026
rect 19854 34974 19906 35026
rect 20302 34974 20354 35026
rect 24334 34974 24386 35026
rect 28366 34974 28418 35026
rect 32958 34974 33010 35026
rect 39006 34974 39058 35026
rect 42142 34974 42194 35026
rect 49646 34974 49698 35026
rect 56926 34974 56978 35026
rect 2830 34862 2882 34914
rect 3502 34862 3554 34914
rect 5070 34862 5122 34914
rect 6302 34862 6354 34914
rect 7870 34862 7922 34914
rect 8094 34862 8146 34914
rect 10110 34862 10162 34914
rect 10670 34862 10722 34914
rect 11342 34862 11394 34914
rect 11790 34862 11842 34914
rect 13694 34862 13746 34914
rect 14814 34862 14866 34914
rect 16942 34862 16994 34914
rect 20526 34862 20578 34914
rect 23214 34862 23266 34914
rect 23774 34862 23826 34914
rect 27358 34862 27410 34914
rect 27806 34862 27858 34914
rect 32510 34862 32562 34914
rect 36094 34862 36146 34914
rect 37774 34862 37826 34914
rect 38558 34862 38610 34914
rect 39230 34862 39282 34914
rect 40574 34862 40626 34914
rect 42030 34862 42082 34914
rect 48526 34862 48578 34914
rect 51662 34862 51714 34914
rect 51998 34862 52050 34914
rect 53790 34862 53842 34914
rect 54462 34862 54514 34914
rect 55358 34862 55410 34914
rect 57038 34862 57090 34914
rect 1934 34750 1986 34802
rect 4510 34750 4562 34802
rect 6078 34750 6130 34802
rect 6638 34750 6690 34802
rect 8430 34750 8482 34802
rect 13806 34750 13858 34802
rect 15822 34750 15874 34802
rect 15934 34750 15986 34802
rect 16046 34750 16098 34802
rect 18846 34750 18898 34802
rect 21982 34750 22034 34802
rect 22430 34750 22482 34802
rect 23886 34750 23938 34802
rect 30046 34750 30098 34802
rect 33630 34750 33682 34802
rect 40686 34750 40738 34802
rect 44382 34750 44434 34802
rect 46062 34750 46114 34802
rect 46398 34750 46450 34802
rect 48638 34750 48690 34802
rect 53454 34750 53506 34802
rect 53566 34750 53618 34802
rect 56590 34750 56642 34802
rect 4062 34638 4114 34690
rect 4734 34638 4786 34690
rect 7758 34638 7810 34690
rect 12910 34638 12962 34690
rect 19294 34638 19346 34690
rect 21646 34638 21698 34690
rect 25118 34638 25170 34690
rect 31838 34638 31890 34690
rect 32398 34638 32450 34690
rect 33742 34638 33794 34690
rect 33966 34638 34018 34690
rect 34414 34638 34466 34690
rect 35646 34638 35698 34690
rect 37550 34638 37602 34690
rect 38782 34638 38834 34690
rect 39006 34638 39058 34690
rect 43934 34638 43986 34690
rect 44830 34638 44882 34690
rect 45502 34638 45554 34690
rect 46846 34638 46898 34690
rect 47294 34638 47346 34690
rect 47742 34638 47794 34690
rect 52446 34638 52498 34690
rect 54686 34638 54738 34690
rect 55694 34638 55746 34690
rect 58046 34638 58098 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4622 34302 4674 34354
rect 6526 34302 6578 34354
rect 6974 34302 7026 34354
rect 10558 34302 10610 34354
rect 11006 34302 11058 34354
rect 14590 34302 14642 34354
rect 16270 34302 16322 34354
rect 16606 34302 16658 34354
rect 24334 34302 24386 34354
rect 24894 34302 24946 34354
rect 29822 34302 29874 34354
rect 30942 34302 30994 34354
rect 31166 34302 31218 34354
rect 31726 34302 31778 34354
rect 37998 34302 38050 34354
rect 40574 34302 40626 34354
rect 46398 34302 46450 34354
rect 47630 34302 47682 34354
rect 49758 34302 49810 34354
rect 51326 34302 51378 34354
rect 52446 34302 52498 34354
rect 55582 34302 55634 34354
rect 55806 34302 55858 34354
rect 6414 34190 6466 34242
rect 7982 34190 8034 34242
rect 9102 34190 9154 34242
rect 11230 34190 11282 34242
rect 11342 34190 11394 34242
rect 13806 34190 13858 34242
rect 14142 34190 14194 34242
rect 17950 34190 18002 34242
rect 20638 34190 20690 34242
rect 26350 34190 26402 34242
rect 27022 34190 27074 34242
rect 30046 34190 30098 34242
rect 34638 34190 34690 34242
rect 38110 34190 38162 34242
rect 40014 34190 40066 34242
rect 40462 34190 40514 34242
rect 42142 34190 42194 34242
rect 47294 34190 47346 34242
rect 49646 34190 49698 34242
rect 50654 34190 50706 34242
rect 52782 34190 52834 34242
rect 53678 34190 53730 34242
rect 55470 34190 55522 34242
rect 56366 34190 56418 34242
rect 57486 34190 57538 34242
rect 5966 34078 6018 34130
rect 6190 34078 6242 34130
rect 7198 34078 7250 34130
rect 9774 34078 9826 34130
rect 9998 34078 10050 34130
rect 10110 34078 10162 34130
rect 18062 34078 18114 34130
rect 18622 34078 18674 34130
rect 19742 34078 19794 34130
rect 21198 34078 21250 34130
rect 21758 34078 21810 34130
rect 25902 34078 25954 34130
rect 26574 34078 26626 34130
rect 27918 34078 27970 34130
rect 30158 34078 30210 34130
rect 30718 34078 30770 34130
rect 30830 34078 30882 34130
rect 33966 34078 34018 34130
rect 36318 34078 36370 34130
rect 37214 34078 37266 34130
rect 38446 34078 38498 34130
rect 40798 34078 40850 34130
rect 41694 34078 41746 34130
rect 41918 34078 41970 34130
rect 43038 34078 43090 34130
rect 44270 34078 44322 34130
rect 44942 34078 44994 34130
rect 45166 34078 45218 34130
rect 46734 34078 46786 34130
rect 49870 34078 49922 34130
rect 50206 34078 50258 34130
rect 51886 34078 51938 34130
rect 53790 34078 53842 34130
rect 54686 34078 54738 34130
rect 56590 34078 56642 34130
rect 5070 33966 5122 34018
rect 5406 33966 5458 34018
rect 8542 33966 8594 34018
rect 12798 33966 12850 34018
rect 13246 33966 13298 34018
rect 15038 33966 15090 34018
rect 15822 33966 15874 34018
rect 20414 33966 20466 34018
rect 26462 33966 26514 34018
rect 29486 33966 29538 34018
rect 33742 33966 33794 34018
rect 35198 33966 35250 34018
rect 35870 33966 35922 34018
rect 37550 33966 37602 34018
rect 38894 33966 38946 34018
rect 43934 33966 43986 34018
rect 45054 33966 45106 34018
rect 48190 33966 48242 34018
rect 48526 33966 48578 34018
rect 54910 33966 54962 34018
rect 58046 33966 58098 34018
rect 7870 33854 7922 33906
rect 34974 33854 35026 33906
rect 35198 33854 35250 33906
rect 44046 33854 44098 33906
rect 53678 33854 53730 33906
rect 54350 33854 54402 33906
rect 57598 33854 57650 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 4398 33518 4450 33570
rect 26910 33518 26962 33570
rect 27918 33518 27970 33570
rect 37438 33518 37490 33570
rect 37886 33518 37938 33570
rect 51438 33518 51490 33570
rect 8318 33406 8370 33458
rect 15150 33406 15202 33458
rect 17614 33406 17666 33458
rect 22094 33406 22146 33458
rect 22542 33406 22594 33458
rect 27358 33406 27410 33458
rect 29710 33406 29762 33458
rect 34190 33406 34242 33458
rect 36766 33406 36818 33458
rect 37438 33406 37490 33458
rect 40574 33406 40626 33458
rect 48414 33406 48466 33458
rect 50430 33406 50482 33458
rect 51550 33406 51602 33458
rect 54350 33406 54402 33458
rect 56254 33406 56306 33458
rect 4510 33294 4562 33346
rect 4734 33294 4786 33346
rect 5742 33294 5794 33346
rect 6750 33294 6802 33346
rect 7982 33294 8034 33346
rect 9214 33294 9266 33346
rect 23662 33294 23714 33346
rect 27582 33294 27634 33346
rect 28478 33294 28530 33346
rect 29934 33294 29986 33346
rect 31950 33294 32002 33346
rect 32510 33294 32562 33346
rect 33294 33294 33346 33346
rect 33518 33294 33570 33346
rect 36318 33294 36370 33346
rect 39790 33294 39842 33346
rect 40014 33294 40066 33346
rect 41582 33294 41634 33346
rect 44158 33294 44210 33346
rect 47966 33294 48018 33346
rect 48526 33294 48578 33346
rect 50990 33294 51042 33346
rect 53902 33294 53954 33346
rect 54238 33294 54290 33346
rect 54574 33294 54626 33346
rect 5854 33182 5906 33234
rect 7310 33182 7362 33234
rect 8318 33182 8370 33234
rect 8542 33182 8594 33234
rect 12462 33182 12514 33234
rect 23102 33182 23154 33234
rect 23438 33182 23490 33234
rect 24446 33182 24498 33234
rect 28814 33182 28866 33234
rect 39678 33182 39730 33234
rect 41806 33182 41858 33234
rect 41918 33182 41970 33234
rect 42030 33182 42082 33234
rect 45502 33182 45554 33234
rect 47182 33182 47234 33234
rect 49086 33182 49138 33234
rect 55918 33182 55970 33234
rect 57150 33182 57202 33234
rect 7198 33070 7250 33122
rect 8206 33070 8258 33122
rect 9662 33070 9714 33122
rect 12126 33070 12178 33122
rect 12350 33070 12402 33122
rect 12910 33070 12962 33122
rect 13694 33070 13746 33122
rect 14030 33070 14082 33122
rect 16158 33070 16210 33122
rect 16270 33070 16322 33122
rect 16382 33070 16434 33122
rect 16606 33070 16658 33122
rect 17278 33070 17330 33122
rect 19182 33070 19234 33122
rect 19854 33070 19906 33122
rect 20862 33070 20914 33122
rect 30270 33070 30322 33122
rect 30830 33070 30882 33122
rect 32398 33070 32450 33122
rect 32622 33070 32674 33122
rect 34750 33070 34802 33122
rect 35422 33070 35474 33122
rect 35982 33070 36034 33122
rect 37886 33070 37938 33122
rect 38446 33070 38498 33122
rect 39230 33070 39282 33122
rect 40910 33070 40962 33122
rect 41694 33070 41746 33122
rect 42926 33070 42978 33122
rect 43262 33070 43314 33122
rect 43710 33070 43762 33122
rect 44606 33070 44658 33122
rect 45614 33070 45666 33122
rect 45726 33070 45778 33122
rect 46398 33070 46450 33122
rect 46734 33070 46786 33122
rect 49534 33070 49586 33122
rect 50318 33070 50370 33122
rect 50542 33070 50594 33122
rect 51662 33070 51714 33122
rect 52334 33070 52386 33122
rect 52670 33070 52722 33122
rect 53342 33070 53394 33122
rect 56142 33070 56194 33122
rect 56366 33070 56418 33122
rect 57486 33070 57538 33122
rect 57934 33070 57986 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 4734 32734 4786 32786
rect 6526 32734 6578 32786
rect 7646 32734 7698 32786
rect 8654 32734 8706 32786
rect 13582 32734 13634 32786
rect 17726 32734 17778 32786
rect 21870 32734 21922 32786
rect 22878 32734 22930 32786
rect 25790 32734 25842 32786
rect 26014 32734 26066 32786
rect 26910 32734 26962 32786
rect 35310 32734 35362 32786
rect 38558 32734 38610 32786
rect 39454 32734 39506 32786
rect 39790 32734 39842 32786
rect 40350 32734 40402 32786
rect 41806 32734 41858 32786
rect 45278 32734 45330 32786
rect 46398 32734 46450 32786
rect 47182 32734 47234 32786
rect 50094 32734 50146 32786
rect 50766 32734 50818 32786
rect 52894 32734 52946 32786
rect 7758 32622 7810 32674
rect 8766 32622 8818 32674
rect 11790 32622 11842 32674
rect 14926 32622 14978 32674
rect 15038 32622 15090 32674
rect 18622 32622 18674 32674
rect 20638 32622 20690 32674
rect 22654 32622 22706 32674
rect 23326 32622 23378 32674
rect 31838 32622 31890 32674
rect 36878 32622 36930 32674
rect 37550 32622 37602 32674
rect 40910 32622 40962 32674
rect 42142 32622 42194 32674
rect 53454 32622 53506 32674
rect 57486 32622 57538 32674
rect 3838 32510 3890 32562
rect 5406 32510 5458 32562
rect 6302 32510 6354 32562
rect 8430 32510 8482 32562
rect 8878 32510 8930 32562
rect 12462 32510 12514 32562
rect 13358 32510 13410 32562
rect 13470 32510 13522 32562
rect 14030 32510 14082 32562
rect 15262 32510 15314 32562
rect 16606 32510 16658 32562
rect 18062 32510 18114 32562
rect 19518 32510 19570 32562
rect 20526 32510 20578 32562
rect 21646 32510 21698 32562
rect 21982 32510 22034 32562
rect 22542 32510 22594 32562
rect 23774 32510 23826 32562
rect 24222 32510 24274 32562
rect 26126 32510 26178 32562
rect 26686 32510 26738 32562
rect 26798 32510 26850 32562
rect 27358 32510 27410 32562
rect 31502 32510 31554 32562
rect 35534 32510 35586 32562
rect 36430 32510 36482 32562
rect 37438 32510 37490 32562
rect 39678 32510 39730 32562
rect 39902 32510 39954 32562
rect 41470 32510 41522 32562
rect 41918 32510 41970 32562
rect 43038 32510 43090 32562
rect 43598 32510 43650 32562
rect 43822 32510 43874 32562
rect 44046 32510 44098 32562
rect 44270 32510 44322 32562
rect 44718 32510 44770 32562
rect 45166 32510 45218 32562
rect 45390 32510 45442 32562
rect 45950 32510 46002 32562
rect 46286 32510 46338 32562
rect 46510 32510 46562 32562
rect 47294 32510 47346 32562
rect 47966 32510 48018 32562
rect 49646 32510 49698 32562
rect 49982 32510 50034 32562
rect 50206 32510 50258 32562
rect 51102 32510 51154 32562
rect 53678 32510 53730 32562
rect 54014 32510 54066 32562
rect 55022 32510 55074 32562
rect 56590 32510 56642 32562
rect 57822 32510 57874 32562
rect 3390 32398 3442 32450
rect 4286 32398 4338 32450
rect 7086 32398 7138 32450
rect 9662 32398 9714 32450
rect 10222 32398 10274 32450
rect 10894 32398 10946 32450
rect 12686 32398 12738 32450
rect 14478 32398 14530 32450
rect 15822 32398 15874 32450
rect 16270 32398 16322 32450
rect 19406 32398 19458 32450
rect 21310 32398 21362 32450
rect 24782 32398 24834 32450
rect 27694 32398 27746 32450
rect 28142 32398 28194 32450
rect 30494 32398 30546 32450
rect 32846 32398 32898 32450
rect 34974 32398 35026 32450
rect 38110 32398 38162 32450
rect 42590 32398 42642 32450
rect 44158 32398 44210 32450
rect 48414 32398 48466 32450
rect 51550 32398 51602 32450
rect 52446 32398 52498 32450
rect 53790 32398 53842 32450
rect 56030 32398 56082 32450
rect 4846 32286 4898 32338
rect 5070 32286 5122 32338
rect 5630 32286 5682 32338
rect 7086 32286 7138 32338
rect 7310 32286 7362 32338
rect 7534 32286 7586 32338
rect 47182 32286 47234 32338
rect 54238 32286 54290 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 14142 31950 14194 32002
rect 14590 31950 14642 32002
rect 22206 31950 22258 32002
rect 23102 31950 23154 32002
rect 44606 31950 44658 32002
rect 48078 31950 48130 32002
rect 6078 31838 6130 31890
rect 8990 31838 9042 31890
rect 10334 31838 10386 31890
rect 11454 31838 11506 31890
rect 12350 31838 12402 31890
rect 13918 31838 13970 31890
rect 15262 31838 15314 31890
rect 16046 31838 16098 31890
rect 17726 31838 17778 31890
rect 20190 31838 20242 31890
rect 20862 31838 20914 31890
rect 21646 31838 21698 31890
rect 33966 31838 34018 31890
rect 34302 31838 34354 31890
rect 36654 31838 36706 31890
rect 40462 31838 40514 31890
rect 46286 31838 46338 31890
rect 46734 31838 46786 31890
rect 48190 31838 48242 31890
rect 53678 31838 53730 31890
rect 55358 31838 55410 31890
rect 56702 31838 56754 31890
rect 8654 31726 8706 31778
rect 8878 31726 8930 31778
rect 9102 31726 9154 31778
rect 9774 31726 9826 31778
rect 12126 31726 12178 31778
rect 13694 31726 13746 31778
rect 15710 31726 15762 31778
rect 18062 31726 18114 31778
rect 21870 31726 21922 31778
rect 23550 31726 23602 31778
rect 23662 31726 23714 31778
rect 24670 31726 24722 31778
rect 33742 31726 33794 31778
rect 34862 31726 34914 31778
rect 35758 31726 35810 31778
rect 37438 31726 37490 31778
rect 39230 31726 39282 31778
rect 39678 31726 39730 31778
rect 41470 31726 41522 31778
rect 42702 31726 42754 31778
rect 43150 31726 43202 31778
rect 44158 31726 44210 31778
rect 44494 31726 44546 31778
rect 46174 31726 46226 31778
rect 46510 31726 46562 31778
rect 47742 31726 47794 31778
rect 48414 31726 48466 31778
rect 49310 31726 49362 31778
rect 51326 31726 51378 31778
rect 51998 31726 52050 31778
rect 52446 31726 52498 31778
rect 52670 31726 52722 31778
rect 54238 31726 54290 31778
rect 54910 31726 54962 31778
rect 55246 31726 55298 31778
rect 56478 31726 56530 31778
rect 57486 31726 57538 31778
rect 57934 31726 57986 31778
rect 4174 31614 4226 31666
rect 7534 31614 7586 31666
rect 18510 31614 18562 31666
rect 20078 31614 20130 31666
rect 23774 31614 23826 31666
rect 24446 31614 24498 31666
rect 26462 31614 26514 31666
rect 31278 31614 31330 31666
rect 35422 31614 35474 31666
rect 37886 31614 37938 31666
rect 38110 31614 38162 31666
rect 44718 31614 44770 31666
rect 49646 31614 49698 31666
rect 50206 31614 50258 31666
rect 50990 31614 51042 31666
rect 53454 31614 53506 31666
rect 53678 31614 53730 31666
rect 56814 31614 56866 31666
rect 2382 31502 2434 31554
rect 2830 31502 2882 31554
rect 3278 31502 3330 31554
rect 3726 31502 3778 31554
rect 4622 31502 4674 31554
rect 5070 31502 5122 31554
rect 5742 31502 5794 31554
rect 6526 31502 6578 31554
rect 6974 31502 7026 31554
rect 10222 31502 10274 31554
rect 10446 31502 10498 31554
rect 10894 31502 10946 31554
rect 13022 31502 13074 31554
rect 19406 31502 19458 31554
rect 20302 31502 20354 31554
rect 28142 31502 28194 31554
rect 30718 31502 30770 31554
rect 31390 31502 31442 31554
rect 35534 31502 35586 31554
rect 36318 31502 36370 31554
rect 36542 31502 36594 31554
rect 36766 31502 36818 31554
rect 37662 31502 37714 31554
rect 38558 31502 38610 31554
rect 40910 31502 40962 31554
rect 42030 31502 42082 31554
rect 44270 31502 44322 31554
rect 49870 31502 49922 31554
rect 52222 31502 52274 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 3726 31166 3778 31218
rect 4622 31166 4674 31218
rect 5070 31166 5122 31218
rect 10894 31166 10946 31218
rect 11902 31166 11954 31218
rect 13134 31166 13186 31218
rect 14702 31166 14754 31218
rect 16494 31166 16546 31218
rect 21646 31166 21698 31218
rect 22430 31166 22482 31218
rect 23662 31166 23714 31218
rect 24782 31166 24834 31218
rect 26014 31166 26066 31218
rect 26126 31166 26178 31218
rect 27358 31166 27410 31218
rect 27582 31166 27634 31218
rect 28254 31166 28306 31218
rect 31950 31166 32002 31218
rect 35758 31166 35810 31218
rect 40910 31166 40962 31218
rect 42926 31166 42978 31218
rect 43038 31166 43090 31218
rect 43822 31166 43874 31218
rect 44830 31166 44882 31218
rect 44942 31166 44994 31218
rect 45054 31166 45106 31218
rect 45838 31166 45890 31218
rect 49422 31166 49474 31218
rect 49758 31166 49810 31218
rect 53118 31166 53170 31218
rect 8318 31054 8370 31106
rect 12686 31054 12738 31106
rect 19406 31054 19458 31106
rect 22766 31054 22818 31106
rect 24894 31054 24946 31106
rect 26238 31054 26290 31106
rect 27694 31054 27746 31106
rect 30382 31054 30434 31106
rect 31166 31054 31218 31106
rect 31502 31054 31554 31106
rect 33630 31054 33682 31106
rect 33966 31054 34018 31106
rect 36542 31054 36594 31106
rect 39790 31054 39842 31106
rect 40798 31054 40850 31106
rect 42814 31054 42866 31106
rect 47070 31054 47122 31106
rect 48638 31054 48690 31106
rect 49534 31054 49586 31106
rect 50878 31054 50930 31106
rect 50990 31054 51042 31106
rect 52334 31054 52386 31106
rect 54798 31054 54850 31106
rect 56366 31054 56418 31106
rect 57486 31054 57538 31106
rect 5294 30942 5346 30994
rect 8094 30942 8146 30994
rect 8542 30942 8594 30994
rect 8766 30942 8818 30994
rect 12238 30942 12290 30994
rect 19854 30942 19906 30994
rect 21534 30942 21586 30994
rect 22318 30942 22370 30994
rect 22542 30942 22594 30994
rect 24558 30942 24610 30994
rect 25566 30942 25618 30994
rect 29934 30942 29986 30994
rect 33854 30942 33906 30994
rect 35646 30942 35698 30994
rect 37886 30942 37938 30994
rect 39678 30942 39730 30994
rect 40350 30942 40402 30994
rect 40574 30942 40626 30994
rect 43934 30942 43986 30994
rect 44158 30942 44210 30994
rect 45502 30942 45554 30994
rect 47518 30942 47570 30994
rect 48302 30942 48354 30994
rect 49982 30942 50034 30994
rect 51662 30942 51714 30994
rect 53678 30942 53730 30994
rect 55358 30942 55410 30994
rect 56702 30942 56754 30994
rect 57710 30942 57762 30994
rect 1934 30830 1986 30882
rect 2270 30830 2322 30882
rect 2830 30830 2882 30882
rect 3166 30830 3218 30882
rect 4174 30830 4226 30882
rect 6190 30830 6242 30882
rect 6638 30830 6690 30882
rect 7086 30830 7138 30882
rect 7534 30830 7586 30882
rect 8430 30830 8482 30882
rect 9662 30830 9714 30882
rect 10558 30830 10610 30882
rect 11454 30830 11506 30882
rect 13918 30830 13970 30882
rect 14366 30830 14418 30882
rect 15262 30830 15314 30882
rect 16046 30830 16098 30882
rect 16942 30830 16994 30882
rect 17726 30830 17778 30882
rect 18398 30830 18450 30882
rect 18846 30830 18898 30882
rect 24110 30830 24162 30882
rect 30158 30830 30210 30882
rect 34190 30830 34242 30882
rect 34974 30830 35026 30882
rect 41470 30830 41522 30882
rect 42590 30830 42642 30882
rect 46286 30830 46338 30882
rect 1934 30718 1986 30770
rect 2830 30718 2882 30770
rect 13918 30718 13970 30770
rect 14702 30718 14754 30770
rect 18510 30718 18562 30770
rect 18846 30718 18898 30770
rect 23550 30718 23602 30770
rect 23774 30718 23826 30770
rect 24110 30718 24162 30770
rect 34414 30718 34466 30770
rect 42142 30718 42194 30770
rect 42366 30718 42418 30770
rect 43822 30718 43874 30770
rect 47406 30718 47458 30770
rect 50878 30718 50930 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 3166 30382 3218 30434
rect 3614 30382 3666 30434
rect 4286 30382 4338 30434
rect 6190 30382 6242 30434
rect 6862 30382 6914 30434
rect 8654 30382 8706 30434
rect 8878 30382 8930 30434
rect 9774 30382 9826 30434
rect 15374 30382 15426 30434
rect 15710 30382 15762 30434
rect 21758 30382 21810 30434
rect 22094 30382 22146 30434
rect 24334 30382 24386 30434
rect 29710 30382 29762 30434
rect 31502 30382 31554 30434
rect 44606 30382 44658 30434
rect 47294 30382 47346 30434
rect 51326 30382 51378 30434
rect 52558 30382 52610 30434
rect 5742 30270 5794 30322
rect 5966 30270 6018 30322
rect 8318 30270 8370 30322
rect 17726 30270 17778 30322
rect 23662 30270 23714 30322
rect 24222 30270 24274 30322
rect 25342 30270 25394 30322
rect 40238 30270 40290 30322
rect 44270 30270 44322 30322
rect 51214 30270 51266 30322
rect 56926 30270 56978 30322
rect 2382 30158 2434 30210
rect 6414 30158 6466 30210
rect 9102 30158 9154 30210
rect 11678 30158 11730 30210
rect 13918 30158 13970 30210
rect 19742 30158 19794 30210
rect 20078 30158 20130 30210
rect 20638 30158 20690 30210
rect 23214 30158 23266 30210
rect 24446 30158 24498 30210
rect 28142 30158 28194 30210
rect 30942 30158 30994 30210
rect 31502 30158 31554 30210
rect 32286 30158 32338 30210
rect 34750 30158 34802 30210
rect 35086 30158 35138 30210
rect 39006 30158 39058 30210
rect 40462 30158 40514 30210
rect 42030 30158 42082 30210
rect 44046 30158 44098 30210
rect 45726 30158 45778 30210
rect 46174 30158 46226 30210
rect 47406 30158 47458 30210
rect 49422 30158 49474 30210
rect 52446 30158 52498 30210
rect 53790 30158 53842 30210
rect 54238 30158 54290 30210
rect 54686 30158 54738 30210
rect 56702 30158 56754 30210
rect 57374 30158 57426 30210
rect 3726 30046 3778 30098
rect 8094 30046 8146 30098
rect 11006 30046 11058 30098
rect 11118 30046 11170 30098
rect 14142 30046 14194 30098
rect 14366 30046 14418 30098
rect 14590 30046 14642 30098
rect 15150 30046 15202 30098
rect 18734 30046 18786 30098
rect 19294 30046 19346 30098
rect 20862 30046 20914 30098
rect 21982 30046 22034 30098
rect 28702 30046 28754 30098
rect 28814 30046 28866 30098
rect 29598 30046 29650 30098
rect 30830 30046 30882 30098
rect 31166 30046 31218 30098
rect 31390 30046 31442 30098
rect 31838 30046 31890 30098
rect 34190 30046 34242 30098
rect 35646 30046 35698 30098
rect 37886 30046 37938 30098
rect 40798 30046 40850 30098
rect 41246 30046 41298 30098
rect 42142 30046 42194 30098
rect 42366 30046 42418 30098
rect 42590 30046 42642 30098
rect 48862 30046 48914 30098
rect 50990 30046 51042 30098
rect 55582 30046 55634 30098
rect 56254 30046 56306 30098
rect 1934 29934 1986 29986
rect 2830 29934 2882 29986
rect 3278 29934 3330 29986
rect 4174 29934 4226 29986
rect 4622 29934 4674 29986
rect 5070 29934 5122 29986
rect 7646 29934 7698 29986
rect 9550 29934 9602 29986
rect 10110 29934 10162 29986
rect 10446 29934 10498 29986
rect 11342 29934 11394 29986
rect 12462 29934 12514 29986
rect 12686 29934 12738 29986
rect 12798 29934 12850 29986
rect 12910 29934 12962 29986
rect 16270 29934 16322 29986
rect 16830 29934 16882 29986
rect 17278 29934 17330 29986
rect 18398 29934 18450 29986
rect 19854 29934 19906 29986
rect 25902 29934 25954 29986
rect 26238 29934 26290 29986
rect 28478 29934 28530 29986
rect 29710 29934 29762 29986
rect 30494 29934 30546 29986
rect 30718 29934 30770 29986
rect 33182 29934 33234 29986
rect 37550 29934 37602 29986
rect 43038 29934 43090 29986
rect 43486 29934 43538 29986
rect 45390 29934 45442 29986
rect 45614 29934 45666 29986
rect 46622 29934 46674 29986
rect 50206 29934 50258 29986
rect 53342 29934 53394 29986
rect 55134 29934 55186 29986
rect 57822 29934 57874 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 2158 29598 2210 29650
rect 2494 29598 2546 29650
rect 2942 29598 2994 29650
rect 5294 29598 5346 29650
rect 7646 29598 7698 29650
rect 8430 29598 8482 29650
rect 8542 29598 8594 29650
rect 8654 29598 8706 29650
rect 18062 29598 18114 29650
rect 20974 29598 21026 29650
rect 21870 29598 21922 29650
rect 26126 29598 26178 29650
rect 26238 29598 26290 29650
rect 29486 29598 29538 29650
rect 32846 29598 32898 29650
rect 33518 29598 33570 29650
rect 35198 29598 35250 29650
rect 38334 29598 38386 29650
rect 38446 29598 38498 29650
rect 39342 29598 39394 29650
rect 44718 29598 44770 29650
rect 47966 29598 48018 29650
rect 54238 29598 54290 29650
rect 55022 29598 55074 29650
rect 56366 29598 56418 29650
rect 57486 29598 57538 29650
rect 4846 29486 4898 29538
rect 7534 29486 7586 29538
rect 11678 29486 11730 29538
rect 13582 29486 13634 29538
rect 16830 29486 16882 29538
rect 20190 29486 20242 29538
rect 22654 29486 22706 29538
rect 23774 29486 23826 29538
rect 27582 29486 27634 29538
rect 29374 29486 29426 29538
rect 30270 29486 30322 29538
rect 32510 29486 32562 29538
rect 37998 29486 38050 29538
rect 38222 29486 38274 29538
rect 39006 29486 39058 29538
rect 41582 29486 41634 29538
rect 44046 29486 44098 29538
rect 46398 29486 46450 29538
rect 48078 29486 48130 29538
rect 50878 29486 50930 29538
rect 53566 29486 53618 29538
rect 5630 29374 5682 29426
rect 6974 29374 7026 29426
rect 7310 29374 7362 29426
rect 9102 29374 9154 29426
rect 10446 29374 10498 29426
rect 11566 29374 11618 29426
rect 13470 29374 13522 29426
rect 14254 29374 14306 29426
rect 15710 29374 15762 29426
rect 16270 29374 16322 29426
rect 18622 29374 18674 29426
rect 19630 29374 19682 29426
rect 20414 29374 20466 29426
rect 23550 29374 23602 29426
rect 24334 29374 24386 29426
rect 25566 29374 25618 29426
rect 26014 29374 26066 29426
rect 26686 29374 26738 29426
rect 27358 29374 27410 29426
rect 30718 29374 30770 29426
rect 31054 29374 31106 29426
rect 34638 29374 34690 29426
rect 36318 29374 36370 29426
rect 36878 29374 36930 29426
rect 39342 29374 39394 29426
rect 39678 29374 39730 29426
rect 40126 29374 40178 29426
rect 40350 29374 40402 29426
rect 40798 29374 40850 29426
rect 41918 29374 41970 29426
rect 43374 29374 43426 29426
rect 44942 29374 44994 29426
rect 46958 29374 47010 29426
rect 48750 29374 48802 29426
rect 49758 29374 49810 29426
rect 53230 29374 53282 29426
rect 54910 29374 54962 29426
rect 55134 29374 55186 29426
rect 56030 29374 56082 29426
rect 56478 29374 56530 29426
rect 56702 29374 56754 29426
rect 57710 29374 57762 29426
rect 3502 29262 3554 29314
rect 3950 29262 4002 29314
rect 4398 29262 4450 29314
rect 5854 29262 5906 29314
rect 6526 29262 6578 29314
rect 9998 29262 10050 29314
rect 11006 29262 11058 29314
rect 19182 29262 19234 29314
rect 21534 29262 21586 29314
rect 22430 29262 22482 29314
rect 22766 29262 22818 29314
rect 23998 29262 24050 29314
rect 24110 29262 24162 29314
rect 28030 29262 28082 29314
rect 30830 29262 30882 29314
rect 31726 29262 31778 29314
rect 34302 29262 34354 29314
rect 36990 29262 37042 29314
rect 40238 29262 40290 29314
rect 42366 29262 42418 29314
rect 48638 29262 48690 29314
rect 49982 29262 50034 29314
rect 52334 29262 52386 29314
rect 55358 29262 55410 29314
rect 10782 29150 10834 29202
rect 29598 29150 29650 29202
rect 36094 29150 36146 29202
rect 47966 29150 48018 29202
rect 50094 29150 50146 29202
rect 50990 29150 51042 29202
rect 51214 29150 51266 29202
rect 51326 29150 51378 29202
rect 55582 29150 55634 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 5854 28814 5906 28866
rect 7758 28814 7810 28866
rect 11230 28814 11282 28866
rect 17950 28814 18002 28866
rect 22206 28814 22258 28866
rect 22766 28814 22818 28866
rect 24110 28814 24162 28866
rect 24670 28814 24722 28866
rect 31278 28814 31330 28866
rect 47406 28814 47458 28866
rect 49422 28814 49474 28866
rect 3726 28702 3778 28754
rect 4174 28702 4226 28754
rect 4622 28702 4674 28754
rect 5070 28702 5122 28754
rect 5966 28702 6018 28754
rect 10894 28702 10946 28754
rect 12910 28702 12962 28754
rect 13806 28702 13858 28754
rect 19406 28702 19458 28754
rect 21758 28702 21810 28754
rect 23774 28702 23826 28754
rect 24782 28702 24834 28754
rect 28702 28702 28754 28754
rect 32286 28702 32338 28754
rect 33070 28702 33122 28754
rect 33966 28702 34018 28754
rect 34974 28702 35026 28754
rect 37550 28702 37602 28754
rect 38894 28702 38946 28754
rect 39230 28702 39282 28754
rect 45390 28702 45442 28754
rect 47070 28702 47122 28754
rect 48974 28702 49026 28754
rect 53678 28702 53730 28754
rect 56142 28702 56194 28754
rect 2942 28590 2994 28642
rect 7086 28590 7138 28642
rect 7310 28590 7362 28642
rect 8654 28590 8706 28642
rect 9326 28590 9378 28642
rect 11230 28590 11282 28642
rect 14030 28590 14082 28642
rect 14254 28590 14306 28642
rect 16270 28590 16322 28642
rect 16830 28590 16882 28642
rect 17278 28590 17330 28642
rect 18174 28590 18226 28642
rect 18510 28590 18562 28642
rect 19294 28590 19346 28642
rect 20974 28590 21026 28642
rect 22206 28590 22258 28642
rect 22654 28590 22706 28642
rect 23102 28590 23154 28642
rect 23550 28590 23602 28642
rect 26686 28590 26738 28642
rect 27918 28590 27970 28642
rect 30606 28590 30658 28642
rect 33518 28590 33570 28642
rect 35534 28590 35586 28642
rect 35870 28590 35922 28642
rect 36430 28590 36482 28642
rect 39678 28590 39730 28642
rect 40686 28590 40738 28642
rect 42814 28590 42866 28642
rect 44382 28590 44434 28642
rect 46510 28590 46562 28642
rect 47518 28590 47570 28642
rect 48638 28590 48690 28642
rect 49534 28590 49586 28642
rect 52334 28590 52386 28642
rect 52558 28590 52610 28642
rect 54014 28590 54066 28642
rect 54238 28590 54290 28642
rect 56030 28590 56082 28642
rect 56702 28590 56754 28642
rect 57710 28590 57762 28642
rect 1934 28478 1986 28530
rect 7198 28478 7250 28530
rect 9998 28478 10050 28530
rect 15598 28478 15650 28530
rect 15822 28478 15874 28530
rect 19742 28478 19794 28530
rect 24894 28478 24946 28530
rect 26350 28478 26402 28530
rect 27358 28478 27410 28530
rect 30270 28478 30322 28530
rect 31278 28478 31330 28530
rect 31390 28478 31442 28530
rect 32174 28478 32226 28530
rect 32398 28478 32450 28530
rect 34526 28478 34578 28530
rect 34750 28478 34802 28530
rect 36766 28478 36818 28530
rect 37774 28478 37826 28530
rect 37998 28478 38050 28530
rect 38334 28478 38386 28530
rect 40574 28478 40626 28530
rect 44718 28478 44770 28530
rect 46062 28478 46114 28530
rect 49870 28478 49922 28530
rect 50654 28478 50706 28530
rect 50990 28478 51042 28530
rect 51214 28478 51266 28530
rect 51774 28478 51826 28530
rect 51998 28478 52050 28530
rect 52110 28478 52162 28530
rect 56254 28478 56306 28530
rect 57150 28478 57202 28530
rect 57374 28478 57426 28530
rect 6078 28366 6130 28418
rect 15710 28366 15762 28418
rect 20526 28366 20578 28418
rect 25902 28366 25954 28418
rect 27134 28366 27186 28418
rect 27246 28366 27298 28418
rect 28254 28366 28306 28418
rect 34974 28366 35026 28418
rect 36654 28366 36706 28418
rect 38110 28366 38162 28418
rect 40798 28366 40850 28418
rect 50878 28366 50930 28418
rect 53566 28366 53618 28418
rect 53790 28366 53842 28418
rect 55134 28366 55186 28418
rect 55470 28366 55522 28418
rect 57598 28366 57650 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 5294 28030 5346 28082
rect 6526 28030 6578 28082
rect 8430 28030 8482 28082
rect 9774 28030 9826 28082
rect 10222 28030 10274 28082
rect 10670 28030 10722 28082
rect 12014 28030 12066 28082
rect 13022 28030 13074 28082
rect 16046 28030 16098 28082
rect 16942 28030 16994 28082
rect 18734 28030 18786 28082
rect 18846 28030 18898 28082
rect 20750 28030 20802 28082
rect 23662 28030 23714 28082
rect 23998 28030 24050 28082
rect 24670 28030 24722 28082
rect 24894 28030 24946 28082
rect 31054 28030 31106 28082
rect 31166 28030 31218 28082
rect 31726 28030 31778 28082
rect 32622 28030 32674 28082
rect 39342 28030 39394 28082
rect 40014 28030 40066 28082
rect 41582 28030 41634 28082
rect 42814 28030 42866 28082
rect 47854 28030 47906 28082
rect 49870 28030 49922 28082
rect 53006 28030 53058 28082
rect 3166 27918 3218 27970
rect 11454 27918 11506 27970
rect 14030 27918 14082 27970
rect 14254 27918 14306 27970
rect 14366 27918 14418 27970
rect 16718 27918 16770 27970
rect 18174 27918 18226 27970
rect 21982 27918 22034 27970
rect 22654 27918 22706 27970
rect 26126 27918 26178 27970
rect 28142 27918 28194 27970
rect 28254 27918 28306 27970
rect 34190 27918 34242 27970
rect 35534 27918 35586 27970
rect 36654 27918 36706 27970
rect 37550 27918 37602 27970
rect 39230 27918 39282 27970
rect 40574 27918 40626 27970
rect 50430 27918 50482 27970
rect 50654 27918 50706 27970
rect 51886 27918 51938 27970
rect 52110 27918 52162 27970
rect 53118 27918 53170 27970
rect 57486 27918 57538 27970
rect 57822 27918 57874 27970
rect 3950 27806 4002 27858
rect 7198 27806 7250 27858
rect 7422 27806 7474 27858
rect 7646 27806 7698 27858
rect 7870 27806 7922 27858
rect 8766 27806 8818 27858
rect 11678 27806 11730 27858
rect 12238 27806 12290 27858
rect 12798 27806 12850 27858
rect 13022 27806 13074 27858
rect 13246 27806 13298 27858
rect 13358 27806 13410 27858
rect 15262 27806 15314 27858
rect 16606 27806 16658 27858
rect 18622 27806 18674 27858
rect 19182 27806 19234 27858
rect 19742 27806 19794 27858
rect 20302 27806 20354 27858
rect 20862 27806 20914 27858
rect 22206 27806 22258 27858
rect 22766 27806 22818 27858
rect 24558 27806 24610 27858
rect 26462 27806 26514 27858
rect 27134 27806 27186 27858
rect 30606 27806 30658 27858
rect 31278 27806 31330 27858
rect 34414 27806 34466 27858
rect 35198 27806 35250 27858
rect 36766 27806 36818 27858
rect 37326 27806 37378 27858
rect 38558 27806 38610 27858
rect 42702 27806 42754 27858
rect 42926 27806 42978 27858
rect 43262 27806 43314 27858
rect 43934 27806 43986 27858
rect 44942 27806 44994 27858
rect 45726 27806 45778 27858
rect 46846 27806 46898 27858
rect 47742 27806 47794 27858
rect 47966 27806 48018 27858
rect 49646 27806 49698 27858
rect 53006 27806 53058 27858
rect 54574 27806 54626 27858
rect 56030 27806 56082 27858
rect 1822 27694 1874 27746
rect 2270 27694 2322 27746
rect 2718 27694 2770 27746
rect 3614 27694 3666 27746
rect 4398 27694 4450 27746
rect 4958 27694 5010 27746
rect 5854 27694 5906 27746
rect 7758 27694 7810 27746
rect 8990 27694 9042 27746
rect 15710 27694 15762 27746
rect 17726 27694 17778 27746
rect 25566 27694 25618 27746
rect 26798 27694 26850 27746
rect 28702 27694 28754 27746
rect 34190 27694 34242 27746
rect 36878 27694 36930 27746
rect 42142 27694 42194 27746
rect 44046 27694 44098 27746
rect 44494 27694 44546 27746
rect 45950 27694 46002 27746
rect 46958 27694 47010 27746
rect 50542 27694 50594 27746
rect 51214 27694 51266 27746
rect 52222 27694 52274 27746
rect 1822 27582 1874 27634
rect 3278 27582 3330 27634
rect 6302 27582 6354 27634
rect 6638 27582 6690 27634
rect 15150 27582 15202 27634
rect 15934 27582 15986 27634
rect 25454 27582 25506 27634
rect 26014 27582 26066 27634
rect 28142 27582 28194 27634
rect 39342 27582 39394 27634
rect 41918 27582 41970 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 7198 27246 7250 27298
rect 8094 27246 8146 27298
rect 8318 27246 8370 27298
rect 15150 27246 15202 27298
rect 15934 27246 15986 27298
rect 16270 27246 16322 27298
rect 20638 27246 20690 27298
rect 23774 27246 23826 27298
rect 33854 27246 33906 27298
rect 34190 27246 34242 27298
rect 40686 27246 40738 27298
rect 43374 27246 43426 27298
rect 47854 27246 47906 27298
rect 48302 27246 48354 27298
rect 51886 27246 51938 27298
rect 53566 27246 53618 27298
rect 55806 27246 55858 27298
rect 56142 27246 56194 27298
rect 4958 27134 5010 27186
rect 6190 27134 6242 27186
rect 8094 27134 8146 27186
rect 8430 27134 8482 27186
rect 10334 27134 10386 27186
rect 14590 27134 14642 27186
rect 14926 27134 14978 27186
rect 16830 27134 16882 27186
rect 17950 27134 18002 27186
rect 18846 27134 18898 27186
rect 20078 27134 20130 27186
rect 21646 27134 21698 27186
rect 22094 27134 22146 27186
rect 22654 27134 22706 27186
rect 23550 27134 23602 27186
rect 25678 27134 25730 27186
rect 26574 27134 26626 27186
rect 27694 27134 27746 27186
rect 28142 27134 28194 27186
rect 31502 27134 31554 27186
rect 32286 27134 32338 27186
rect 35198 27134 35250 27186
rect 36094 27134 36146 27186
rect 39118 27134 39170 27186
rect 42254 27134 42306 27186
rect 44270 27134 44322 27186
rect 46398 27134 46450 27186
rect 47294 27134 47346 27186
rect 47854 27134 47906 27186
rect 48302 27134 48354 27186
rect 50766 27134 50818 27186
rect 52334 27134 52386 27186
rect 57934 27134 57986 27186
rect 2606 27022 2658 27074
rect 5742 27022 5794 27074
rect 6078 27022 6130 27074
rect 6302 27022 6354 27074
rect 7310 27022 7362 27074
rect 9886 27022 9938 27074
rect 10446 27022 10498 27074
rect 12350 27022 12402 27074
rect 12574 27022 12626 27074
rect 12910 27022 12962 27074
rect 14702 27022 14754 27074
rect 15374 27022 15426 27074
rect 16718 27022 16770 27074
rect 17166 27022 17218 27074
rect 18510 27022 18562 27074
rect 20190 27022 20242 27074
rect 20302 27022 20354 27074
rect 20862 27022 20914 27074
rect 23326 27022 23378 27074
rect 24334 27022 24386 27074
rect 24782 27022 24834 27074
rect 25006 27022 25058 27074
rect 26126 27022 26178 27074
rect 27022 27022 27074 27074
rect 28590 27022 28642 27074
rect 30158 27022 30210 27074
rect 30494 27022 30546 27074
rect 30942 27022 30994 27074
rect 31166 27022 31218 27074
rect 31390 27022 31442 27074
rect 38446 27022 38498 27074
rect 38782 27022 38834 27074
rect 40238 27022 40290 27074
rect 40686 27022 40738 27074
rect 41470 27022 41522 27074
rect 41694 27022 41746 27074
rect 43374 27022 43426 27074
rect 43710 27022 43762 27074
rect 49982 27022 50034 27074
rect 51550 27022 51602 27074
rect 51886 27022 51938 27074
rect 53678 27022 53730 27074
rect 54350 27022 54402 27074
rect 54910 27022 54962 27074
rect 56030 27022 56082 27074
rect 3502 26910 3554 26962
rect 4398 26910 4450 26962
rect 9326 26910 9378 26962
rect 10334 26910 10386 26962
rect 11118 26910 11170 26962
rect 11454 26910 11506 26962
rect 13806 26910 13858 26962
rect 14478 26910 14530 26962
rect 16942 26910 16994 26962
rect 19294 26910 19346 26962
rect 26574 26910 26626 26962
rect 30270 26910 30322 26962
rect 32398 26910 32450 26962
rect 32622 26910 32674 26962
rect 34414 26910 34466 26962
rect 37886 26910 37938 26962
rect 45838 26910 45890 26962
rect 46958 26910 47010 26962
rect 49422 26910 49474 26962
rect 55134 26910 55186 26962
rect 55694 26910 55746 26962
rect 2158 26798 2210 26850
rect 2942 26798 2994 26850
rect 3838 26798 3890 26850
rect 7198 26798 7250 26850
rect 8990 26798 9042 26850
rect 10110 26798 10162 26850
rect 12798 26798 12850 26850
rect 15934 26798 15986 26850
rect 16606 26798 16658 26850
rect 19966 26798 20018 26850
rect 24558 26798 24610 26850
rect 31614 26798 31666 26850
rect 33182 26798 33234 26850
rect 35758 26798 35810 26850
rect 36542 26798 36594 26850
rect 37550 26798 37602 26850
rect 38558 26798 38610 26850
rect 45502 26798 45554 26850
rect 47182 26798 47234 26850
rect 47406 26798 47458 26850
rect 49086 26798 49138 26850
rect 50094 26798 50146 26850
rect 50318 26798 50370 26850
rect 57150 26798 57202 26850
rect 57486 26798 57538 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 2494 26462 2546 26514
rect 3502 26462 3554 26514
rect 3838 26462 3890 26514
rect 7870 26462 7922 26514
rect 9662 26462 9714 26514
rect 10894 26462 10946 26514
rect 12798 26462 12850 26514
rect 12910 26462 12962 26514
rect 14702 26462 14754 26514
rect 16830 26462 16882 26514
rect 17838 26462 17890 26514
rect 19294 26462 19346 26514
rect 25902 26462 25954 26514
rect 27134 26462 27186 26514
rect 28254 26462 28306 26514
rect 34750 26462 34802 26514
rect 35870 26462 35922 26514
rect 39118 26462 39170 26514
rect 40238 26462 40290 26514
rect 43710 26462 43762 26514
rect 44046 26462 44098 26514
rect 44830 26462 44882 26514
rect 46622 26462 46674 26514
rect 49870 26462 49922 26514
rect 50766 26462 50818 26514
rect 52110 26462 52162 26514
rect 52782 26462 52834 26514
rect 4398 26350 4450 26402
rect 4734 26350 4786 26402
rect 5406 26350 5458 26402
rect 7086 26350 7138 26402
rect 9886 26350 9938 26402
rect 10558 26350 10610 26402
rect 13022 26350 13074 26402
rect 13134 26350 13186 26402
rect 13358 26350 13410 26402
rect 14590 26350 14642 26402
rect 15486 26350 15538 26402
rect 15598 26350 15650 26402
rect 20414 26350 20466 26402
rect 22206 26350 22258 26402
rect 23550 26350 23602 26402
rect 29486 26350 29538 26402
rect 31726 26350 31778 26402
rect 32174 26350 32226 26402
rect 34414 26350 34466 26402
rect 35422 26350 35474 26402
rect 37998 26350 38050 26402
rect 39342 26350 39394 26402
rect 41582 26350 41634 26402
rect 42702 26350 42754 26402
rect 43822 26350 43874 26402
rect 44270 26350 44322 26402
rect 45054 26350 45106 26402
rect 45166 26350 45218 26402
rect 47742 26350 47794 26402
rect 50094 26350 50146 26402
rect 6750 26238 6802 26290
rect 7198 26238 7250 26290
rect 8430 26238 8482 26290
rect 9998 26238 10050 26290
rect 10894 26238 10946 26290
rect 11118 26238 11170 26290
rect 16270 26238 16322 26290
rect 16718 26238 16770 26290
rect 16942 26238 16994 26290
rect 17614 26238 17666 26290
rect 17950 26238 18002 26290
rect 19182 26238 19234 26290
rect 19406 26238 19458 26290
rect 20302 26238 20354 26290
rect 22654 26238 22706 26290
rect 24222 26238 24274 26290
rect 25678 26238 25730 26290
rect 25902 26238 25954 26290
rect 26238 26238 26290 26290
rect 28590 26238 28642 26290
rect 31278 26238 31330 26290
rect 32062 26238 32114 26290
rect 34638 26238 34690 26290
rect 34862 26238 34914 26290
rect 35646 26238 35698 26290
rect 36094 26238 36146 26290
rect 36430 26238 36482 26290
rect 37438 26238 37490 26290
rect 37774 26238 37826 26290
rect 38222 26238 38274 26290
rect 38670 26238 38722 26290
rect 40014 26238 40066 26290
rect 40462 26238 40514 26290
rect 40686 26238 40738 26290
rect 41806 26238 41858 26290
rect 42814 26238 42866 26290
rect 43150 26238 43202 26290
rect 46846 26238 46898 26290
rect 48078 26238 48130 26290
rect 49758 26238 49810 26290
rect 50318 26238 50370 26290
rect 52894 26238 52946 26290
rect 54014 26238 54066 26290
rect 54910 26238 54962 26290
rect 2158 26126 2210 26178
rect 2942 26126 2994 26178
rect 5854 26126 5906 26178
rect 6302 26126 6354 26178
rect 6862 26126 6914 26178
rect 11790 26126 11842 26178
rect 12238 26126 12290 26178
rect 14478 26126 14530 26178
rect 18958 26126 19010 26178
rect 24894 26126 24946 26178
rect 27694 26126 27746 26178
rect 29038 26126 29090 26178
rect 30046 26126 30098 26178
rect 31726 26126 31778 26178
rect 33518 26126 33570 26178
rect 36878 26126 36930 26178
rect 37886 26126 37938 26178
rect 39230 26126 39282 26178
rect 40798 26126 40850 26178
rect 45614 26126 45666 26178
rect 46062 26126 46114 26178
rect 48526 26126 48578 26178
rect 51214 26126 51266 26178
rect 51662 26126 51714 26178
rect 53454 26126 53506 26178
rect 56030 26126 56082 26178
rect 56590 26126 56642 26178
rect 58046 26126 58098 26178
rect 5182 26014 5234 26066
rect 5854 26014 5906 26066
rect 8654 26014 8706 26066
rect 8990 26014 9042 26066
rect 15486 26014 15538 26066
rect 18510 26014 18562 26066
rect 18734 26014 18786 26066
rect 27470 26014 27522 26066
rect 42142 26014 42194 26066
rect 43038 26014 43090 26066
rect 51102 26014 51154 26066
rect 51774 26014 51826 26066
rect 52782 26014 52834 26066
rect 57486 26014 57538 26066
rect 57822 26014 57874 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 3614 25678 3666 25730
rect 5182 25678 5234 25730
rect 7198 25678 7250 25730
rect 19854 25678 19906 25730
rect 21534 25678 21586 25730
rect 25454 25678 25506 25730
rect 27694 25678 27746 25730
rect 38334 25678 38386 25730
rect 40574 25678 40626 25730
rect 43934 25678 43986 25730
rect 46622 25678 46674 25730
rect 49198 25678 49250 25730
rect 51662 25678 51714 25730
rect 51998 25678 52050 25730
rect 2270 25566 2322 25618
rect 4958 25566 5010 25618
rect 7310 25566 7362 25618
rect 10110 25566 10162 25618
rect 12574 25566 12626 25618
rect 12910 25566 12962 25618
rect 14478 25566 14530 25618
rect 16942 25566 16994 25618
rect 17614 25566 17666 25618
rect 18398 25566 18450 25618
rect 19518 25566 19570 25618
rect 22654 25566 22706 25618
rect 24334 25566 24386 25618
rect 32062 25566 32114 25618
rect 34526 25566 34578 25618
rect 38782 25566 38834 25618
rect 41470 25566 41522 25618
rect 41918 25566 41970 25618
rect 44494 25566 44546 25618
rect 45614 25566 45666 25618
rect 51102 25566 51154 25618
rect 52334 25566 52386 25618
rect 54574 25566 54626 25618
rect 1934 25454 1986 25506
rect 6862 25454 6914 25506
rect 7198 25454 7250 25506
rect 7982 25454 8034 25506
rect 8430 25454 8482 25506
rect 11454 25454 11506 25506
rect 11566 25454 11618 25506
rect 14366 25454 14418 25506
rect 15262 25454 15314 25506
rect 19742 25454 19794 25506
rect 20078 25454 20130 25506
rect 20862 25454 20914 25506
rect 23438 25454 23490 25506
rect 24446 25454 24498 25506
rect 24782 25454 24834 25506
rect 31278 25454 31330 25506
rect 31950 25454 32002 25506
rect 34414 25454 34466 25506
rect 34862 25454 34914 25506
rect 35086 25454 35138 25506
rect 35870 25454 35922 25506
rect 36430 25454 36482 25506
rect 37774 25454 37826 25506
rect 37886 25454 37938 25506
rect 39566 25454 39618 25506
rect 40126 25454 40178 25506
rect 40798 25454 40850 25506
rect 42590 25454 42642 25506
rect 45726 25454 45778 25506
rect 46622 25454 46674 25506
rect 48078 25454 48130 25506
rect 49982 25454 50034 25506
rect 51214 25454 51266 25506
rect 53678 25454 53730 25506
rect 55246 25454 55298 25506
rect 56590 25454 56642 25506
rect 57934 25454 57986 25506
rect 2830 25342 2882 25394
rect 9998 25342 10050 25394
rect 14030 25342 14082 25394
rect 15038 25342 15090 25394
rect 17502 25342 17554 25394
rect 17726 25342 17778 25394
rect 19406 25342 19458 25394
rect 22094 25342 22146 25394
rect 23102 25342 23154 25394
rect 23214 25342 23266 25394
rect 23662 25342 23714 25394
rect 25566 25342 25618 25394
rect 26014 25342 26066 25394
rect 26238 25342 26290 25394
rect 26350 25342 26402 25394
rect 27694 25342 27746 25394
rect 27806 25342 27858 25394
rect 30942 25342 30994 25394
rect 31390 25342 31442 25394
rect 32286 25342 32338 25394
rect 33742 25342 33794 25394
rect 35534 25342 35586 25394
rect 36654 25342 36706 25394
rect 36766 25342 36818 25394
rect 37662 25342 37714 25394
rect 40350 25342 40402 25394
rect 41022 25342 41074 25394
rect 42926 25342 42978 25394
rect 3278 25230 3330 25282
rect 3726 25230 3778 25282
rect 4174 25230 4226 25282
rect 4622 25230 4674 25282
rect 5742 25230 5794 25282
rect 6078 25230 6130 25282
rect 9438 25230 9490 25282
rect 10222 25230 10274 25282
rect 10446 25230 10498 25282
rect 11230 25230 11282 25282
rect 11678 25230 11730 25282
rect 13694 25230 13746 25282
rect 13918 25230 13970 25282
rect 15486 25230 15538 25282
rect 15598 25230 15650 25282
rect 16046 25230 16098 25282
rect 16382 25230 16434 25282
rect 18958 25230 19010 25282
rect 21646 25230 21698 25282
rect 21870 25230 21922 25282
rect 24222 25230 24274 25282
rect 25454 25230 25506 25282
rect 26798 25230 26850 25282
rect 28254 25230 28306 25282
rect 28814 25230 28866 25282
rect 29486 25230 29538 25282
rect 29934 25230 29986 25282
rect 31166 25230 31218 25282
rect 32734 25230 32786 25282
rect 33406 25230 33458 25282
rect 34638 25230 34690 25282
rect 35758 25230 35810 25282
rect 39454 25230 39506 25282
rect 40462 25230 40514 25282
rect 42814 25230 42866 25282
rect 43038 25230 43090 25282
rect 43150 25230 43202 25282
rect 43934 25230 43986 25282
rect 44046 25286 44098 25338
rect 45502 25342 45554 25394
rect 46062 25342 46114 25394
rect 46958 25342 47010 25394
rect 48974 25342 49026 25394
rect 49086 25342 49138 25394
rect 49758 25342 49810 25394
rect 50766 25342 50818 25394
rect 53790 25342 53842 25394
rect 47406 25230 47458 25282
rect 48190 25230 48242 25282
rect 48414 25230 48466 25282
rect 51886 25230 51938 25282
rect 57710 25230 57762 25282
rect 58606 25230 58658 25282
rect 59614 25230 59666 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 1934 24894 1986 24946
rect 12126 24894 12178 24946
rect 16942 24894 16994 24946
rect 19294 24894 19346 24946
rect 21198 24894 21250 24946
rect 27022 24894 27074 24946
rect 28142 24894 28194 24946
rect 32510 24894 32562 24946
rect 32958 24894 33010 24946
rect 33966 24894 34018 24946
rect 37326 24894 37378 24946
rect 38334 24894 38386 24946
rect 38782 24894 38834 24946
rect 39454 24894 39506 24946
rect 41582 24894 41634 24946
rect 45278 24894 45330 24946
rect 52558 24894 52610 24946
rect 53454 24894 53506 24946
rect 54014 24894 54066 24946
rect 54798 24894 54850 24946
rect 56142 24894 56194 24946
rect 56590 24894 56642 24946
rect 2830 24782 2882 24834
rect 9886 24782 9938 24834
rect 18174 24782 18226 24834
rect 21086 24782 21138 24834
rect 24334 24782 24386 24834
rect 26014 24782 26066 24834
rect 27246 24782 27298 24834
rect 29262 24782 29314 24834
rect 34414 24782 34466 24834
rect 35086 24782 35138 24834
rect 35982 24782 36034 24834
rect 42814 24782 42866 24834
rect 45166 24782 45218 24834
rect 45838 24782 45890 24834
rect 47070 24782 47122 24834
rect 50878 24782 50930 24834
rect 52446 24782 52498 24834
rect 55134 24782 55186 24834
rect 55806 24782 55858 24834
rect 57486 24782 57538 24834
rect 57598 24782 57650 24834
rect 4062 24670 4114 24722
rect 4286 24670 4338 24722
rect 5854 24670 5906 24722
rect 6974 24670 7026 24722
rect 8430 24670 8482 24722
rect 10446 24670 10498 24722
rect 10782 24670 10834 24722
rect 12014 24670 12066 24722
rect 12350 24670 12402 24722
rect 12798 24670 12850 24722
rect 13470 24670 13522 24722
rect 14030 24670 14082 24722
rect 17838 24670 17890 24722
rect 19070 24670 19122 24722
rect 20190 24670 20242 24722
rect 21982 24670 22034 24722
rect 23998 24670 24050 24722
rect 25790 24670 25842 24722
rect 26910 24670 26962 24722
rect 2382 24558 2434 24610
rect 6638 24558 6690 24610
rect 9102 24558 9154 24610
rect 10110 24558 10162 24610
rect 11566 24558 11618 24610
rect 14814 24558 14866 24610
rect 15150 24558 15202 24610
rect 15598 24558 15650 24610
rect 16046 24558 16098 24610
rect 16494 24558 16546 24610
rect 18734 24558 18786 24610
rect 3054 24446 3106 24498
rect 3390 24446 3442 24498
rect 12462 24446 12514 24498
rect 18398 24446 18450 24498
rect 27358 24670 27410 24722
rect 28030 24670 28082 24722
rect 28254 24670 28306 24722
rect 28590 24670 28642 24722
rect 37214 24670 37266 24722
rect 37550 24670 37602 24722
rect 37774 24670 37826 24722
rect 39902 24670 39954 24722
rect 43150 24670 43202 24722
rect 44158 24670 44210 24722
rect 45054 24670 45106 24722
rect 45614 24670 45666 24722
rect 46734 24670 46786 24722
rect 47518 24670 47570 24722
rect 47966 24670 48018 24722
rect 49534 24670 49586 24722
rect 49870 24670 49922 24722
rect 50430 24670 50482 24722
rect 51102 24670 51154 24722
rect 51214 24670 51266 24722
rect 52782 24670 52834 24722
rect 53006 24670 53058 24722
rect 53566 24670 53618 24722
rect 53790 24670 53842 24722
rect 54126 24670 54178 24722
rect 57710 24670 57762 24722
rect 58046 24670 58098 24722
rect 19630 24558 19682 24610
rect 24894 24558 24946 24610
rect 29150 24558 29202 24610
rect 29934 24558 29986 24610
rect 30382 24558 30434 24610
rect 30830 24558 30882 24610
rect 31614 24558 31666 24610
rect 33518 24558 33570 24610
rect 35534 24558 35586 24610
rect 36430 24558 36482 24610
rect 37662 24558 37714 24610
rect 40798 24558 40850 24610
rect 41918 24558 41970 24610
rect 46958 24558 47010 24610
rect 48638 24558 48690 24610
rect 19630 24446 19682 24498
rect 29486 24446 29538 24498
rect 35982 24446 36034 24498
rect 36430 24446 36482 24498
rect 40126 24446 40178 24498
rect 40238 24446 40290 24498
rect 48414 24446 48466 24498
rect 48638 24446 48690 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 3166 24110 3218 24162
rect 7982 24110 8034 24162
rect 11566 24110 11618 24162
rect 11790 24110 11842 24162
rect 16382 24110 16434 24162
rect 16942 24110 16994 24162
rect 18398 24110 18450 24162
rect 28590 24110 28642 24162
rect 31166 24110 31218 24162
rect 37662 24110 37714 24162
rect 38334 24110 38386 24162
rect 41134 24110 41186 24162
rect 42030 24110 42082 24162
rect 49310 24110 49362 24162
rect 50766 24110 50818 24162
rect 4510 23998 4562 24050
rect 5966 23998 6018 24050
rect 6974 23998 7026 24050
rect 7870 23998 7922 24050
rect 8878 23998 8930 24050
rect 12014 23998 12066 24050
rect 12350 23998 12402 24050
rect 13806 23998 13858 24050
rect 16606 23998 16658 24050
rect 21646 23998 21698 24050
rect 24110 23998 24162 24050
rect 26798 23998 26850 24050
rect 33070 23998 33122 24050
rect 36206 23998 36258 24050
rect 37438 23998 37490 24050
rect 40238 23998 40290 24050
rect 40686 23998 40738 24050
rect 41246 23998 41298 24050
rect 41694 23998 41746 24050
rect 42030 23998 42082 24050
rect 42702 23998 42754 24050
rect 43598 23998 43650 24050
rect 44494 23998 44546 24050
rect 45614 23998 45666 24050
rect 47182 23998 47234 24050
rect 48526 23998 48578 24050
rect 52334 23998 52386 24050
rect 54462 23998 54514 24050
rect 55918 23998 55970 24050
rect 57150 23998 57202 24050
rect 57822 23998 57874 24050
rect 2158 23886 2210 23938
rect 2494 23886 2546 23938
rect 4846 23886 4898 23938
rect 6526 23886 6578 23938
rect 2942 23830 2994 23882
rect 6750 23886 6802 23938
rect 7198 23886 7250 23938
rect 7422 23886 7474 23938
rect 9662 23886 9714 23938
rect 10222 23886 10274 23938
rect 14702 23886 14754 23938
rect 15374 23886 15426 23938
rect 2270 23774 2322 23826
rect 16494 23886 16546 23938
rect 17166 23886 17218 23938
rect 18510 23886 18562 23938
rect 19294 23886 19346 23938
rect 19630 23886 19682 23938
rect 19742 23886 19794 23938
rect 20526 23886 20578 23938
rect 20862 23886 20914 23938
rect 23214 23886 23266 23938
rect 24222 23886 24274 23938
rect 24782 23886 24834 23938
rect 25342 23886 25394 23938
rect 25454 23886 25506 23938
rect 27694 23886 27746 23938
rect 30942 23886 30994 23938
rect 31502 23886 31554 23938
rect 33854 23886 33906 23938
rect 38894 23886 38946 23938
rect 44046 23886 44098 23938
rect 45726 23886 45778 23938
rect 46174 23886 46226 23938
rect 48190 23886 48242 23938
rect 48750 23886 48802 23938
rect 49982 23886 50034 23938
rect 51550 23886 51602 23938
rect 53454 23886 53506 23938
rect 55246 23886 55298 23938
rect 55582 23886 55634 23938
rect 56590 23886 56642 23938
rect 9774 23774 9826 23826
rect 13806 23774 13858 23826
rect 14030 23774 14082 23826
rect 15710 23774 15762 23826
rect 17838 23774 17890 23826
rect 18062 23774 18114 23826
rect 20078 23774 20130 23826
rect 20750 23774 20802 23826
rect 22318 23774 22370 23826
rect 22878 23774 22930 23826
rect 23774 23774 23826 23826
rect 27246 23774 27298 23826
rect 28030 23774 28082 23826
rect 28702 23774 28754 23826
rect 29934 23774 29986 23826
rect 33294 23774 33346 23826
rect 33518 23774 33570 23826
rect 34302 23774 34354 23826
rect 34638 23774 34690 23826
rect 35646 23774 35698 23826
rect 37886 23774 37938 23826
rect 39342 23774 39394 23826
rect 47294 23774 47346 23826
rect 49422 23774 49474 23826
rect 50542 23774 50594 23826
rect 51886 23774 51938 23826
rect 54014 23774 54066 23826
rect 57038 23830 57090 23882
rect 3502 23662 3554 23714
rect 7422 23662 7474 23714
rect 7758 23662 7810 23714
rect 10446 23662 10498 23714
rect 10558 23662 10610 23714
rect 12238 23662 12290 23714
rect 12462 23662 12514 23714
rect 14926 23662 14978 23714
rect 15598 23662 15650 23714
rect 18286 23662 18338 23714
rect 19294 23662 19346 23714
rect 22430 23662 22482 23714
rect 27918 23662 27970 23714
rect 29486 23662 29538 23714
rect 32510 23662 32562 23714
rect 33630 23662 33682 23714
rect 34526 23662 34578 23714
rect 35310 23662 35362 23714
rect 36542 23662 36594 23714
rect 38334 23662 38386 23714
rect 39790 23662 39842 23714
rect 43150 23662 43202 23714
rect 45502 23662 45554 23714
rect 46846 23662 46898 23714
rect 47070 23662 47122 23714
rect 48414 23662 48466 23714
rect 48638 23662 48690 23714
rect 49646 23662 49698 23714
rect 50654 23662 50706 23714
rect 57150 23662 57202 23714
rect 57374 23662 57426 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 5742 23326 5794 23378
rect 8206 23326 8258 23378
rect 8542 23326 8594 23378
rect 11342 23326 11394 23378
rect 17838 23326 17890 23378
rect 20862 23326 20914 23378
rect 23214 23326 23266 23378
rect 25006 23326 25058 23378
rect 28702 23326 28754 23378
rect 29486 23326 29538 23378
rect 32286 23326 32338 23378
rect 32622 23326 32674 23378
rect 33966 23326 34018 23378
rect 36206 23326 36258 23378
rect 36318 23326 36370 23378
rect 39006 23326 39058 23378
rect 40014 23326 40066 23378
rect 40910 23326 40962 23378
rect 42478 23326 42530 23378
rect 44718 23326 44770 23378
rect 45838 23326 45890 23378
rect 46622 23326 46674 23378
rect 47294 23326 47346 23378
rect 48638 23326 48690 23378
rect 51550 23326 51602 23378
rect 54238 23326 54290 23378
rect 55246 23326 55298 23378
rect 57486 23326 57538 23378
rect 6190 23214 6242 23266
rect 10670 23214 10722 23266
rect 13022 23214 13074 23266
rect 14590 23214 14642 23266
rect 15262 23214 15314 23266
rect 15710 23214 15762 23266
rect 18062 23214 18114 23266
rect 18286 23214 18338 23266
rect 19518 23214 19570 23266
rect 20414 23214 20466 23266
rect 20638 23214 20690 23266
rect 21758 23214 21810 23266
rect 25678 23214 25730 23266
rect 27806 23214 27858 23266
rect 31838 23214 31890 23266
rect 32398 23214 32450 23266
rect 33518 23214 33570 23266
rect 40350 23214 40402 23266
rect 41694 23214 41746 23266
rect 41918 23214 41970 23266
rect 44494 23214 44546 23266
rect 45278 23214 45330 23266
rect 48190 23214 48242 23266
rect 3054 23102 3106 23154
rect 4062 23102 4114 23154
rect 4398 23102 4450 23154
rect 5070 23102 5122 23154
rect 7534 23102 7586 23154
rect 10446 23102 10498 23154
rect 11790 23102 11842 23154
rect 13582 23102 13634 23154
rect 14814 23102 14866 23154
rect 17726 23102 17778 23154
rect 21198 23102 21250 23154
rect 21982 23102 22034 23154
rect 22206 23102 22258 23154
rect 23662 23102 23714 23154
rect 26238 23102 26290 23154
rect 27022 23102 27074 23154
rect 27918 23102 27970 23154
rect 29038 23102 29090 23154
rect 29934 23102 29986 23154
rect 31166 23102 31218 23154
rect 31726 23102 31778 23154
rect 32958 23102 33010 23154
rect 34526 23102 34578 23154
rect 34750 23102 34802 23154
rect 35086 23102 35138 23154
rect 35870 23102 35922 23154
rect 36094 23102 36146 23154
rect 36542 23102 36594 23154
rect 37550 23102 37602 23154
rect 37886 23102 37938 23154
rect 38110 23102 38162 23154
rect 39790 23102 39842 23154
rect 40126 23102 40178 23154
rect 43150 23102 43202 23154
rect 43486 23102 43538 23154
rect 43710 23102 43762 23154
rect 44382 23102 44434 23154
rect 45054 23102 45106 23154
rect 49534 23214 49586 23266
rect 49758 23214 49810 23266
rect 50654 23214 50706 23266
rect 52446 23214 52498 23266
rect 54462 23214 54514 23266
rect 57822 23214 57874 23266
rect 45390 23102 45442 23154
rect 46846 23102 46898 23154
rect 49310 23102 49362 23154
rect 50990 23102 51042 23154
rect 52782 23102 52834 23154
rect 53902 23102 53954 23154
rect 54574 23102 54626 23154
rect 55134 23102 55186 23154
rect 55918 23102 55970 23154
rect 56478 23102 56530 23154
rect 1822 22990 1874 23042
rect 2270 22990 2322 23042
rect 8990 22990 9042 23042
rect 16494 22990 16546 23042
rect 16942 22990 16994 23042
rect 19070 22990 19122 23042
rect 22094 22990 22146 23042
rect 22766 22990 22818 23042
rect 24222 22990 24274 23042
rect 27470 22990 27522 23042
rect 34638 22990 34690 23042
rect 36990 22990 37042 23042
rect 37662 22990 37714 23042
rect 38558 22990 38610 23042
rect 41582 22990 41634 23042
rect 43262 22990 43314 23042
rect 47742 22990 47794 23042
rect 51886 22990 51938 23042
rect 53230 22990 53282 23042
rect 25790 22878 25842 22930
rect 26014 22878 26066 22930
rect 46510 22878 46562 22930
rect 47518 22878 47570 22930
rect 48638 22878 48690 22930
rect 49646 22878 49698 22930
rect 49982 22878 50034 22930
rect 55246 22878 55298 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 9214 22542 9266 22594
rect 10782 22542 10834 22594
rect 16046 22542 16098 22594
rect 26798 22542 26850 22594
rect 29934 22542 29986 22594
rect 34526 22542 34578 22594
rect 35758 22542 35810 22594
rect 42814 22542 42866 22594
rect 46958 22542 47010 22594
rect 51326 22542 51378 22594
rect 56590 22542 56642 22594
rect 1934 22430 1986 22482
rect 3726 22430 3778 22482
rect 7534 22430 7586 22482
rect 8542 22430 8594 22482
rect 11790 22430 11842 22482
rect 12574 22430 12626 22482
rect 13022 22430 13074 22482
rect 13806 22430 13858 22482
rect 18734 22430 18786 22482
rect 18958 22430 19010 22482
rect 21646 22430 21698 22482
rect 25566 22430 25618 22482
rect 29598 22430 29650 22482
rect 31390 22430 31442 22482
rect 31950 22430 32002 22482
rect 37998 22430 38050 22482
rect 39006 22430 39058 22482
rect 40126 22430 40178 22482
rect 41022 22430 41074 22482
rect 41470 22430 41522 22482
rect 47294 22430 47346 22482
rect 48862 22430 48914 22482
rect 55806 22430 55858 22482
rect 2830 22318 2882 22370
rect 3614 22318 3666 22370
rect 4286 22318 4338 22370
rect 4958 22318 5010 22370
rect 6302 22318 6354 22370
rect 6638 22318 6690 22370
rect 6974 22318 7026 22370
rect 7422 22318 7474 22370
rect 9326 22318 9378 22370
rect 10110 22318 10162 22370
rect 14254 22318 14306 22370
rect 15374 22318 15426 22370
rect 16606 22318 16658 22370
rect 16942 22318 16994 22370
rect 18174 22318 18226 22370
rect 18622 22318 18674 22370
rect 19182 22318 19234 22370
rect 20078 22318 20130 22370
rect 20638 22318 20690 22370
rect 22878 22318 22930 22370
rect 25678 22318 25730 22370
rect 26350 22318 26402 22370
rect 27470 22318 27522 22370
rect 28590 22318 28642 22370
rect 31838 22318 31890 22370
rect 32286 22318 32338 22370
rect 35870 22318 35922 22370
rect 36430 22318 36482 22370
rect 36542 22318 36594 22370
rect 40014 22318 40066 22370
rect 42478 22318 42530 22370
rect 43038 22318 43090 22370
rect 47070 22318 47122 22370
rect 47518 22318 47570 22370
rect 48974 22318 49026 22370
rect 49758 22318 49810 22370
rect 50206 22318 50258 22370
rect 51438 22318 51490 22370
rect 52110 22318 52162 22370
rect 52334 22318 52386 22370
rect 55022 22318 55074 22370
rect 55246 22318 55298 22370
rect 55470 22318 55522 22370
rect 55694 22318 55746 22370
rect 57598 22318 57650 22370
rect 3838 22206 3890 22258
rect 5854 22206 5906 22258
rect 6414 22206 6466 22258
rect 9214 22206 9266 22258
rect 10670 22206 10722 22258
rect 14590 22206 14642 22258
rect 15934 22206 15986 22258
rect 21982 22206 22034 22258
rect 22766 22206 22818 22258
rect 23550 22206 23602 22258
rect 28254 22206 28306 22258
rect 28478 22206 28530 22258
rect 30158 22206 30210 22258
rect 30606 22206 30658 22258
rect 32510 22206 32562 22258
rect 33518 22206 33570 22258
rect 34302 22206 34354 22258
rect 36654 22206 36706 22258
rect 37886 22206 37938 22258
rect 37998 22206 38050 22258
rect 40462 22206 40514 22258
rect 42254 22206 42306 22258
rect 44046 22206 44098 22258
rect 45838 22206 45890 22258
rect 46174 22206 46226 22258
rect 46398 22206 46450 22258
rect 48414 22206 48466 22258
rect 48638 22206 48690 22258
rect 50766 22206 50818 22258
rect 51998 22206 52050 22258
rect 53454 22206 53506 22258
rect 56926 22206 56978 22258
rect 57822 22206 57874 22258
rect 7646 22094 7698 22146
rect 8094 22094 8146 22146
rect 10446 22094 10498 22146
rect 11230 22094 11282 22146
rect 15150 22094 15202 22146
rect 16046 22094 16098 22146
rect 16830 22094 16882 22146
rect 17838 22094 17890 22146
rect 19294 22094 19346 22146
rect 23886 22094 23938 22146
rect 32062 22094 32114 22146
rect 33182 22094 33234 22146
rect 34414 22094 34466 22146
rect 34974 22094 35026 22146
rect 36206 22094 36258 22146
rect 38110 22094 38162 22146
rect 38334 22094 38386 22146
rect 39454 22094 39506 22146
rect 40238 22094 40290 22146
rect 43150 22094 43202 22146
rect 43710 22094 43762 22146
rect 44494 22094 44546 22146
rect 46062 22094 46114 22146
rect 49758 22094 49810 22146
rect 51774 22094 51826 22146
rect 53790 22094 53842 22146
rect 54238 22094 54290 22146
rect 55918 22094 55970 22146
rect 56702 22094 56754 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 2158 21758 2210 21810
rect 3838 21758 3890 21810
rect 5518 21758 5570 21810
rect 6638 21758 6690 21810
rect 7982 21758 8034 21810
rect 10558 21758 10610 21810
rect 12686 21758 12738 21810
rect 16830 21758 16882 21810
rect 17838 21758 17890 21810
rect 19182 21758 19234 21810
rect 20078 21758 20130 21810
rect 21646 21758 21698 21810
rect 22542 21758 22594 21810
rect 26014 21758 26066 21810
rect 27694 21758 27746 21810
rect 30830 21758 30882 21810
rect 35422 21758 35474 21810
rect 36654 21758 36706 21810
rect 37662 21758 37714 21810
rect 40126 21758 40178 21810
rect 41470 21758 41522 21810
rect 41918 21758 41970 21810
rect 47518 21758 47570 21810
rect 49422 21758 49474 21810
rect 50542 21758 50594 21810
rect 54350 21758 54402 21810
rect 57486 21758 57538 21810
rect 2830 21646 2882 21698
rect 3278 21646 3330 21698
rect 4958 21646 5010 21698
rect 10110 21646 10162 21698
rect 12238 21646 12290 21698
rect 12910 21646 12962 21698
rect 15822 21646 15874 21698
rect 16158 21646 16210 21698
rect 17054 21646 17106 21698
rect 17950 21646 18002 21698
rect 18062 21646 18114 21698
rect 18174 21646 18226 21698
rect 20862 21646 20914 21698
rect 22094 21646 22146 21698
rect 22318 21646 22370 21698
rect 23438 21646 23490 21698
rect 23662 21646 23714 21698
rect 26686 21646 26738 21698
rect 27806 21646 27858 21698
rect 30046 21646 30098 21698
rect 32510 21646 32562 21698
rect 32846 21646 32898 21698
rect 34078 21646 34130 21698
rect 36206 21646 36258 21698
rect 42478 21646 42530 21698
rect 44942 21646 44994 21698
rect 45838 21646 45890 21698
rect 47742 21646 47794 21698
rect 47966 21646 48018 21698
rect 51662 21646 51714 21698
rect 55582 21646 55634 21698
rect 56366 21646 56418 21698
rect 4510 21534 4562 21586
rect 5406 21534 5458 21586
rect 6414 21534 6466 21586
rect 7870 21534 7922 21586
rect 8094 21534 8146 21586
rect 10334 21534 10386 21586
rect 11118 21534 11170 21586
rect 12126 21534 12178 21586
rect 13022 21534 13074 21586
rect 14702 21534 14754 21586
rect 14926 21534 14978 21586
rect 15374 21534 15426 21586
rect 16718 21534 16770 21586
rect 17726 21534 17778 21586
rect 19406 21534 19458 21586
rect 20526 21534 20578 21586
rect 21310 21534 21362 21586
rect 21534 21534 21586 21586
rect 22654 21534 22706 21586
rect 23326 21534 23378 21586
rect 24446 21534 24498 21586
rect 26574 21534 26626 21586
rect 27022 21534 27074 21586
rect 27582 21534 27634 21586
rect 28366 21534 28418 21586
rect 28926 21534 28978 21586
rect 30270 21534 30322 21586
rect 31278 21534 31330 21586
rect 33966 21534 34018 21586
rect 34526 21534 34578 21586
rect 35422 21534 35474 21586
rect 35982 21534 36034 21586
rect 40014 21534 40066 21586
rect 40350 21534 40402 21586
rect 40574 21534 40626 21586
rect 42702 21534 42754 21586
rect 44158 21534 44210 21586
rect 46398 21534 46450 21586
rect 47406 21534 47458 21586
rect 47518 21534 47570 21586
rect 50318 21534 50370 21586
rect 50542 21534 50594 21586
rect 50878 21534 50930 21586
rect 51886 21534 51938 21586
rect 52222 21534 52274 21586
rect 53790 21534 53842 21586
rect 55246 21534 55298 21586
rect 56702 21534 56754 21586
rect 57710 21534 57762 21586
rect 3502 21422 3554 21474
rect 7646 21422 7698 21474
rect 9102 21422 9154 21474
rect 10558 21422 10610 21474
rect 14142 21422 14194 21474
rect 14814 21422 14866 21474
rect 19070 21422 19122 21474
rect 23998 21422 24050 21474
rect 24894 21422 24946 21474
rect 26910 21422 26962 21474
rect 28030 21422 28082 21474
rect 31950 21422 32002 21474
rect 34190 21422 34242 21474
rect 37102 21422 37154 21474
rect 38110 21422 38162 21474
rect 38558 21422 38610 21474
rect 39006 21422 39058 21474
rect 39454 21422 39506 21474
rect 48414 21422 48466 21474
rect 51774 21422 51826 21474
rect 52670 21422 52722 21474
rect 53342 21422 53394 21474
rect 54686 21422 54738 21474
rect 7198 21310 7250 21362
rect 7422 21310 7474 21362
rect 14254 21310 14306 21362
rect 14478 21310 14530 21362
rect 21086 21310 21138 21362
rect 29150 21310 29202 21362
rect 29486 21310 29538 21362
rect 35758 21310 35810 21362
rect 37326 21310 37378 21362
rect 37886 21310 37938 21362
rect 38558 21310 38610 21362
rect 41470 21310 41522 21362
rect 41918 21310 41970 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 18846 20974 18898 21026
rect 19854 20974 19906 21026
rect 20078 20974 20130 21026
rect 23102 20974 23154 21026
rect 23774 20974 23826 21026
rect 31950 20974 32002 21026
rect 32622 20974 32674 21026
rect 34302 20974 34354 21026
rect 34862 20974 34914 21026
rect 37662 20974 37714 21026
rect 40462 20974 40514 21026
rect 41470 20974 41522 21026
rect 41806 20974 41858 21026
rect 42478 20974 42530 21026
rect 46622 20974 46674 21026
rect 47742 20974 47794 21026
rect 47966 20974 48018 21026
rect 48638 20974 48690 21026
rect 48974 20974 49026 21026
rect 49422 20974 49474 21026
rect 1934 20862 1986 20914
rect 2382 20862 2434 20914
rect 2830 20862 2882 20914
rect 4174 20862 4226 20914
rect 6078 20862 6130 20914
rect 8318 20862 8370 20914
rect 12462 20862 12514 20914
rect 13582 20862 13634 20914
rect 14254 20862 14306 20914
rect 15374 20862 15426 20914
rect 15822 20862 15874 20914
rect 16494 20862 16546 20914
rect 18622 20862 18674 20914
rect 20638 20862 20690 20914
rect 24670 20862 24722 20914
rect 25342 20862 25394 20914
rect 26462 20862 26514 20914
rect 27582 20862 27634 20914
rect 29486 20862 29538 20914
rect 32286 20862 32338 20914
rect 32734 20862 32786 20914
rect 33070 20862 33122 20914
rect 34862 20862 34914 20914
rect 36654 20862 36706 20914
rect 38894 20862 38946 20914
rect 45390 20862 45442 20914
rect 48190 20862 48242 20914
rect 6302 20750 6354 20802
rect 6638 20750 6690 20802
rect 7646 20750 7698 20802
rect 8990 20750 9042 20802
rect 10334 20750 10386 20802
rect 12350 20750 12402 20802
rect 14590 20750 14642 20802
rect 16942 20750 16994 20802
rect 18174 20750 18226 20802
rect 20302 20750 20354 20802
rect 22878 20750 22930 20802
rect 23326 20750 23378 20802
rect 24334 20750 24386 20802
rect 25118 20750 25170 20802
rect 25566 20750 25618 20802
rect 27694 20750 27746 20802
rect 28142 20750 28194 20802
rect 30270 20750 30322 20802
rect 30830 20750 30882 20802
rect 33406 20750 33458 20802
rect 33854 20750 33906 20802
rect 35870 20750 35922 20802
rect 37774 20750 37826 20802
rect 38110 20750 38162 20802
rect 38334 20750 38386 20802
rect 40126 20750 40178 20802
rect 41246 20750 41298 20802
rect 42814 20750 42866 20802
rect 43038 20750 43090 20802
rect 4622 20638 4674 20690
rect 7534 20638 7586 20690
rect 12798 20638 12850 20690
rect 14254 20638 14306 20690
rect 14814 20638 14866 20690
rect 17726 20638 17778 20690
rect 19182 20638 19234 20690
rect 19518 20638 19570 20690
rect 25790 20638 25842 20690
rect 27134 20638 27186 20690
rect 28702 20638 28754 20690
rect 33182 20638 33234 20690
rect 37550 20638 37602 20690
rect 39902 20638 39954 20690
rect 43598 20638 43650 20690
rect 46622 20638 46674 20690
rect 46734 20638 46786 20690
rect 50430 20974 50482 21026
rect 57262 20974 57314 21026
rect 50878 20862 50930 20914
rect 53342 20862 53394 20914
rect 56590 20862 56642 20914
rect 57822 20862 57874 20914
rect 54014 20750 54066 20802
rect 55022 20750 55074 20802
rect 57374 20750 57426 20802
rect 47406 20638 47458 20690
rect 50318 20638 50370 20690
rect 51550 20638 51602 20690
rect 51886 20638 51938 20690
rect 54350 20638 54402 20690
rect 56030 20638 56082 20690
rect 3278 20526 3330 20578
rect 3726 20526 3778 20578
rect 5070 20526 5122 20578
rect 11566 20526 11618 20578
rect 12238 20526 12290 20578
rect 12574 20526 12626 20578
rect 14366 20526 14418 20578
rect 16382 20526 16434 20578
rect 16606 20526 16658 20578
rect 20526 20526 20578 20578
rect 20750 20526 20802 20578
rect 21870 20526 21922 20578
rect 22318 20526 22370 20578
rect 24558 20526 24610 20578
rect 30046 20526 30098 20578
rect 31838 20526 31890 20578
rect 33630 20526 33682 20578
rect 34302 20526 34354 20578
rect 35310 20526 35362 20578
rect 36206 20526 36258 20578
rect 39342 20526 39394 20578
rect 40350 20526 40402 20578
rect 43934 20526 43986 20578
rect 44382 20526 44434 20578
rect 45838 20526 45890 20578
rect 47630 20526 47682 20578
rect 48638 20526 48690 20578
rect 49086 20526 49138 20578
rect 49534 20526 49586 20578
rect 49982 20526 50034 20578
rect 50430 20526 50482 20578
rect 51774 20526 51826 20578
rect 52334 20526 52386 20578
rect 54238 20526 54290 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 3054 20190 3106 20242
rect 4286 20190 4338 20242
rect 12350 20190 12402 20242
rect 18510 20190 18562 20242
rect 20190 20190 20242 20242
rect 23662 20190 23714 20242
rect 26238 20190 26290 20242
rect 27358 20190 27410 20242
rect 29934 20190 29986 20242
rect 33630 20190 33682 20242
rect 35758 20190 35810 20242
rect 38446 20190 38498 20242
rect 39566 20190 39618 20242
rect 40126 20190 40178 20242
rect 44270 20190 44322 20242
rect 45838 20190 45890 20242
rect 48526 20190 48578 20242
rect 51550 20190 51602 20242
rect 53566 20190 53618 20242
rect 54574 20190 54626 20242
rect 55582 20190 55634 20242
rect 57822 20190 57874 20242
rect 2158 20078 2210 20130
rect 10670 20078 10722 20130
rect 12238 20078 12290 20130
rect 15038 20078 15090 20130
rect 16158 20078 16210 20130
rect 19854 20078 19906 20130
rect 22430 20078 22482 20130
rect 23774 20078 23826 20130
rect 24334 20078 24386 20130
rect 29038 20078 29090 20130
rect 32510 20078 32562 20130
rect 34078 20078 34130 20130
rect 34862 20078 34914 20130
rect 35198 20078 35250 20130
rect 36766 20078 36818 20130
rect 36990 20078 37042 20130
rect 41582 20078 41634 20130
rect 42814 20078 42866 20130
rect 43038 20078 43090 20130
rect 45278 20078 45330 20130
rect 48414 20078 48466 20130
rect 53006 20078 53058 20130
rect 56702 20078 56754 20130
rect 57486 20078 57538 20130
rect 3390 19966 3442 20018
rect 4510 19966 4562 20018
rect 4958 19966 5010 20018
rect 7310 19966 7362 20018
rect 8094 19966 8146 20018
rect 8430 19966 8482 20018
rect 9662 19966 9714 20018
rect 10446 19966 10498 20018
rect 11790 19966 11842 20018
rect 12462 19966 12514 20018
rect 14030 19966 14082 20018
rect 19070 19966 19122 20018
rect 19742 19966 19794 20018
rect 20974 19966 21026 20018
rect 23550 19966 23602 20018
rect 25902 19966 25954 20018
rect 26014 19966 26066 20018
rect 26238 19966 26290 20018
rect 26462 19966 26514 20018
rect 28142 19966 28194 20018
rect 29710 19966 29762 20018
rect 30158 19966 30210 20018
rect 30382 19966 30434 20018
rect 33854 19966 33906 20018
rect 36094 19966 36146 20018
rect 37550 19966 37602 20018
rect 39118 19966 39170 20018
rect 39342 19966 39394 20018
rect 41806 19966 41858 20018
rect 42030 19966 42082 20018
rect 44270 19966 44322 20018
rect 45166 19966 45218 20018
rect 46174 19966 46226 20018
rect 46734 19966 46786 20018
rect 47182 19966 47234 20018
rect 48302 19966 48354 20018
rect 48862 19966 48914 20018
rect 49758 19966 49810 20018
rect 50318 19966 50370 20018
rect 51886 19966 51938 20018
rect 52782 19966 52834 20018
rect 53230 19966 53282 20018
rect 53454 19966 53506 20018
rect 54350 19966 54402 20018
rect 55470 19966 55522 20018
rect 2606 19854 2658 19906
rect 4734 19854 4786 19906
rect 5742 19854 5794 19906
rect 6078 19854 6130 19906
rect 7198 19854 7250 19906
rect 7646 19854 7698 19906
rect 8990 19854 9042 19906
rect 10334 19854 10386 19906
rect 13694 19854 13746 19906
rect 13806 19854 13858 19906
rect 16606 19854 16658 19906
rect 17950 19854 18002 19906
rect 20526 19854 20578 19906
rect 21870 19854 21922 19906
rect 22990 19854 23042 19906
rect 26910 19854 26962 19906
rect 28590 19854 28642 19906
rect 30830 19854 30882 19906
rect 31278 19854 31330 19906
rect 31726 19854 31778 19906
rect 32958 19854 33010 19906
rect 37998 19854 38050 19906
rect 39230 19854 39282 19906
rect 40574 19854 40626 19906
rect 41694 19854 41746 19906
rect 43486 19854 43538 19906
rect 47406 19854 47458 19906
rect 50542 19854 50594 19906
rect 56590 19854 56642 19906
rect 22766 19742 22818 19794
rect 26910 19742 26962 19794
rect 27246 19742 27298 19794
rect 30494 19742 30546 19794
rect 30830 19742 30882 19794
rect 33518 19742 33570 19794
rect 37102 19742 37154 19794
rect 42702 19742 42754 19794
rect 47518 19742 47570 19794
rect 50654 19742 50706 19794
rect 55694 19742 55746 19794
rect 55918 19742 55970 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 5742 19406 5794 19458
rect 12350 19406 12402 19458
rect 12686 19406 12738 19458
rect 14254 19406 14306 19458
rect 15486 19406 15538 19458
rect 21646 19406 21698 19458
rect 21982 19406 22034 19458
rect 23998 19406 24050 19458
rect 24222 19406 24274 19458
rect 27358 19406 27410 19458
rect 35982 19406 36034 19458
rect 36430 19406 36482 19458
rect 45614 19406 45666 19458
rect 46174 19406 46226 19458
rect 53454 19406 53506 19458
rect 54126 19406 54178 19458
rect 7758 19294 7810 19346
rect 10334 19294 10386 19346
rect 13918 19294 13970 19346
rect 15374 19294 15426 19346
rect 16158 19294 16210 19346
rect 16606 19294 16658 19346
rect 17166 19294 17218 19346
rect 18062 19294 18114 19346
rect 19630 19294 19682 19346
rect 20750 19294 20802 19346
rect 22990 19294 23042 19346
rect 23550 19294 23602 19346
rect 24894 19294 24946 19346
rect 25342 19294 25394 19346
rect 25790 19294 25842 19346
rect 31166 19294 31218 19346
rect 33406 19294 33458 19346
rect 33854 19294 33906 19346
rect 34302 19294 34354 19346
rect 41470 19294 41522 19346
rect 42590 19294 42642 19346
rect 42926 19294 42978 19346
rect 44158 19294 44210 19346
rect 45950 19294 46002 19346
rect 47854 19294 47906 19346
rect 48974 19294 49026 19346
rect 50654 19294 50706 19346
rect 51662 19294 51714 19346
rect 54014 19294 54066 19346
rect 57710 19294 57762 19346
rect 2382 19182 2434 19234
rect 3614 19182 3666 19234
rect 6862 19182 6914 19234
rect 8990 19182 9042 19234
rect 10222 19182 10274 19234
rect 10894 19182 10946 19234
rect 12462 19182 12514 19234
rect 12910 19182 12962 19234
rect 13806 19182 13858 19234
rect 14142 19182 14194 19234
rect 17614 19182 17666 19234
rect 18286 19182 18338 19234
rect 19518 19182 19570 19234
rect 20302 19182 20354 19234
rect 23326 19182 23378 19234
rect 26350 19182 26402 19234
rect 26574 19182 26626 19234
rect 27022 19182 27074 19234
rect 28030 19182 28082 19234
rect 30718 19182 30770 19234
rect 32958 19182 33010 19234
rect 34750 19182 34802 19234
rect 35310 19182 35362 19234
rect 36094 19182 36146 19234
rect 36654 19182 36706 19234
rect 37662 19182 37714 19234
rect 38334 19182 38386 19234
rect 38894 19182 38946 19234
rect 40014 19182 40066 19234
rect 42030 19182 42082 19234
rect 43822 19182 43874 19234
rect 44046 19182 44098 19234
rect 46398 19182 46450 19234
rect 48750 19182 48802 19234
rect 49086 19182 49138 19234
rect 49870 19182 49922 19234
rect 51438 19182 51490 19234
rect 52222 19182 52274 19234
rect 53566 19182 53618 19234
rect 53790 19182 53842 19234
rect 3278 19070 3330 19122
rect 4062 19070 4114 19122
rect 4958 19070 5010 19122
rect 6638 19070 6690 19122
rect 8654 19070 8706 19122
rect 9662 19070 9714 19122
rect 15262 19070 15314 19122
rect 17838 19070 17890 19122
rect 19294 19070 19346 19122
rect 27470 19070 27522 19122
rect 27694 19070 27746 19122
rect 28478 19070 28530 19122
rect 28814 19070 28866 19122
rect 29598 19070 29650 19122
rect 29934 19070 29986 19122
rect 30606 19070 30658 19122
rect 34862 19070 34914 19122
rect 35086 19070 35138 19122
rect 35534 19070 35586 19122
rect 35758 19070 35810 19122
rect 35870 19070 35922 19122
rect 37886 19070 37938 19122
rect 39118 19070 39170 19122
rect 39678 19070 39730 19122
rect 40462 19070 40514 19122
rect 40798 19070 40850 19122
rect 45838 19070 45890 19122
rect 47630 19070 47682 19122
rect 52110 19070 52162 19122
rect 55806 19070 55858 19122
rect 56926 19070 56978 19122
rect 57262 19070 57314 19122
rect 1934 18958 1986 19010
rect 2830 18958 2882 19010
rect 4622 18958 4674 19010
rect 5854 18958 5906 19010
rect 5966 18958 6018 19010
rect 8094 18958 8146 19010
rect 11342 18958 11394 19010
rect 11790 18958 11842 19010
rect 18622 18958 18674 19010
rect 21758 18958 21810 19010
rect 22878 18958 22930 19010
rect 23102 18958 23154 19010
rect 24222 18958 24274 19010
rect 26462 18958 26514 19010
rect 30382 18958 30434 19010
rect 31838 18958 31890 19010
rect 32510 18958 32562 19010
rect 37774 18958 37826 19010
rect 44718 18958 44770 19010
rect 46958 18958 47010 19010
rect 50206 18958 50258 19010
rect 54686 18958 54738 19010
rect 55470 18958 55522 19010
rect 56254 18958 56306 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 3614 18622 3666 18674
rect 3726 18622 3778 18674
rect 4958 18622 5010 18674
rect 5966 18622 6018 18674
rect 6078 18622 6130 18674
rect 8542 18622 8594 18674
rect 13918 18622 13970 18674
rect 14702 18622 14754 18674
rect 6190 18510 6242 18562
rect 6974 18510 7026 18562
rect 7870 18510 7922 18562
rect 8094 18510 8146 18562
rect 13806 18510 13858 18562
rect 14814 18566 14866 18618
rect 20750 18622 20802 18674
rect 20862 18622 20914 18674
rect 21982 18622 22034 18674
rect 23998 18622 24050 18674
rect 24110 18622 24162 18674
rect 24894 18622 24946 18674
rect 26238 18622 26290 18674
rect 27022 18622 27074 18674
rect 27582 18622 27634 18674
rect 29710 18622 29762 18674
rect 30158 18622 30210 18674
rect 31278 18622 31330 18674
rect 31502 18622 31554 18674
rect 34302 18622 34354 18674
rect 35870 18622 35922 18674
rect 37438 18622 37490 18674
rect 38222 18622 38274 18674
rect 38782 18622 38834 18674
rect 39566 18622 39618 18674
rect 40686 18622 40738 18674
rect 42030 18622 42082 18674
rect 45614 18622 45666 18674
rect 46622 18622 46674 18674
rect 48526 18622 48578 18674
rect 49534 18622 49586 18674
rect 49870 18622 49922 18674
rect 50318 18622 50370 18674
rect 51550 18622 51602 18674
rect 52782 18622 52834 18674
rect 54798 18622 54850 18674
rect 56478 18622 56530 18674
rect 57822 18622 57874 18674
rect 15374 18510 15426 18562
rect 15598 18510 15650 18562
rect 15710 18510 15762 18562
rect 15934 18510 15986 18562
rect 21870 18510 21922 18562
rect 24222 18510 24274 18562
rect 32174 18510 32226 18562
rect 32510 18510 32562 18562
rect 35982 18510 36034 18562
rect 36878 18510 36930 18562
rect 37102 18510 37154 18562
rect 37214 18510 37266 18562
rect 37326 18510 37378 18562
rect 39118 18510 39170 18562
rect 40574 18510 40626 18562
rect 40798 18510 40850 18562
rect 41022 18510 41074 18562
rect 42254 18510 42306 18562
rect 3054 18398 3106 18450
rect 3502 18398 3554 18450
rect 4622 18398 4674 18450
rect 5518 18398 5570 18450
rect 7310 18398 7362 18450
rect 8318 18398 8370 18450
rect 8542 18398 8594 18450
rect 8990 18398 9042 18450
rect 9774 18398 9826 18450
rect 10782 18398 10834 18450
rect 12350 18398 12402 18450
rect 14142 18398 14194 18450
rect 18062 18398 18114 18450
rect 18286 18398 18338 18450
rect 19182 18398 19234 18450
rect 19406 18398 19458 18450
rect 20638 18398 20690 18450
rect 21310 18398 21362 18450
rect 23550 18398 23602 18450
rect 23886 18398 23938 18450
rect 26574 18398 26626 18450
rect 27918 18398 27970 18450
rect 28366 18398 28418 18450
rect 28926 18398 28978 18450
rect 29374 18398 29426 18450
rect 31166 18398 31218 18450
rect 32622 18398 32674 18450
rect 35646 18398 35698 18450
rect 40126 18398 40178 18450
rect 1822 18286 1874 18338
rect 2270 18286 2322 18338
rect 2718 18286 2770 18338
rect 4846 18286 4898 18338
rect 10334 18286 10386 18338
rect 11454 18286 11506 18338
rect 11902 18286 11954 18338
rect 12798 18286 12850 18338
rect 13358 18286 13410 18338
rect 16158 18286 16210 18338
rect 17054 18286 17106 18338
rect 18174 18286 18226 18338
rect 22878 18286 22930 18338
rect 25678 18286 25730 18338
rect 31390 18286 31442 18338
rect 32286 18286 32338 18338
rect 42478 18510 42530 18562
rect 44158 18510 44210 18562
rect 44270 18510 44322 18562
rect 46062 18510 46114 18562
rect 46958 18510 47010 18562
rect 48638 18510 48690 18562
rect 51886 18510 51938 18562
rect 52446 18510 52498 18562
rect 54910 18510 54962 18562
rect 55918 18510 55970 18562
rect 57486 18510 57538 18562
rect 41806 18398 41858 18450
rect 44718 18398 44770 18450
rect 45390 18398 45442 18450
rect 45726 18398 45778 18450
rect 47630 18398 47682 18450
rect 54238 18398 54290 18450
rect 54686 18398 54738 18450
rect 55806 18398 55858 18450
rect 56366 18398 56418 18450
rect 34862 18286 34914 18338
rect 41022 18286 41074 18338
rect 43038 18286 43090 18338
rect 43374 18286 43426 18338
rect 50766 18286 50818 18338
rect 53342 18286 53394 18338
rect 53790 18286 53842 18338
rect 1710 18174 1762 18226
rect 2718 18174 2770 18226
rect 12910 18174 12962 18226
rect 13246 18174 13298 18226
rect 14702 18174 14754 18226
rect 18734 18174 18786 18226
rect 22094 18174 22146 18226
rect 23326 18174 23378 18226
rect 30830 18174 30882 18226
rect 33742 18174 33794 18226
rect 33966 18174 34018 18226
rect 34190 18174 34242 18226
rect 34302 18174 34354 18226
rect 41918 18174 41970 18226
rect 44158 18174 44210 18226
rect 48414 18174 48466 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 3950 17838 4002 17890
rect 4846 17838 4898 17890
rect 7534 17838 7586 17890
rect 9214 17838 9266 17890
rect 10222 17838 10274 17890
rect 11678 17838 11730 17890
rect 17950 17838 18002 17890
rect 18286 17838 18338 17890
rect 25454 17838 25506 17890
rect 25678 17838 25730 17890
rect 27246 17838 27298 17890
rect 31166 17838 31218 17890
rect 34862 17838 34914 17890
rect 35086 17838 35138 17890
rect 35534 17838 35586 17890
rect 36094 17838 36146 17890
rect 36654 17838 36706 17890
rect 40350 17838 40402 17890
rect 42478 17838 42530 17890
rect 46062 17838 46114 17890
rect 46734 17838 46786 17890
rect 50318 17838 50370 17890
rect 51326 17838 51378 17890
rect 55582 17838 55634 17890
rect 56814 17838 56866 17890
rect 3054 17726 3106 17778
rect 6526 17726 6578 17778
rect 8206 17726 8258 17778
rect 9662 17726 9714 17778
rect 12462 17726 12514 17778
rect 12910 17726 12962 17778
rect 15486 17726 15538 17778
rect 16270 17726 16322 17778
rect 17278 17726 17330 17778
rect 20414 17726 20466 17778
rect 24446 17726 24498 17778
rect 32510 17726 32562 17778
rect 33966 17726 34018 17778
rect 34638 17726 34690 17778
rect 36430 17726 36482 17778
rect 36878 17726 36930 17778
rect 37438 17726 37490 17778
rect 39006 17726 39058 17778
rect 39678 17726 39730 17778
rect 40798 17726 40850 17778
rect 41022 17726 41074 17778
rect 42142 17726 42194 17778
rect 42926 17726 42978 17778
rect 46734 17726 46786 17778
rect 47182 17726 47234 17778
rect 48750 17726 48802 17778
rect 49198 17726 49250 17778
rect 49646 17726 49698 17778
rect 50878 17726 50930 17778
rect 52334 17726 52386 17778
rect 52670 17726 52722 17778
rect 7646 17614 7698 17666
rect 8766 17614 8818 17666
rect 9886 17614 9938 17666
rect 10782 17614 10834 17666
rect 11006 17614 11058 17666
rect 11118 17614 11170 17666
rect 11790 17614 11842 17666
rect 13806 17614 13858 17666
rect 14030 17614 14082 17666
rect 14366 17614 14418 17666
rect 15150 17614 15202 17666
rect 16158 17614 16210 17666
rect 17726 17614 17778 17666
rect 19742 17614 19794 17666
rect 21982 17614 22034 17666
rect 23326 17614 23378 17666
rect 23886 17614 23938 17666
rect 25006 17614 25058 17666
rect 25342 17614 25394 17666
rect 27358 17614 27410 17666
rect 28254 17614 28306 17666
rect 29822 17614 29874 17666
rect 32734 17614 32786 17666
rect 33518 17614 33570 17666
rect 35310 17614 35362 17666
rect 35758 17614 35810 17666
rect 38110 17614 38162 17666
rect 40574 17614 40626 17666
rect 41918 17614 41970 17666
rect 44270 17614 44322 17666
rect 44718 17614 44770 17666
rect 53454 17614 53506 17666
rect 56478 17614 56530 17666
rect 2046 17502 2098 17554
rect 7534 17502 7586 17554
rect 8318 17502 8370 17554
rect 8542 17502 8594 17554
rect 16494 17502 16546 17554
rect 19182 17502 19234 17554
rect 19854 17502 19906 17554
rect 21646 17502 21698 17554
rect 23214 17502 23266 17554
rect 23438 17502 23490 17554
rect 25118 17502 25170 17554
rect 26238 17502 26290 17554
rect 26462 17502 26514 17554
rect 26574 17502 26626 17554
rect 31166 17502 31218 17554
rect 31278 17502 31330 17554
rect 32062 17502 32114 17554
rect 32286 17502 32338 17554
rect 38446 17502 38498 17554
rect 41022 17502 41074 17554
rect 53790 17502 53842 17554
rect 55694 17502 55746 17554
rect 56254 17502 56306 17554
rect 57374 17502 57426 17554
rect 4174 17390 4226 17442
rect 4622 17390 4674 17442
rect 4958 17390 5010 17442
rect 5966 17390 6018 17442
rect 11342 17390 11394 17442
rect 18846 17390 18898 17442
rect 20078 17390 20130 17442
rect 20862 17390 20914 17442
rect 21758 17390 21810 17442
rect 22542 17390 22594 17442
rect 25678 17390 25730 17442
rect 27246 17390 27298 17442
rect 27918 17390 27970 17442
rect 28814 17390 28866 17442
rect 29486 17390 29538 17442
rect 29710 17390 29762 17442
rect 30494 17390 30546 17442
rect 33182 17390 33234 17442
rect 35422 17390 35474 17442
rect 38334 17390 38386 17442
rect 41246 17390 41298 17442
rect 43374 17390 43426 17442
rect 45502 17390 45554 17442
rect 45838 17390 45890 17442
rect 46286 17390 46338 17442
rect 47966 17390 48018 17442
rect 48302 17390 48354 17442
rect 50430 17390 50482 17442
rect 51326 17390 51378 17442
rect 51774 17390 51826 17442
rect 54574 17390 54626 17442
rect 54910 17390 54962 17442
rect 55582 17390 55634 17442
rect 57710 17390 57762 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 2158 17054 2210 17106
rect 2494 17054 2546 17106
rect 2942 17054 2994 17106
rect 5630 17054 5682 17106
rect 9102 17054 9154 17106
rect 10110 17054 10162 17106
rect 11006 17054 11058 17106
rect 11902 17054 11954 17106
rect 15038 17054 15090 17106
rect 15374 17054 15426 17106
rect 16606 17054 16658 17106
rect 17054 17054 17106 17106
rect 18174 17054 18226 17106
rect 20190 17054 20242 17106
rect 25566 17054 25618 17106
rect 28142 17054 28194 17106
rect 28590 17054 28642 17106
rect 29934 17054 29986 17106
rect 30718 17054 30770 17106
rect 31726 17054 31778 17106
rect 32174 17054 32226 17106
rect 33966 17054 34018 17106
rect 34750 17054 34802 17106
rect 36318 17054 36370 17106
rect 36654 17054 36706 17106
rect 37102 17054 37154 17106
rect 37550 17054 37602 17106
rect 39118 17054 39170 17106
rect 41918 17054 41970 17106
rect 42366 17054 42418 17106
rect 43374 17054 43426 17106
rect 44270 17054 44322 17106
rect 45726 17054 45778 17106
rect 46846 17054 46898 17106
rect 51998 17054 52050 17106
rect 53566 17054 53618 17106
rect 54910 17054 54962 17106
rect 56702 17054 56754 17106
rect 4398 16942 4450 16994
rect 5742 16942 5794 16994
rect 6078 16942 6130 16994
rect 6974 16942 7026 16994
rect 7310 16942 7362 16994
rect 12238 16942 12290 16994
rect 13582 16942 13634 16994
rect 14478 16942 14530 16994
rect 17726 16942 17778 16994
rect 19966 16942 20018 16994
rect 26574 16942 26626 16994
rect 29150 16942 29202 16994
rect 34414 16942 34466 16994
rect 35534 16942 35586 16994
rect 45390 16942 45442 16994
rect 47854 16942 47906 16994
rect 49646 16942 49698 16994
rect 51550 16942 51602 16994
rect 54462 16942 54514 16994
rect 54686 16942 54738 16994
rect 55918 16942 55970 16994
rect 57486 16942 57538 16994
rect 3390 16830 3442 16882
rect 4622 16830 4674 16882
rect 6414 16830 6466 16882
rect 7198 16830 7250 16882
rect 8654 16830 8706 16882
rect 9774 16830 9826 16882
rect 10670 16830 10722 16882
rect 12798 16830 12850 16882
rect 13246 16830 13298 16882
rect 13918 16830 13970 16882
rect 17950 16830 18002 16882
rect 18846 16830 18898 16882
rect 19406 16830 19458 16882
rect 19742 16830 19794 16882
rect 20750 16830 20802 16882
rect 21310 16830 21362 16882
rect 21646 16830 21698 16882
rect 21870 16830 21922 16882
rect 22654 16830 22706 16882
rect 23102 16830 23154 16882
rect 23774 16830 23826 16882
rect 26462 16830 26514 16882
rect 27694 16830 27746 16882
rect 29486 16830 29538 16882
rect 32510 16830 32562 16882
rect 32734 16830 32786 16882
rect 35646 16830 35698 16882
rect 36094 16830 36146 16882
rect 37998 16830 38050 16882
rect 38894 16830 38946 16882
rect 40014 16830 40066 16882
rect 40350 16830 40402 16882
rect 41470 16830 41522 16882
rect 42814 16830 42866 16882
rect 44606 16830 44658 16882
rect 46174 16830 46226 16882
rect 47182 16830 47234 16882
rect 48190 16830 48242 16882
rect 48414 16830 48466 16882
rect 49982 16830 50034 16882
rect 50542 16830 50594 16882
rect 53006 16830 53058 16882
rect 53230 16830 53282 16882
rect 55022 16830 55074 16882
rect 56254 16830 56306 16882
rect 57710 16830 57762 16882
rect 3950 16718 4002 16770
rect 7534 16718 7586 16770
rect 16046 16718 16098 16770
rect 18286 16718 18338 16770
rect 19854 16718 19906 16770
rect 21422 16718 21474 16770
rect 23662 16718 23714 16770
rect 24894 16718 24946 16770
rect 27358 16718 27410 16770
rect 35310 16718 35362 16770
rect 40574 16718 40626 16770
rect 49758 16718 49810 16770
rect 50318 16718 50370 16770
rect 53566 16718 53618 16770
rect 2158 16606 2210 16658
rect 2942 16606 2994 16658
rect 7758 16606 7810 16658
rect 23438 16606 23490 16658
rect 26574 16606 26626 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 12126 16270 12178 16322
rect 12574 16270 12626 16322
rect 23774 16270 23826 16322
rect 33630 16270 33682 16322
rect 40910 16270 40962 16322
rect 41022 16270 41074 16322
rect 41358 16270 41410 16322
rect 45502 16270 45554 16322
rect 54126 16270 54178 16322
rect 3278 16158 3330 16210
rect 3614 16158 3666 16210
rect 4622 16158 4674 16210
rect 6526 16158 6578 16210
rect 7870 16158 7922 16210
rect 8430 16158 8482 16210
rect 10334 16158 10386 16210
rect 12910 16158 12962 16210
rect 14478 16158 14530 16210
rect 15374 16158 15426 16210
rect 17502 16158 17554 16210
rect 18174 16158 18226 16210
rect 20974 16158 21026 16210
rect 23214 16158 23266 16210
rect 26126 16158 26178 16210
rect 27022 16158 27074 16210
rect 28254 16158 28306 16210
rect 28814 16158 28866 16210
rect 30830 16158 30882 16210
rect 33518 16158 33570 16210
rect 34526 16158 34578 16210
rect 35534 16158 35586 16210
rect 44158 16158 44210 16210
rect 44494 16158 44546 16210
rect 48302 16158 48354 16210
rect 50206 16158 50258 16210
rect 52222 16158 52274 16210
rect 54686 16158 54738 16210
rect 57374 16158 57426 16210
rect 4174 16046 4226 16098
rect 5070 16046 5122 16098
rect 9550 16046 9602 16098
rect 11118 16046 11170 16098
rect 15822 16046 15874 16098
rect 16046 16046 16098 16098
rect 17054 16046 17106 16098
rect 18286 16046 18338 16098
rect 19070 16046 19122 16098
rect 20526 16046 20578 16098
rect 23438 16046 23490 16098
rect 24558 16046 24610 16098
rect 25118 16046 25170 16098
rect 26350 16046 26402 16098
rect 26574 16046 26626 16098
rect 27918 16046 27970 16098
rect 29934 16046 29986 16098
rect 30382 16046 30434 16098
rect 32062 16046 32114 16098
rect 35086 16046 35138 16098
rect 35310 16046 35362 16098
rect 35758 16046 35810 16098
rect 37998 16046 38050 16098
rect 38110 16046 38162 16098
rect 38446 16046 38498 16098
rect 39118 16046 39170 16098
rect 41246 16046 41298 16098
rect 42254 16046 42306 16098
rect 43598 16046 43650 16098
rect 45838 16046 45890 16098
rect 46062 16046 46114 16098
rect 47630 16046 47682 16098
rect 49310 16046 49362 16098
rect 49646 16046 49698 16098
rect 50766 16046 50818 16098
rect 51214 16046 51266 16098
rect 52110 16046 52162 16098
rect 53678 16046 53730 16098
rect 54126 16046 54178 16098
rect 55470 16046 55522 16098
rect 55806 16046 55858 16098
rect 5742 15934 5794 15986
rect 7310 15934 7362 15986
rect 7422 15934 7474 15986
rect 7534 15934 7586 15986
rect 9326 15934 9378 15986
rect 13918 15934 13970 15986
rect 16270 15934 16322 15986
rect 16382 15934 16434 15986
rect 17838 15934 17890 15986
rect 21758 15934 21810 15986
rect 21982 15934 22034 15986
rect 22318 15934 22370 15986
rect 25454 15934 25506 15986
rect 26014 15934 26066 15986
rect 29598 15934 29650 15986
rect 31950 15934 32002 15986
rect 32622 15934 32674 15986
rect 32958 15934 33010 15986
rect 34078 15934 34130 15986
rect 36318 15934 36370 15986
rect 36430 15934 36482 15986
rect 36654 15934 36706 15986
rect 37662 15934 37714 15986
rect 39454 15934 39506 15986
rect 42030 15934 42082 15986
rect 46622 15934 46674 15986
rect 46958 15934 47010 15986
rect 47854 15934 47906 15986
rect 52558 15934 52610 15986
rect 56590 15934 56642 15986
rect 1934 15822 1986 15874
rect 2382 15822 2434 15874
rect 2830 15822 2882 15874
rect 6078 15822 6130 15874
rect 7086 15822 7138 15874
rect 8878 15822 8930 15874
rect 10894 15822 10946 15874
rect 11006 15822 11058 15874
rect 11342 15822 11394 15874
rect 12014 15822 12066 15874
rect 12574 15822 12626 15874
rect 13582 15822 13634 15874
rect 13806 15822 13858 15874
rect 19182 15822 19234 15874
rect 19294 15822 19346 15874
rect 19518 15822 19570 15874
rect 22094 15822 22146 15874
rect 23102 15822 23154 15874
rect 23326 15822 23378 15874
rect 31278 15822 31330 15874
rect 31726 15822 31778 15874
rect 37774 15822 37826 15874
rect 39902 15822 39954 15874
rect 43262 15822 43314 15874
rect 48974 15822 49026 15874
rect 49086 15822 49138 15874
rect 50094 15822 50146 15874
rect 50318 15822 50370 15874
rect 55358 15822 55410 15874
rect 56926 15822 56978 15874
rect 57822 15822 57874 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 2158 15486 2210 15538
rect 2606 15486 2658 15538
rect 3390 15486 3442 15538
rect 3950 15486 4002 15538
rect 5406 15486 5458 15538
rect 6750 15486 6802 15538
rect 8654 15486 8706 15538
rect 9662 15486 9714 15538
rect 11454 15486 11506 15538
rect 13022 15486 13074 15538
rect 16158 15486 16210 15538
rect 16942 15486 16994 15538
rect 18174 15486 18226 15538
rect 22430 15486 22482 15538
rect 22990 15486 23042 15538
rect 23774 15486 23826 15538
rect 24558 15486 24610 15538
rect 24782 15486 24834 15538
rect 25790 15486 25842 15538
rect 28030 15486 28082 15538
rect 29262 15486 29314 15538
rect 29934 15486 29986 15538
rect 31726 15486 31778 15538
rect 32510 15486 32562 15538
rect 33742 15486 33794 15538
rect 34302 15486 34354 15538
rect 34862 15486 34914 15538
rect 35422 15486 35474 15538
rect 36206 15486 36258 15538
rect 36990 15486 37042 15538
rect 38110 15486 38162 15538
rect 38670 15486 38722 15538
rect 39230 15486 39282 15538
rect 39566 15486 39618 15538
rect 40014 15486 40066 15538
rect 40686 15486 40738 15538
rect 41582 15486 41634 15538
rect 44382 15486 44434 15538
rect 45054 15486 45106 15538
rect 45950 15486 46002 15538
rect 46286 15486 46338 15538
rect 46846 15486 46898 15538
rect 51326 15486 51378 15538
rect 51886 15486 51938 15538
rect 53342 15486 53394 15538
rect 53790 15486 53842 15538
rect 54574 15486 54626 15538
rect 56590 15486 56642 15538
rect 57486 15486 57538 15538
rect 9886 15374 9938 15426
rect 10558 15374 10610 15426
rect 10782 15374 10834 15426
rect 16046 15374 16098 15426
rect 16382 15374 16434 15426
rect 17950 15374 18002 15426
rect 21646 15374 21698 15426
rect 26462 15374 26514 15426
rect 26686 15374 26738 15426
rect 33854 15374 33906 15426
rect 35870 15374 35922 15426
rect 37886 15374 37938 15426
rect 42142 15374 42194 15426
rect 42366 15374 42418 15426
rect 45390 15374 45442 15426
rect 46958 15374 47010 15426
rect 48190 15374 48242 15426
rect 48526 15374 48578 15426
rect 53006 15374 53058 15426
rect 54686 15374 54738 15426
rect 54910 15374 54962 15426
rect 55470 15374 55522 15426
rect 3054 15262 3106 15314
rect 4174 15262 4226 15314
rect 4846 15262 4898 15314
rect 5742 15262 5794 15314
rect 6862 15262 6914 15314
rect 7198 15262 7250 15314
rect 8094 15262 8146 15314
rect 9998 15262 10050 15314
rect 12350 15262 12402 15314
rect 12910 15262 12962 15314
rect 13694 15262 13746 15314
rect 14030 15262 14082 15314
rect 15038 15262 15090 15314
rect 15934 15262 15986 15314
rect 18398 15262 18450 15314
rect 18510 15262 18562 15314
rect 19518 15262 19570 15314
rect 19854 15262 19906 15314
rect 20526 15262 20578 15314
rect 21086 15262 21138 15314
rect 23326 15262 23378 15314
rect 24894 15262 24946 15314
rect 27246 15262 27298 15314
rect 27806 15262 27858 15314
rect 28814 15262 28866 15314
rect 30158 15262 30210 15314
rect 30382 15262 30434 15314
rect 30606 15262 30658 15314
rect 32286 15262 32338 15314
rect 32958 15262 33010 15314
rect 33518 15262 33570 15314
rect 36094 15262 36146 15314
rect 36542 15262 36594 15314
rect 37214 15262 37266 15314
rect 37998 15262 38050 15314
rect 42030 15262 42082 15314
rect 42702 15262 42754 15314
rect 43486 15262 43538 15314
rect 43710 15262 43762 15314
rect 50430 15262 50482 15314
rect 52222 15262 52274 15314
rect 54238 15262 54290 15314
rect 55918 15262 55970 15314
rect 57710 15262 57762 15314
rect 7310 15150 7362 15202
rect 8990 15150 9042 15202
rect 11118 15150 11170 15202
rect 12014 15150 12066 15202
rect 20974 15150 21026 15202
rect 26350 15150 26402 15202
rect 30046 15150 30098 15202
rect 31278 15150 31330 15202
rect 32398 15150 32450 15202
rect 43038 15150 43090 15202
rect 43934 15150 43986 15202
rect 47406 15150 47458 15202
rect 49422 15150 49474 15202
rect 50206 15150 50258 15202
rect 50878 15150 50930 15202
rect 52446 15150 52498 15202
rect 56142 15150 56194 15202
rect 11342 15038 11394 15090
rect 18062 15038 18114 15090
rect 25566 15038 25618 15090
rect 26126 15038 26178 15090
rect 30830 15038 30882 15090
rect 55694 15038 55746 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 1822 14702 1874 14754
rect 2270 14702 2322 14754
rect 4174 14702 4226 14754
rect 4958 14702 5010 14754
rect 9550 14702 9602 14754
rect 12126 14702 12178 14754
rect 12910 14702 12962 14754
rect 17054 14702 17106 14754
rect 17390 14702 17442 14754
rect 20414 14702 20466 14754
rect 20974 14702 21026 14754
rect 26238 14702 26290 14754
rect 36094 14702 36146 14754
rect 45950 14702 46002 14754
rect 46286 14702 46338 14754
rect 47854 14702 47906 14754
rect 48078 14702 48130 14754
rect 1934 14590 1986 14642
rect 3614 14590 3666 14642
rect 4062 14590 4114 14642
rect 5854 14590 5906 14642
rect 7646 14590 7698 14642
rect 15598 14590 15650 14642
rect 17054 14590 17106 14642
rect 18062 14590 18114 14642
rect 19070 14590 19122 14642
rect 19854 14590 19906 14642
rect 21870 14590 21922 14642
rect 23102 14590 23154 14642
rect 25230 14590 25282 14642
rect 29598 14590 29650 14642
rect 30270 14590 30322 14642
rect 31278 14590 31330 14642
rect 34638 14590 34690 14642
rect 38446 14590 38498 14642
rect 39790 14590 39842 14642
rect 41246 14590 41298 14642
rect 42926 14590 42978 14642
rect 47182 14590 47234 14642
rect 48190 14590 48242 14642
rect 48750 14590 48802 14642
rect 50318 14590 50370 14642
rect 51102 14590 51154 14642
rect 52222 14590 52274 14642
rect 55358 14590 55410 14642
rect 4510 14478 4562 14530
rect 6862 14478 6914 14530
rect 7758 14478 7810 14530
rect 8654 14478 8706 14530
rect 9102 14478 9154 14530
rect 9326 14478 9378 14530
rect 10334 14478 10386 14530
rect 11454 14478 11506 14530
rect 11790 14478 11842 14530
rect 12910 14478 12962 14530
rect 13694 14478 13746 14530
rect 17390 14478 17442 14530
rect 19630 14478 19682 14530
rect 23774 14478 23826 14530
rect 30046 14478 30098 14530
rect 35534 14478 35586 14530
rect 35982 14478 36034 14530
rect 36318 14478 36370 14530
rect 40462 14478 40514 14530
rect 43150 14478 43202 14530
rect 52334 14478 52386 14530
rect 56030 14478 56082 14530
rect 57934 14478 57986 14530
rect 6414 14366 6466 14418
rect 6638 14366 6690 14418
rect 6974 14366 7026 14418
rect 7534 14366 7586 14418
rect 8094 14366 8146 14418
rect 9774 14366 9826 14418
rect 10446 14366 10498 14418
rect 11006 14366 11058 14418
rect 12014 14366 12066 14418
rect 12574 14366 12626 14418
rect 13918 14366 13970 14418
rect 14478 14366 14530 14418
rect 16046 14366 16098 14418
rect 18734 14366 18786 14418
rect 20078 14366 20130 14418
rect 20302 14366 20354 14418
rect 23326 14366 23378 14418
rect 24670 14366 24722 14418
rect 25566 14366 25618 14418
rect 26574 14366 26626 14418
rect 28814 14366 28866 14418
rect 36542 14366 36594 14418
rect 37550 14366 37602 14418
rect 37886 14366 37938 14418
rect 39006 14366 39058 14418
rect 41694 14366 41746 14418
rect 42478 14366 42530 14418
rect 42926 14366 42978 14418
rect 43710 14366 43762 14418
rect 44046 14366 44098 14418
rect 45502 14366 45554 14418
rect 45614 14366 45666 14418
rect 49422 14366 49474 14418
rect 51326 14366 51378 14418
rect 51662 14366 51714 14418
rect 51774 14366 51826 14418
rect 53902 14366 53954 14418
rect 56702 14366 56754 14418
rect 57038 14366 57090 14418
rect 57598 14366 57650 14418
rect 2382 14254 2434 14306
rect 2830 14254 2882 14306
rect 3278 14254 3330 14306
rect 4958 14254 5010 14306
rect 13806 14254 13858 14306
rect 16382 14254 16434 14306
rect 18958 14254 19010 14306
rect 19182 14254 19234 14306
rect 20862 14254 20914 14306
rect 22430 14254 22482 14306
rect 22990 14254 23042 14306
rect 23214 14254 23266 14306
rect 24334 14254 24386 14306
rect 26350 14254 26402 14306
rect 27022 14254 27074 14306
rect 27582 14254 27634 14306
rect 27918 14254 27970 14306
rect 28478 14254 28530 14306
rect 30494 14254 30546 14306
rect 30606 14254 30658 14306
rect 30718 14254 30770 14306
rect 31726 14254 31778 14306
rect 34302 14254 34354 14306
rect 35086 14254 35138 14306
rect 36654 14254 36706 14306
rect 39342 14254 39394 14306
rect 40798 14254 40850 14306
rect 42702 14254 42754 14306
rect 44494 14254 44546 14306
rect 45838 14254 45890 14306
rect 46286 14254 46338 14306
rect 46734 14254 46786 14306
rect 47630 14254 47682 14306
rect 49534 14254 49586 14306
rect 49646 14254 49698 14306
rect 50654 14254 50706 14306
rect 53566 14254 53618 14306
rect 54350 14254 54402 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 1822 13918 1874 13970
rect 2270 13918 2322 13970
rect 2718 13918 2770 13970
rect 3166 13918 3218 13970
rect 3614 13918 3666 13970
rect 4510 13918 4562 13970
rect 6750 13918 6802 13970
rect 14702 13918 14754 13970
rect 16494 13918 16546 13970
rect 16830 13918 16882 13970
rect 18174 13918 18226 13970
rect 19518 13918 19570 13970
rect 21198 13918 21250 13970
rect 22654 13918 22706 13970
rect 24222 13918 24274 13970
rect 24782 13918 24834 13970
rect 30158 13918 30210 13970
rect 30942 13918 30994 13970
rect 33630 13918 33682 13970
rect 34414 13918 34466 13970
rect 35758 13918 35810 13970
rect 37662 13918 37714 13970
rect 38222 13918 38274 13970
rect 40126 13918 40178 13970
rect 40350 13918 40402 13970
rect 43038 13918 43090 13970
rect 43486 13918 43538 13970
rect 44270 13918 44322 13970
rect 46510 13918 46562 13970
rect 47070 13918 47122 13970
rect 47854 13918 47906 13970
rect 48414 13918 48466 13970
rect 51326 13918 51378 13970
rect 57486 13918 57538 13970
rect 5854 13806 5906 13858
rect 6190 13806 6242 13858
rect 7870 13806 7922 13858
rect 8878 13806 8930 13858
rect 9774 13806 9826 13858
rect 18734 13806 18786 13858
rect 23438 13806 23490 13858
rect 25902 13806 25954 13858
rect 33966 13806 34018 13858
rect 37550 13806 37602 13858
rect 41806 13806 41858 13858
rect 45390 13806 45442 13858
rect 53230 13806 53282 13858
rect 7758 13694 7810 13746
rect 8094 13694 8146 13746
rect 8542 13694 8594 13746
rect 11230 13694 11282 13746
rect 12126 13694 12178 13746
rect 13470 13694 13522 13746
rect 14142 13694 14194 13746
rect 15262 13694 15314 13746
rect 15822 13694 15874 13746
rect 16382 13694 16434 13746
rect 16606 13694 16658 13746
rect 21198 13694 21250 13746
rect 21534 13694 21586 13746
rect 23774 13694 23826 13746
rect 24110 13694 24162 13746
rect 27358 13694 27410 13746
rect 28254 13694 28306 13746
rect 28478 13694 28530 13746
rect 29486 13694 29538 13746
rect 30382 13694 30434 13746
rect 35310 13694 35362 13746
rect 36318 13694 36370 13746
rect 36542 13694 36594 13746
rect 4062 13582 4114 13634
rect 4846 13582 4898 13634
rect 5294 13582 5346 13634
rect 7310 13582 7362 13634
rect 17726 13582 17778 13634
rect 19182 13582 19234 13634
rect 20302 13582 20354 13634
rect 21086 13582 21138 13634
rect 25566 13582 25618 13634
rect 25790 13582 25842 13634
rect 29934 13582 29986 13634
rect 30270 13582 30322 13634
rect 31390 13582 31442 13634
rect 37214 13582 37266 13634
rect 38670 13694 38722 13746
rect 38894 13694 38946 13746
rect 39342 13694 39394 13746
rect 42030 13694 42082 13746
rect 45614 13694 45666 13746
rect 47630 13694 47682 13746
rect 48750 13694 48802 13746
rect 49982 13694 50034 13746
rect 50542 13694 50594 13746
rect 52334 13694 52386 13746
rect 52782 13694 52834 13746
rect 54462 13694 54514 13746
rect 54910 13694 54962 13746
rect 55694 13694 55746 13746
rect 57822 13694 57874 13746
rect 38782 13582 38834 13634
rect 40238 13582 40290 13634
rect 40574 13582 40626 13634
rect 42702 13582 42754 13634
rect 44718 13582 44770 13634
rect 49646 13582 49698 13634
rect 51662 13582 51714 13634
rect 54238 13582 54290 13634
rect 56030 13582 56082 13634
rect 2270 13470 2322 13522
rect 3054 13470 3106 13522
rect 10334 13470 10386 13522
rect 15486 13470 15538 13522
rect 26350 13470 26402 13522
rect 28254 13470 28306 13522
rect 29710 13470 29762 13522
rect 37550 13470 37602 13522
rect 40798 13470 40850 13522
rect 53902 13470 53954 13522
rect 55582 13470 55634 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 16494 13134 16546 13186
rect 16830 13134 16882 13186
rect 22430 13134 22482 13186
rect 24670 13134 24722 13186
rect 24894 13134 24946 13186
rect 27358 13134 27410 13186
rect 28142 13134 28194 13186
rect 28366 13134 28418 13186
rect 40910 13134 40962 13186
rect 48302 13134 48354 13186
rect 55134 13134 55186 13186
rect 1934 13022 1986 13074
rect 4622 13022 4674 13074
rect 7758 13022 7810 13074
rect 10110 13022 10162 13074
rect 15038 13022 15090 13074
rect 18622 13022 18674 13074
rect 20190 13022 20242 13074
rect 21534 13022 21586 13074
rect 22318 13022 22370 13074
rect 22990 13022 23042 13074
rect 27358 13022 27410 13074
rect 29598 13022 29650 13074
rect 30382 13022 30434 13074
rect 30830 13022 30882 13074
rect 32846 13022 32898 13074
rect 35198 13022 35250 13074
rect 36318 13022 36370 13074
rect 36766 13022 36818 13074
rect 38558 13022 38610 13074
rect 41806 13022 41858 13074
rect 44158 13022 44210 13074
rect 44606 13022 44658 13074
rect 45502 13022 45554 13074
rect 48974 13022 49026 13074
rect 49534 13022 49586 13074
rect 53342 13022 53394 13074
rect 55694 13022 55746 13074
rect 56142 13022 56194 13074
rect 57822 13022 57874 13074
rect 2382 12910 2434 12962
rect 6078 12910 6130 12962
rect 7198 12910 7250 12962
rect 9102 12910 9154 12962
rect 11566 12910 11618 12962
rect 12910 12910 12962 12962
rect 16046 12910 16098 12962
rect 16606 12910 16658 12962
rect 16942 12910 16994 12962
rect 17950 12910 18002 12962
rect 18734 12910 18786 12962
rect 19070 12910 19122 12962
rect 19742 12910 19794 12962
rect 20862 12910 20914 12962
rect 22094 12910 22146 12962
rect 25342 12910 25394 12962
rect 26462 12910 26514 12962
rect 31278 12910 31330 12962
rect 33294 12910 33346 12962
rect 33630 12910 33682 12962
rect 37774 12910 37826 12962
rect 39118 12910 39170 12962
rect 39902 12910 39954 12962
rect 40238 12910 40290 12962
rect 41022 12910 41074 12962
rect 42030 12910 42082 12962
rect 46174 12910 46226 12962
rect 46398 12910 46450 12962
rect 47742 12910 47794 12962
rect 47966 12910 48018 12962
rect 49198 12910 49250 12962
rect 51774 12910 51826 12962
rect 3614 12798 3666 12850
rect 8766 12798 8818 12850
rect 10894 12798 10946 12850
rect 12798 12798 12850 12850
rect 14254 12798 14306 12850
rect 14590 12798 14642 12850
rect 17614 12798 17666 12850
rect 20750 12798 20802 12850
rect 23662 12798 23714 12850
rect 23998 12798 24050 12850
rect 25566 12798 25618 12850
rect 28478 12798 28530 12850
rect 33966 12798 34018 12850
rect 34526 12798 34578 12850
rect 34638 12798 34690 12850
rect 39454 12798 39506 12850
rect 40910 12798 40962 12850
rect 42590 12798 42642 12850
rect 43262 12798 43314 12850
rect 49646 12798 49698 12850
rect 51438 12798 51490 12850
rect 52334 12798 52386 12850
rect 52670 12798 52722 12850
rect 54126 12798 54178 12850
rect 54462 12798 54514 12850
rect 55134 12798 55186 12850
rect 55246 12798 55298 12850
rect 57038 12798 57090 12850
rect 57374 12798 57426 12850
rect 2718 12686 2770 12738
rect 3950 12686 4002 12738
rect 5070 12686 5122 12738
rect 13806 12686 13858 12738
rect 15598 12686 15650 12738
rect 18622 12686 18674 12738
rect 18958 12686 19010 12738
rect 24670 12686 24722 12738
rect 26686 12686 26738 12738
rect 27806 12686 27858 12738
rect 29934 12686 29986 12738
rect 33630 12686 33682 12738
rect 34862 12686 34914 12738
rect 35646 12686 35698 12738
rect 37998 12686 38050 12738
rect 40126 12686 40178 12738
rect 43598 12686 43650 12738
rect 47070 12686 47122 12738
rect 49422 12686 49474 12738
rect 50318 12686 50370 12738
rect 50654 12686 50706 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 4398 12350 4450 12402
rect 6078 12350 6130 12402
rect 6190 12350 6242 12402
rect 8654 12350 8706 12402
rect 11678 12350 11730 12402
rect 12238 12350 12290 12402
rect 12574 12350 12626 12402
rect 13134 12350 13186 12402
rect 14030 12350 14082 12402
rect 15150 12350 15202 12402
rect 15710 12350 15762 12402
rect 16046 12350 16098 12402
rect 16606 12350 16658 12402
rect 17950 12350 18002 12402
rect 18734 12350 18786 12402
rect 19854 12350 19906 12402
rect 20638 12350 20690 12402
rect 21422 12350 21474 12402
rect 22878 12350 22930 12402
rect 23662 12350 23714 12402
rect 24222 12350 24274 12402
rect 24558 12350 24610 12402
rect 25566 12350 25618 12402
rect 27582 12350 27634 12402
rect 28590 12350 28642 12402
rect 29822 12350 29874 12402
rect 37550 12350 37602 12402
rect 38334 12350 38386 12402
rect 38670 12350 38722 12402
rect 39230 12350 39282 12402
rect 40014 12350 40066 12402
rect 40574 12350 40626 12402
rect 41470 12350 41522 12402
rect 42254 12350 42306 12402
rect 43374 12350 43426 12402
rect 44830 12350 44882 12402
rect 45726 12350 45778 12402
rect 46174 12350 46226 12402
rect 46734 12350 46786 12402
rect 47294 12350 47346 12402
rect 48750 12350 48802 12402
rect 50878 12350 50930 12402
rect 51662 12350 51714 12402
rect 52558 12350 52610 12402
rect 53118 12350 53170 12402
rect 56030 12350 56082 12402
rect 56590 12350 56642 12402
rect 57374 12350 57426 12402
rect 57822 12350 57874 12402
rect 4062 12238 4114 12290
rect 5070 12238 5122 12290
rect 8094 12238 8146 12290
rect 9662 12238 9714 12290
rect 11118 12238 11170 12290
rect 13470 12238 13522 12290
rect 18958 12238 19010 12290
rect 19518 12238 19570 12290
rect 21870 12238 21922 12290
rect 22094 12238 22146 12290
rect 22206 12238 22258 12290
rect 26462 12238 26514 12290
rect 27470 12238 27522 12290
rect 31166 12238 31218 12290
rect 33966 12238 34018 12290
rect 34414 12238 34466 12290
rect 36318 12238 36370 12290
rect 36878 12238 36930 12290
rect 42702 12238 42754 12290
rect 48638 12238 48690 12290
rect 49870 12238 49922 12290
rect 55134 12238 55186 12290
rect 2830 12126 2882 12178
rect 5182 12126 5234 12178
rect 5854 12126 5906 12178
rect 6974 12126 7026 12178
rect 7646 12126 7698 12178
rect 8990 12126 9042 12178
rect 9886 12126 9938 12178
rect 10446 12126 10498 12178
rect 11006 12126 11058 12178
rect 14366 12126 14418 12178
rect 16830 12126 16882 12178
rect 18510 12126 18562 12178
rect 19854 12126 19906 12178
rect 20078 12126 20130 12178
rect 20862 12126 20914 12178
rect 23214 12126 23266 12178
rect 28926 12126 28978 12178
rect 29598 12126 29650 12178
rect 36094 12126 36146 12178
rect 44606 12126 44658 12178
rect 45390 12126 45442 12178
rect 49646 12126 49698 12178
rect 52222 12126 52274 12178
rect 53342 12126 53394 12178
rect 54238 12126 54290 12178
rect 55694 12126 55746 12178
rect 1934 12014 1986 12066
rect 3614 12014 3666 12066
rect 7982 12014 8034 12066
rect 18846 12014 18898 12066
rect 26014 12014 26066 12066
rect 30270 12014 30322 12066
rect 30718 12014 30770 12066
rect 32846 12014 32898 12066
rect 43710 12014 43762 12066
rect 47742 12014 47794 12066
rect 50318 12014 50370 12066
rect 51214 12014 51266 12066
rect 54350 12014 54402 12066
rect 25454 11902 25506 11954
rect 26014 11902 26066 11954
rect 27694 11902 27746 11954
rect 34638 11902 34690 11954
rect 34974 11902 35026 11954
rect 35758 11902 35810 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 11230 11566 11282 11618
rect 16942 11566 16994 11618
rect 26126 11566 26178 11618
rect 33854 11566 33906 11618
rect 41806 11566 41858 11618
rect 46286 11566 46338 11618
rect 46846 11566 46898 11618
rect 55694 11566 55746 11618
rect 56366 11566 56418 11618
rect 57262 11566 57314 11618
rect 4846 11454 4898 11506
rect 6974 11454 7026 11506
rect 8318 11454 8370 11506
rect 13806 11454 13858 11506
rect 14254 11454 14306 11506
rect 15934 11454 15986 11506
rect 17278 11454 17330 11506
rect 21646 11454 21698 11506
rect 28030 11454 28082 11506
rect 28590 11454 28642 11506
rect 30494 11454 30546 11506
rect 34078 11454 34130 11506
rect 35758 11454 35810 11506
rect 36878 11454 36930 11506
rect 37774 11454 37826 11506
rect 42254 11454 42306 11506
rect 43038 11454 43090 11506
rect 43486 11454 43538 11506
rect 44046 11454 44098 11506
rect 46286 11454 46338 11506
rect 46622 11454 46674 11506
rect 47070 11454 47122 11506
rect 47630 11454 47682 11506
rect 47966 11454 48018 11506
rect 49422 11454 49474 11506
rect 49870 11454 49922 11506
rect 52110 11454 52162 11506
rect 55358 11454 55410 11506
rect 55806 11454 55858 11506
rect 56254 11454 56306 11506
rect 57150 11454 57202 11506
rect 58046 11566 58098 11618
rect 58270 11566 58322 11618
rect 57598 11454 57650 11506
rect 57934 11454 57986 11506
rect 58046 11454 58098 11506
rect 4958 11342 5010 11394
rect 7422 11342 7474 11394
rect 8878 11342 8930 11394
rect 10446 11342 10498 11394
rect 10670 11342 10722 11394
rect 13582 11342 13634 11394
rect 14702 11342 14754 11394
rect 17502 11342 17554 11394
rect 18958 11342 19010 11394
rect 19182 11342 19234 11394
rect 19630 11342 19682 11394
rect 23214 11342 23266 11394
rect 24894 11342 24946 11394
rect 25790 11342 25842 11394
rect 27246 11342 27298 11394
rect 27470 11342 27522 11394
rect 28366 11342 28418 11394
rect 38110 11342 38162 11394
rect 38670 11342 38722 11394
rect 51326 11342 51378 11394
rect 54350 11342 54402 11394
rect 56702 11342 56754 11394
rect 1822 11230 1874 11282
rect 2270 11230 2322 11282
rect 2606 11230 2658 11282
rect 11790 11230 11842 11282
rect 12350 11230 12402 11282
rect 22654 11230 22706 11282
rect 22878 11230 22930 11282
rect 24110 11230 24162 11282
rect 24670 11230 24722 11282
rect 25566 11230 25618 11282
rect 29598 11230 29650 11282
rect 29934 11230 29986 11282
rect 48526 11230 48578 11282
rect 48862 11230 48914 11282
rect 51662 11230 51714 11282
rect 52782 11230 52834 11282
rect 53342 11230 53394 11282
rect 54126 11230 54178 11282
rect 3166 11118 3218 11170
rect 3502 11118 3554 11170
rect 4510 11118 4562 11170
rect 4734 11118 4786 11170
rect 5742 11118 5794 11170
rect 11342 11118 11394 11170
rect 11566 11118 11618 11170
rect 12686 11118 12738 11170
rect 22094 11118 22146 11170
rect 23102 11118 23154 11170
rect 23774 11118 23826 11170
rect 26910 11118 26962 11170
rect 30830 11118 30882 11170
rect 34078 11118 34130 11170
rect 34638 11118 34690 11170
rect 35310 11118 35362 11170
rect 36318 11118 36370 11170
rect 41022 11118 41074 11170
rect 42590 11118 42642 11170
rect 44718 11118 44770 11170
rect 45502 11118 45554 11170
rect 50206 11118 50258 11170
rect 50654 11118 50706 11170
rect 54910 11118 54962 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 2830 10782 2882 10834
rect 3838 10782 3890 10834
rect 4286 10782 4338 10834
rect 4622 10782 4674 10834
rect 6750 10782 6802 10834
rect 12014 10782 12066 10834
rect 12798 10782 12850 10834
rect 14702 10782 14754 10834
rect 15262 10782 15314 10834
rect 17950 10782 18002 10834
rect 18286 10782 18338 10834
rect 24222 10782 24274 10834
rect 25790 10782 25842 10834
rect 26126 10782 26178 10834
rect 27022 10782 27074 10834
rect 29822 10782 29874 10834
rect 37326 10782 37378 10834
rect 38670 10782 38722 10834
rect 39118 10782 39170 10834
rect 40126 10782 40178 10834
rect 40574 10782 40626 10834
rect 41582 10782 41634 10834
rect 42590 10782 42642 10834
rect 43150 10782 43202 10834
rect 47966 10782 48018 10834
rect 49422 10782 49474 10834
rect 49870 10782 49922 10834
rect 50766 10782 50818 10834
rect 51774 10782 51826 10834
rect 52670 10782 52722 10834
rect 53566 10782 53618 10834
rect 53902 10782 53954 10834
rect 54350 10782 54402 10834
rect 54798 10782 54850 10834
rect 55358 10782 55410 10834
rect 55694 10782 55746 10834
rect 57374 10782 57426 10834
rect 57934 10782 57986 10834
rect 2158 10670 2210 10722
rect 2270 10670 2322 10722
rect 3166 10670 3218 10722
rect 5182 10670 5234 10722
rect 6302 10670 6354 10722
rect 7870 10670 7922 10722
rect 8318 10670 8370 10722
rect 8878 10670 8930 10722
rect 14590 10670 14642 10722
rect 14814 10670 14866 10722
rect 15822 10670 15874 10722
rect 18846 10670 18898 10722
rect 20414 10670 20466 10722
rect 22206 10670 22258 10722
rect 27582 10670 27634 10722
rect 28478 10670 28530 10722
rect 30158 10670 30210 10722
rect 34974 10670 35026 10722
rect 36094 10670 36146 10722
rect 5518 10558 5570 10610
rect 6414 10558 6466 10610
rect 7758 10558 7810 10610
rect 10110 10558 10162 10610
rect 10782 10558 10834 10610
rect 11342 10558 11394 10610
rect 12350 10558 12402 10610
rect 13358 10558 13410 10610
rect 16046 10558 16098 10610
rect 16942 10558 16994 10610
rect 19182 10558 19234 10610
rect 19966 10558 20018 10610
rect 20302 10558 20354 10610
rect 22094 10558 22146 10610
rect 23102 10558 23154 10610
rect 23886 10558 23938 10610
rect 23998 10558 24050 10610
rect 24334 10558 24386 10610
rect 27358 10558 27410 10610
rect 28142 10558 28194 10610
rect 34750 10558 34802 10610
rect 35870 10558 35922 10610
rect 45054 10558 45106 10610
rect 45390 10558 45442 10610
rect 51214 10558 51266 10610
rect 10446 10446 10498 10498
rect 13918 10446 13970 10498
rect 16270 10446 16322 10498
rect 20190 10446 20242 10498
rect 21534 10446 21586 10498
rect 22542 10446 22594 10498
rect 24782 10446 24834 10498
rect 29262 10446 29314 10498
rect 37662 10446 37714 10498
rect 38222 10446 38274 10498
rect 39454 10446 39506 10498
rect 41918 10446 41970 10498
rect 43598 10446 43650 10498
rect 44046 10446 44098 10498
rect 44382 10446 44434 10498
rect 50430 10446 50482 10498
rect 52110 10446 52162 10498
rect 53006 10446 53058 10498
rect 56478 10446 56530 10498
rect 43934 10334 43986 10386
rect 44382 10334 44434 10386
rect 44718 10334 44770 10386
rect 48526 10334 48578 10386
rect 50430 10334 50482 10386
rect 51662 10334 51714 10386
rect 53902 10334 53954 10386
rect 54462 10334 54514 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 1934 9998 1986 10050
rect 3166 9998 3218 10050
rect 5966 9998 6018 10050
rect 25678 9998 25730 10050
rect 26574 9998 26626 10050
rect 41694 9998 41746 10050
rect 49086 9998 49138 10050
rect 1934 9886 1986 9938
rect 2382 9886 2434 9938
rect 4062 9886 4114 9938
rect 6414 9886 6466 9938
rect 8094 9886 8146 9938
rect 8878 9886 8930 9938
rect 9998 9886 10050 9938
rect 11342 9886 11394 9938
rect 14142 9886 14194 9938
rect 19854 9886 19906 9938
rect 20414 9886 20466 9938
rect 22206 9886 22258 9938
rect 28254 9886 28306 9938
rect 29486 9886 29538 9938
rect 43038 9886 43090 9938
rect 43374 9886 43426 9938
rect 44382 9886 44434 9938
rect 49422 9886 49474 9938
rect 52446 9886 52498 9938
rect 53342 9886 53394 9938
rect 53790 9886 53842 9938
rect 55134 9886 55186 9938
rect 55582 9886 55634 9938
rect 56254 9886 56306 9938
rect 56702 9886 56754 9938
rect 57262 9886 57314 9938
rect 57598 9886 57650 9938
rect 58046 9886 58098 9938
rect 4958 9774 5010 9826
rect 6190 9774 6242 9826
rect 7086 9774 7138 9826
rect 8990 9774 9042 9826
rect 9662 9774 9714 9826
rect 13806 9774 13858 9826
rect 14366 9774 14418 9826
rect 14926 9774 14978 9826
rect 15262 9774 15314 9826
rect 15934 9774 15986 9826
rect 16158 9774 16210 9826
rect 17502 9774 17554 9826
rect 17838 9774 17890 9826
rect 18958 9774 19010 9826
rect 22318 9774 22370 9826
rect 22542 9774 22594 9826
rect 25902 9774 25954 9826
rect 26126 9774 26178 9826
rect 27022 9774 27074 9826
rect 38222 9774 38274 9826
rect 38670 9774 38722 9826
rect 45502 9774 45554 9826
rect 45950 9774 46002 9826
rect 4622 9662 4674 9714
rect 7310 9662 7362 9714
rect 7422 9662 7474 9714
rect 8542 9662 8594 9714
rect 12910 9662 12962 9714
rect 13918 9662 13970 9714
rect 15374 9662 15426 9714
rect 18622 9662 18674 9714
rect 24110 9662 24162 9714
rect 25454 9662 25506 9714
rect 27358 9662 27410 9714
rect 48302 9662 48354 9714
rect 51886 9662 51938 9714
rect 2830 9550 2882 9602
rect 3166 9550 3218 9602
rect 3726 9550 3778 9602
rect 10782 9550 10834 9602
rect 12014 9550 12066 9602
rect 12574 9550 12626 9602
rect 17950 9550 18002 9602
rect 20862 9550 20914 9602
rect 23214 9550 23266 9602
rect 23774 9550 23826 9602
rect 24558 9550 24610 9602
rect 27806 9550 27858 9602
rect 28702 9550 28754 9602
rect 37550 9550 37602 9602
rect 41022 9550 41074 9602
rect 42142 9550 42194 9602
rect 42478 9550 42530 9602
rect 43934 9550 43986 9602
rect 44718 9550 44770 9602
rect 54238 9550 54290 9602
rect 54686 9550 54738 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 3726 9214 3778 9266
rect 4062 9214 4114 9266
rect 5070 9214 5122 9266
rect 6302 9214 6354 9266
rect 7198 9214 7250 9266
rect 8206 9214 8258 9266
rect 9102 9214 9154 9266
rect 11678 9214 11730 9266
rect 13246 9214 13298 9266
rect 13694 9214 13746 9266
rect 14702 9214 14754 9266
rect 14814 9214 14866 9266
rect 15934 9214 15986 9266
rect 16158 9214 16210 9266
rect 17054 9214 17106 9266
rect 19966 9214 20018 9266
rect 21310 9214 21362 9266
rect 21758 9214 21810 9266
rect 22542 9214 22594 9266
rect 23998 9214 24050 9266
rect 28366 9214 28418 9266
rect 40350 9214 40402 9266
rect 40910 9214 40962 9266
rect 41806 9214 41858 9266
rect 46062 9214 46114 9266
rect 46846 9214 46898 9266
rect 47406 9214 47458 9266
rect 47854 9214 47906 9266
rect 48302 9214 48354 9266
rect 48638 9214 48690 9266
rect 49534 9214 49586 9266
rect 49982 9214 50034 9266
rect 51102 9214 51154 9266
rect 51550 9214 51602 9266
rect 52894 9214 52946 9266
rect 53678 9214 53730 9266
rect 54350 9214 54402 9266
rect 54686 9214 54738 9266
rect 55134 9214 55186 9266
rect 55694 9214 55746 9266
rect 56142 9214 56194 9266
rect 1934 9102 1986 9154
rect 6526 9102 6578 9154
rect 9774 9102 9826 9154
rect 12574 9102 12626 9154
rect 14030 9102 14082 9154
rect 14926 9102 14978 9154
rect 15822 9102 15874 9154
rect 18174 9102 18226 9154
rect 42590 9102 42642 9154
rect 57486 9102 57538 9154
rect 2830 8990 2882 9042
rect 6414 8990 6466 9042
rect 10334 8990 10386 9042
rect 10894 8990 10946 9042
rect 12238 8990 12290 9042
rect 15262 8990 15314 9042
rect 18062 8990 18114 9042
rect 19182 8990 19234 9042
rect 19630 8990 19682 9042
rect 22094 8990 22146 9042
rect 25790 8990 25842 9042
rect 26014 8990 26066 9042
rect 26350 8990 26402 9042
rect 26910 8990 26962 9042
rect 27134 8990 27186 9042
rect 37438 8990 37490 9042
rect 37774 8990 37826 9042
rect 44830 8990 44882 9042
rect 45502 8990 45554 9042
rect 57710 8990 57762 9042
rect 2382 8878 2434 8930
rect 3278 8878 3330 8930
rect 4510 8878 4562 8930
rect 5518 8878 5570 8930
rect 7758 8878 7810 8930
rect 8542 8878 8594 8930
rect 16494 8878 16546 8930
rect 18286 8878 18338 8930
rect 20750 8878 20802 8930
rect 22990 8878 23042 8930
rect 23438 8878 23490 8930
rect 23662 8878 23714 8930
rect 24558 8878 24610 8930
rect 2942 8766 2994 8818
rect 3278 8766 3330 8818
rect 25902 8878 25954 8930
rect 27918 8878 27970 8930
rect 36878 8878 36930 8930
rect 46398 8878 46450 8930
rect 50430 8878 50482 8930
rect 51886 8878 51938 8930
rect 52334 8878 52386 8930
rect 53230 8878 53282 8930
rect 56702 8878 56754 8930
rect 24558 8766 24610 8818
rect 27470 8766 27522 8818
rect 27918 8766 27970 8818
rect 28254 8766 28306 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 57822 8430 57874 8482
rect 58046 8430 58098 8482
rect 1822 8318 1874 8370
rect 2830 8318 2882 8370
rect 3614 8318 3666 8370
rect 4062 8318 4114 8370
rect 4510 8318 4562 8370
rect 5070 8318 5122 8370
rect 6862 8318 6914 8370
rect 11678 8318 11730 8370
rect 12798 8318 12850 8370
rect 15822 8318 15874 8370
rect 16158 8318 16210 8370
rect 16718 8318 16770 8370
rect 17950 8318 18002 8370
rect 18398 8318 18450 8370
rect 20638 8318 20690 8370
rect 21758 8318 21810 8370
rect 24670 8318 24722 8370
rect 42254 8318 42306 8370
rect 42814 8318 42866 8370
rect 43262 8318 43314 8370
rect 43598 8318 43650 8370
rect 44158 8318 44210 8370
rect 44830 8318 44882 8370
rect 50430 8318 50482 8370
rect 50878 8318 50930 8370
rect 51662 8318 51714 8370
rect 52558 8318 52610 8370
rect 53342 8318 53394 8370
rect 53790 8318 53842 8370
rect 55358 8318 55410 8370
rect 56590 8318 56642 8370
rect 57150 8318 57202 8370
rect 6414 8206 6466 8258
rect 6750 8206 6802 8258
rect 7646 8206 7698 8258
rect 8766 8206 8818 8258
rect 10222 8206 10274 8258
rect 10782 8206 10834 8258
rect 17502 8206 17554 8258
rect 18622 8206 18674 8258
rect 19294 8206 19346 8258
rect 26686 8206 26738 8258
rect 38222 8206 38274 8258
rect 38670 8206 38722 8258
rect 45502 8206 45554 8258
rect 45950 8206 46002 8258
rect 49982 8206 50034 8258
rect 51214 8206 51266 8258
rect 56142 8206 56194 8258
rect 7422 8094 7474 8146
rect 11790 8094 11842 8146
rect 14030 8094 14082 8146
rect 14702 8094 14754 8146
rect 23102 8094 23154 8146
rect 23438 8094 23490 8146
rect 25566 8094 25618 8146
rect 26462 8094 26514 8146
rect 41022 8094 41074 8146
rect 41806 8094 41858 8146
rect 52110 8094 52162 8146
rect 2382 7982 2434 8034
rect 3166 7982 3218 8034
rect 13694 7982 13746 8034
rect 15038 7982 15090 8034
rect 19518 7982 19570 8034
rect 20078 7982 20130 8034
rect 22206 7982 22258 8034
rect 22542 7982 22594 8034
rect 23886 7982 23938 8034
rect 25230 7982 25282 8034
rect 27246 7982 27298 8034
rect 27694 7982 27746 8034
rect 37662 7982 37714 8034
rect 48302 7982 48354 8034
rect 49086 7982 49138 8034
rect 49422 7982 49474 8034
rect 54238 7982 54290 8034
rect 57598 7982 57650 8034
rect 58046 7982 58098 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 2494 7646 2546 7698
rect 2942 7646 2994 7698
rect 4286 7646 4338 7698
rect 4622 7646 4674 7698
rect 5182 7646 5234 7698
rect 6526 7646 6578 7698
rect 7310 7646 7362 7698
rect 8990 7646 9042 7698
rect 13582 7646 13634 7698
rect 14254 7646 14306 7698
rect 15150 7646 15202 7698
rect 17838 7646 17890 7698
rect 19854 7646 19906 7698
rect 20862 7646 20914 7698
rect 23886 7646 23938 7698
rect 24894 7646 24946 7698
rect 25678 7646 25730 7698
rect 26910 7646 26962 7698
rect 37998 7646 38050 7698
rect 38334 7646 38386 7698
rect 39118 7646 39170 7698
rect 39566 7646 39618 7698
rect 40462 7646 40514 7698
rect 40910 7646 40962 7698
rect 47294 7646 47346 7698
rect 47854 7646 47906 7698
rect 48526 7646 48578 7698
rect 49534 7646 49586 7698
rect 49870 7646 49922 7698
rect 50318 7646 50370 7698
rect 51662 7646 51714 7698
rect 52334 7646 52386 7698
rect 52782 7646 52834 7698
rect 53230 7646 53282 7698
rect 54014 7646 54066 7698
rect 54350 7646 54402 7698
rect 54798 7646 54850 7698
rect 56590 7646 56642 7698
rect 57374 7646 57426 7698
rect 2046 7534 2098 7586
rect 6638 7534 6690 7586
rect 7534 7534 7586 7586
rect 7758 7534 7810 7586
rect 8654 7534 8706 7586
rect 12126 7534 12178 7586
rect 21870 7534 21922 7586
rect 26126 7534 26178 7586
rect 26462 7534 26514 7586
rect 55246 7534 55298 7586
rect 5518 7422 5570 7474
rect 6078 7422 6130 7474
rect 6414 7422 6466 7474
rect 7086 7422 7138 7474
rect 10334 7422 10386 7474
rect 11454 7422 11506 7474
rect 13694 7422 13746 7474
rect 14590 7422 14642 7474
rect 16382 7422 16434 7474
rect 16942 7422 16994 7474
rect 18174 7422 18226 7474
rect 19070 7422 19122 7474
rect 19294 7422 19346 7474
rect 21646 7422 21698 7474
rect 22766 7422 22818 7474
rect 24558 7422 24610 7474
rect 45726 7422 45778 7474
rect 3390 7310 3442 7362
rect 3838 7310 3890 7362
rect 10558 7310 10610 7362
rect 12686 7310 12738 7362
rect 13022 7310 13074 7362
rect 15710 7310 15762 7362
rect 20302 7310 20354 7362
rect 22542 7310 22594 7362
rect 23438 7310 23490 7362
rect 40014 7310 40066 7362
rect 42142 7310 42194 7362
rect 50878 7310 50930 7362
rect 55694 7310 55746 7362
rect 57822 7310 57874 7362
rect 3390 7198 3442 7250
rect 4510 7198 4562 7250
rect 18734 7198 18786 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 6750 6862 6802 6914
rect 9550 6862 9602 6914
rect 9886 6862 9938 6914
rect 15038 6862 15090 6914
rect 19294 6862 19346 6914
rect 5742 6750 5794 6802
rect 8430 6750 8482 6802
rect 11566 6750 11618 6802
rect 12238 6750 12290 6802
rect 17278 6750 17330 6802
rect 20974 6750 21026 6802
rect 24334 6750 24386 6802
rect 43710 6750 43762 6802
rect 51774 6750 51826 6802
rect 52558 6750 52610 6802
rect 56254 6750 56306 6802
rect 1934 6638 1986 6690
rect 2606 6638 2658 6690
rect 3278 6638 3330 6690
rect 4174 6638 4226 6690
rect 6414 6638 6466 6690
rect 7086 6638 7138 6690
rect 12126 6638 12178 6690
rect 12910 6638 12962 6690
rect 13582 6638 13634 6690
rect 16606 6638 16658 6690
rect 17838 6638 17890 6690
rect 19518 6638 19570 6690
rect 22990 6638 23042 6690
rect 23550 6638 23602 6690
rect 23774 6638 23826 6690
rect 38222 6638 38274 6690
rect 38782 6638 38834 6690
rect 45502 6638 45554 6690
rect 45950 6638 46002 6690
rect 50318 6638 50370 6690
rect 50766 6638 50818 6690
rect 51214 6638 51266 6690
rect 53454 6638 53506 6690
rect 54014 6638 54066 6690
rect 54910 6638 54962 6690
rect 55806 6638 55858 6690
rect 56702 6638 56754 6690
rect 57262 6638 57314 6690
rect 58046 6638 58098 6690
rect 4510 6526 4562 6578
rect 10110 6526 10162 6578
rect 10670 6526 10722 6578
rect 11006 6526 11058 6578
rect 14030 6526 14082 6578
rect 14254 6526 14306 6578
rect 15150 6526 15202 6578
rect 16382 6526 16434 6578
rect 18062 6526 18114 6578
rect 20078 6526 20130 6578
rect 20414 6526 20466 6578
rect 21758 6526 21810 6578
rect 22094 6526 22146 6578
rect 23886 6526 23938 6578
rect 24894 6526 24946 6578
rect 25230 6526 25282 6578
rect 25678 6526 25730 6578
rect 26126 6526 26178 6578
rect 42590 6526 42642 6578
rect 44494 6526 44546 6578
rect 48302 6526 48354 6578
rect 49422 6526 49474 6578
rect 49870 6526 49922 6578
rect 54462 6526 54514 6578
rect 55358 6526 55410 6578
rect 2382 6414 2434 6466
rect 3726 6414 3778 6466
rect 5070 6414 5122 6466
rect 7870 6414 7922 6466
rect 8990 6414 9042 6466
rect 13918 6414 13970 6466
rect 15710 6414 15762 6466
rect 18958 6414 19010 6466
rect 22542 6414 22594 6466
rect 26574 6414 26626 6466
rect 37774 6414 37826 6466
rect 41358 6414 41410 6466
rect 41918 6414 41970 6466
rect 49086 6414 49138 6466
rect 52222 6414 52274 6466
rect 57598 6414 57650 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 3950 6078 4002 6130
rect 4510 6078 4562 6130
rect 4958 6078 5010 6130
rect 5294 6078 5346 6130
rect 5742 6078 5794 6130
rect 6302 6078 6354 6130
rect 6750 6078 6802 6130
rect 7310 6078 7362 6130
rect 8542 6078 8594 6130
rect 10334 6078 10386 6130
rect 11342 6078 11394 6130
rect 12238 6078 12290 6130
rect 12798 6078 12850 6130
rect 13694 6078 13746 6130
rect 14142 6078 14194 6130
rect 15150 6078 15202 6130
rect 15710 6078 15762 6130
rect 16270 6078 16322 6130
rect 18398 6078 18450 6130
rect 19406 6078 19458 6130
rect 20638 6078 20690 6130
rect 21086 6078 21138 6130
rect 22318 6078 22370 6130
rect 22766 6078 22818 6130
rect 23438 6078 23490 6130
rect 25566 6078 25618 6130
rect 36318 6078 36370 6130
rect 40350 6078 40402 6130
rect 44606 6078 44658 6130
rect 45166 6078 45218 6130
rect 46510 6078 46562 6130
rect 46958 6078 47010 6130
rect 48190 6078 48242 6130
rect 48526 6078 48578 6130
rect 53118 6078 53170 6130
rect 53566 6078 53618 6130
rect 54238 6078 54290 6130
rect 54686 6078 54738 6130
rect 55134 6078 55186 6130
rect 55582 6078 55634 6130
rect 56478 6078 56530 6130
rect 57486 6078 57538 6130
rect 57822 6078 57874 6130
rect 10782 5966 10834 6018
rect 13134 5966 13186 6018
rect 24334 5966 24386 6018
rect 45950 5966 46002 6018
rect 52334 5966 52386 6018
rect 2830 5854 2882 5906
rect 12014 5854 12066 5906
rect 19630 5854 19682 5906
rect 23774 5854 23826 5906
rect 24670 5854 24722 5906
rect 37438 5854 37490 5906
rect 37774 5854 37826 5906
rect 41470 5854 41522 5906
rect 42030 5854 42082 5906
rect 45614 5854 45666 5906
rect 49422 5854 49474 5906
rect 49982 5854 50034 5906
rect 1934 5742 1986 5794
rect 3502 5742 3554 5794
rect 7646 5742 7698 5794
rect 8206 5742 8258 5794
rect 9102 5742 9154 5794
rect 9886 5742 9938 5794
rect 14590 5742 14642 5794
rect 16942 5742 16994 5794
rect 17950 5742 18002 5794
rect 18846 5742 18898 5794
rect 21646 5742 21698 5794
rect 36878 5742 36930 5794
rect 47294 5742 47346 5794
rect 55918 5742 55970 5794
rect 13470 5630 13522 5682
rect 14590 5630 14642 5682
rect 40910 5630 40962 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 11118 5294 11170 5346
rect 11342 5294 11394 5346
rect 41134 5294 41186 5346
rect 49086 5294 49138 5346
rect 50766 5294 50818 5346
rect 51214 5294 51266 5346
rect 2158 5182 2210 5234
rect 3390 5182 3442 5234
rect 3726 5182 3778 5234
rect 4510 5182 4562 5234
rect 4958 5182 5010 5234
rect 5854 5182 5906 5234
rect 6302 5182 6354 5234
rect 7310 5182 7362 5234
rect 8206 5182 8258 5234
rect 8766 5182 8818 5234
rect 9214 5182 9266 5234
rect 9662 5182 9714 5234
rect 10110 5182 10162 5234
rect 10558 5182 10610 5234
rect 11118 5182 11170 5234
rect 11566 5182 11618 5234
rect 12910 5182 12962 5234
rect 14030 5182 14082 5234
rect 14814 5182 14866 5234
rect 15374 5182 15426 5234
rect 15822 5182 15874 5234
rect 16270 5182 16322 5234
rect 17838 5182 17890 5234
rect 18286 5182 18338 5234
rect 19070 5182 19122 5234
rect 19518 5182 19570 5234
rect 19966 5182 20018 5234
rect 20862 5182 20914 5234
rect 21534 5182 21586 5234
rect 22094 5182 22146 5234
rect 22990 5182 23042 5234
rect 23662 5182 23714 5234
rect 28814 5182 28866 5234
rect 36430 5182 36482 5234
rect 43934 5182 43986 5234
rect 44718 5182 44770 5234
rect 49870 5182 49922 5234
rect 50318 5182 50370 5234
rect 50766 5182 50818 5234
rect 51102 5182 51154 5234
rect 51662 5182 51714 5234
rect 52110 5182 52162 5234
rect 53342 5182 53394 5234
rect 54238 5182 54290 5234
rect 54574 5182 54626 5234
rect 56702 5182 56754 5234
rect 57150 5182 57202 5234
rect 57598 5182 57650 5234
rect 2606 5070 2658 5122
rect 6862 5070 6914 5122
rect 7870 5070 7922 5122
rect 12238 5070 12290 5122
rect 17278 5070 17330 5122
rect 22430 5070 22482 5122
rect 24110 5070 24162 5122
rect 24894 5070 24946 5122
rect 33854 5070 33906 5122
rect 34638 5070 34690 5122
rect 37438 5070 37490 5122
rect 37998 5070 38050 5122
rect 45614 5070 45666 5122
rect 45950 5070 46002 5122
rect 52446 5070 52498 5122
rect 28366 4958 28418 5010
rect 41918 4958 41970 5010
rect 56254 4958 56306 5010
rect 16830 4846 16882 4898
rect 20302 4846 20354 4898
rect 28030 4846 28082 4898
rect 34190 4846 34242 4898
rect 36878 4846 36930 4898
rect 40574 4846 40626 4898
rect 48526 4846 48578 4898
rect 55022 4846 55074 4898
rect 55918 4846 55970 4898
rect 58046 4846 58098 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 3278 4510 3330 4562
rect 4062 4510 4114 4562
rect 4622 4510 4674 4562
rect 4958 4510 5010 4562
rect 5518 4510 5570 4562
rect 5966 4510 6018 4562
rect 6414 4510 6466 4562
rect 6862 4510 6914 4562
rect 7310 4510 7362 4562
rect 8654 4510 8706 4562
rect 9998 4510 10050 4562
rect 10446 4510 10498 4562
rect 10894 4510 10946 4562
rect 12350 4510 12402 4562
rect 13022 4510 13074 4562
rect 14142 4510 14194 4562
rect 14590 4510 14642 4562
rect 15822 4510 15874 4562
rect 16494 4510 16546 4562
rect 16942 4510 16994 4562
rect 18398 4510 18450 4562
rect 18846 4510 18898 4562
rect 19294 4510 19346 4562
rect 19966 4510 20018 4562
rect 20414 4510 20466 4562
rect 21310 4510 21362 4562
rect 22430 4510 22482 4562
rect 40462 4510 40514 4562
rect 40798 4510 40850 4562
rect 47742 4510 47794 4562
rect 48078 4510 48130 4562
rect 49982 4510 50034 4562
rect 53790 4510 53842 4562
rect 2382 4398 2434 4450
rect 2718 4398 2770 4450
rect 3614 4398 3666 4450
rect 13806 4398 13858 4450
rect 17726 4398 17778 4450
rect 36878 4398 36930 4450
rect 57486 4398 57538 4450
rect 11230 4286 11282 4338
rect 39566 4286 39618 4338
rect 42142 4286 42194 4338
rect 52558 4286 52610 4338
rect 52894 4286 52946 4338
rect 56142 4286 56194 4338
rect 57710 4286 57762 4338
rect 7758 4174 7810 4226
rect 8094 4174 8146 4226
rect 8990 4174 9042 4226
rect 11678 4174 11730 4226
rect 15374 4174 15426 4226
rect 46734 4174 46786 4226
rect 48750 4174 48802 4226
rect 54126 4174 54178 4226
rect 55358 4174 55410 4226
rect 56590 4174 56642 4226
rect 7758 4062 7810 4114
rect 8094 4062 8146 4114
rect 10558 4062 10610 4114
rect 11678 4062 11730 4114
rect 49422 4062 49474 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 18958 3726 19010 3778
rect 19742 3726 19794 3778
rect 5070 3614 5122 3666
rect 7198 3614 7250 3666
rect 7758 3614 7810 3666
rect 8206 3614 8258 3666
rect 8654 3614 8706 3666
rect 9774 3614 9826 3666
rect 10110 3614 10162 3666
rect 10670 3614 10722 3666
rect 11118 3614 11170 3666
rect 13582 3614 13634 3666
rect 14254 3614 14306 3666
rect 14702 3614 14754 3666
rect 15150 3614 15202 3666
rect 15598 3614 15650 3666
rect 16158 3614 16210 3666
rect 16830 3614 16882 3666
rect 19294 3614 19346 3666
rect 19742 3614 19794 3666
rect 20190 3614 20242 3666
rect 25342 3614 25394 3666
rect 31054 3614 31106 3666
rect 35198 3614 35250 3666
rect 38446 3614 38498 3666
rect 41358 3614 41410 3666
rect 41694 3614 41746 3666
rect 43822 3614 43874 3666
rect 45838 3614 45890 3666
rect 46174 3614 46226 3666
rect 46734 3614 46786 3666
rect 47070 3614 47122 3666
rect 47518 3614 47570 3666
rect 48078 3614 48130 3666
rect 48862 3614 48914 3666
rect 49310 3614 49362 3666
rect 51102 3614 51154 3666
rect 51438 3614 51490 3666
rect 51998 3614 52050 3666
rect 53454 3614 53506 3666
rect 55246 3614 55298 3666
rect 56702 3614 56754 3666
rect 57038 3614 57090 3666
rect 57486 3614 57538 3666
rect 57934 3614 57986 3666
rect 2830 3502 2882 3554
rect 12798 3502 12850 3554
rect 18734 3502 18786 3554
rect 24334 3502 24386 3554
rect 30494 3502 30546 3554
rect 34526 3502 34578 3554
rect 39230 3502 39282 3554
rect 45278 3502 45330 3554
rect 49758 3502 49810 3554
rect 50206 3502 50258 3554
rect 52782 3502 52834 3554
rect 55918 3502 55970 3554
rect 1934 3390 1986 3442
rect 4622 3390 4674 3442
rect 5854 3390 5906 3442
rect 11678 3390 11730 3442
rect 17614 3390 17666 3442
rect 23214 3390 23266 3442
rect 29374 3390 29426 3442
rect 40126 3390 40178 3442
rect 42478 3390 42530 3442
rect 44942 3390 44994 3442
rect 37662 3278 37714 3330
rect 38110 3278 38162 3330
rect 50542 3278 50594 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 2688 59200 2800 59800
rect 8064 59200 8176 59800
rect 14112 59200 14224 59800
rect 19488 59200 19600 59800
rect 25536 59200 25648 59800
rect 31584 59200 31696 59800
rect 36960 59200 37072 59800
rect 43008 59200 43120 59800
rect 48384 59200 48496 59800
rect 54432 59200 54544 59800
rect 59808 59200 59920 59800
rect 1932 57204 1988 57214
rect 1932 55410 1988 57148
rect 2716 56196 2772 59200
rect 4172 56308 4228 56318
rect 3052 56196 3108 56206
rect 2716 56194 3108 56196
rect 2716 56142 3054 56194
rect 3106 56142 3108 56194
rect 2716 56140 3108 56142
rect 3052 56130 3108 56140
rect 4172 56082 4228 56252
rect 4732 56308 4788 56318
rect 4732 56214 4788 56252
rect 4172 56030 4174 56082
rect 4226 56030 4228 56082
rect 4172 56018 4228 56030
rect 8092 55970 8148 59200
rect 8092 55918 8094 55970
rect 8146 55918 8148 55970
rect 8092 55906 8148 55918
rect 8876 56082 8932 56094
rect 8876 56030 8878 56082
rect 8930 56030 8932 56082
rect 4476 55692 4740 55702
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4476 55626 4740 55636
rect 1932 55358 1934 55410
rect 1986 55358 1988 55410
rect 1932 55346 1988 55358
rect 3052 55298 3108 55310
rect 3052 55246 3054 55298
rect 3106 55246 3108 55298
rect 3052 55076 3108 55246
rect 3052 55010 3108 55020
rect 3500 55076 3556 55086
rect 3500 54982 3556 55020
rect 4060 55076 4116 55086
rect 2716 53620 2772 53630
rect 2716 53526 2772 53564
rect 3164 53620 3220 53630
rect 3164 53526 3220 53564
rect 2380 53506 2436 53518
rect 2380 53454 2382 53506
rect 2434 53454 2436 53506
rect 2380 52164 2436 53454
rect 2828 52164 2884 52174
rect 2380 52162 2884 52164
rect 2380 52110 2830 52162
rect 2882 52110 2884 52162
rect 2380 52108 2884 52110
rect 2828 52098 2884 52108
rect 1932 52050 1988 52062
rect 1932 51998 1934 52050
rect 1986 51998 1988 52050
rect 1932 51828 1988 51998
rect 1932 51762 1988 51772
rect 3276 49924 3332 49934
rect 3276 48468 3332 49868
rect 2716 48466 3332 48468
rect 2716 48414 3278 48466
rect 3330 48414 3332 48466
rect 2716 48412 3332 48414
rect 2380 48356 2436 48366
rect 2268 48354 2436 48356
rect 2268 48302 2382 48354
rect 2434 48302 2436 48354
rect 2268 48300 2436 48302
rect 1148 48132 1204 48142
rect 1036 41076 1092 41086
rect 1036 4452 1092 41020
rect 1148 6692 1204 48076
rect 1932 45780 1988 45790
rect 1932 45686 1988 45724
rect 1820 42084 1876 42094
rect 1372 42082 1876 42084
rect 1372 42030 1822 42082
rect 1874 42030 1876 42082
rect 1372 42028 1876 42030
rect 1260 27188 1316 27198
rect 1260 16212 1316 27132
rect 1260 16146 1316 16156
rect 1260 15204 1316 15214
rect 1260 10836 1316 15148
rect 1372 12964 1428 42028
rect 1820 42018 1876 42028
rect 1932 40290 1988 40302
rect 1932 40238 1934 40290
rect 1986 40238 1988 40290
rect 1932 39732 1988 40238
rect 1932 39666 1988 39676
rect 2268 34916 2324 48300
rect 2380 48290 2436 48300
rect 2716 48354 2772 48412
rect 3276 48402 3332 48412
rect 2716 48302 2718 48354
rect 2770 48302 2772 48354
rect 2716 48290 2772 48302
rect 3388 46116 3444 46126
rect 2828 45892 2884 45902
rect 2380 45890 2884 45892
rect 2380 45838 2830 45890
rect 2882 45838 2884 45890
rect 2380 45836 2884 45838
rect 2380 45330 2436 45836
rect 2828 45826 2884 45836
rect 2380 45278 2382 45330
rect 2434 45278 2436 45330
rect 2380 45266 2436 45278
rect 3164 45668 3220 45678
rect 2716 45220 2772 45230
rect 2716 45126 2772 45164
rect 2828 43540 2884 43550
rect 2828 43446 2884 43484
rect 3164 43538 3220 45612
rect 3276 45332 3332 45342
rect 3388 45332 3444 46060
rect 3276 45330 3444 45332
rect 3276 45278 3278 45330
rect 3330 45278 3444 45330
rect 3276 45276 3444 45278
rect 3500 45892 3556 45902
rect 3276 45220 3332 45276
rect 3276 45154 3332 45164
rect 3500 43708 3556 45836
rect 3500 43652 3668 43708
rect 3164 43486 3166 43538
rect 3218 43486 3220 43538
rect 3164 43474 3220 43486
rect 3052 42868 3108 42878
rect 2492 42866 3108 42868
rect 2492 42814 3054 42866
rect 3106 42814 3108 42866
rect 2492 42812 3108 42814
rect 2492 41970 2548 42812
rect 3052 42802 3108 42812
rect 2492 41918 2494 41970
rect 2546 41918 2548 41970
rect 2492 41906 2548 41918
rect 2940 42642 2996 42654
rect 2940 42590 2942 42642
rect 2994 42590 2996 42642
rect 2940 41300 2996 42590
rect 3276 42642 3332 42654
rect 3276 42590 3278 42642
rect 3330 42590 3332 42642
rect 2604 41188 2660 41198
rect 2604 41094 2660 41132
rect 2940 41186 2996 41244
rect 2940 41134 2942 41186
rect 2994 41134 2996 41186
rect 2940 41122 2996 41134
rect 3164 42308 3220 42318
rect 3052 41076 3108 41086
rect 3052 40982 3108 41020
rect 3164 40852 3220 42252
rect 3276 41188 3332 42590
rect 3276 41122 3332 41132
rect 3500 42642 3556 42654
rect 3500 42590 3502 42642
rect 3554 42590 3556 42642
rect 3500 41076 3556 42590
rect 3500 41010 3556 41020
rect 3164 40796 3332 40852
rect 3164 40628 3220 40638
rect 2828 40404 2884 40414
rect 2380 40402 2884 40404
rect 2380 40350 2830 40402
rect 2882 40350 2884 40402
rect 2380 40348 2884 40350
rect 2380 39506 2436 40348
rect 2828 40338 2884 40348
rect 3164 39732 3220 40572
rect 2716 39730 3220 39732
rect 2716 39678 3166 39730
rect 3218 39678 3220 39730
rect 2716 39676 3220 39678
rect 2716 39618 2772 39676
rect 3164 39666 3220 39676
rect 2716 39566 2718 39618
rect 2770 39566 2772 39618
rect 2716 39554 2772 39566
rect 2380 39454 2382 39506
rect 2434 39454 2436 39506
rect 2380 39442 2436 39454
rect 2940 35812 2996 35822
rect 2268 34850 2324 34860
rect 2828 34916 2884 34926
rect 2828 34822 2884 34860
rect 1932 34802 1988 34814
rect 1932 34750 1934 34802
rect 1986 34750 1988 34802
rect 1932 34356 1988 34750
rect 1932 34290 1988 34300
rect 1596 32564 1652 32574
rect 1596 21700 1652 32508
rect 2492 32452 2548 32462
rect 2380 31556 2436 31566
rect 2380 31462 2436 31500
rect 2268 31444 2324 31454
rect 1932 30882 1988 30894
rect 2268 30884 2324 31388
rect 1932 30830 1934 30882
rect 1986 30830 1988 30882
rect 1932 30770 1988 30830
rect 1932 30718 1934 30770
rect 1986 30718 1988 30770
rect 1932 30706 1988 30718
rect 2044 30882 2324 30884
rect 2044 30830 2270 30882
rect 2322 30830 2324 30882
rect 2044 30828 2324 30830
rect 1932 29988 1988 29998
rect 2044 29988 2100 30828
rect 2268 30818 2324 30828
rect 2380 30212 2436 30222
rect 2492 30212 2548 32396
rect 2828 31556 2884 31566
rect 2828 31462 2884 31500
rect 2828 30882 2884 30894
rect 2828 30830 2830 30882
rect 2882 30830 2884 30882
rect 2828 30772 2884 30830
rect 2380 30210 2548 30212
rect 2380 30158 2382 30210
rect 2434 30158 2548 30210
rect 2380 30156 2548 30158
rect 2380 30146 2436 30156
rect 1932 29986 2100 29988
rect 1932 29934 1934 29986
rect 1986 29934 2100 29986
rect 1932 29932 2100 29934
rect 1932 29922 1988 29932
rect 1932 28530 1988 28542
rect 1932 28478 1934 28530
rect 1986 28478 1988 28530
rect 1932 28308 1988 28478
rect 1932 28242 1988 28252
rect 1596 21634 1652 21644
rect 1708 27748 1764 27758
rect 1708 20916 1764 27692
rect 1820 27746 1876 27758
rect 1820 27694 1822 27746
rect 1874 27694 1876 27746
rect 1820 27634 1876 27694
rect 1820 27582 1822 27634
rect 1874 27582 1876 27634
rect 1820 26292 1876 27582
rect 1820 26226 1876 26236
rect 1820 25620 1876 25630
rect 1820 24948 1876 25564
rect 1932 25508 1988 25518
rect 1932 25414 1988 25452
rect 1932 24948 1988 24958
rect 1820 24946 1988 24948
rect 1820 24894 1934 24946
rect 1986 24894 1988 24946
rect 1820 24892 1988 24894
rect 1932 24882 1988 24892
rect 2044 24052 2100 29932
rect 2156 29652 2212 29662
rect 2156 29558 2212 29596
rect 2492 29650 2548 30156
rect 2492 29598 2494 29650
rect 2546 29598 2548 29650
rect 2380 28084 2436 28094
rect 2268 27746 2324 27758
rect 2268 27694 2270 27746
rect 2322 27694 2324 27746
rect 2268 26964 2324 27694
rect 2268 26898 2324 26908
rect 2156 26852 2212 26862
rect 2156 26758 2212 26796
rect 2156 26180 2212 26190
rect 2156 26086 2212 26124
rect 2268 25620 2324 25630
rect 2268 25526 2324 25564
rect 2380 24836 2436 28028
rect 2492 26514 2548 29598
rect 2716 30770 2884 30772
rect 2716 30718 2830 30770
rect 2882 30718 2884 30770
rect 2716 30716 2884 30718
rect 2716 28084 2772 30716
rect 2828 30706 2884 30716
rect 2716 28018 2772 28028
rect 2828 29986 2884 29998
rect 2828 29934 2830 29986
rect 2882 29934 2884 29986
rect 2716 27746 2772 27758
rect 2716 27694 2718 27746
rect 2770 27694 2772 27746
rect 2604 27076 2660 27086
rect 2604 26982 2660 27020
rect 2716 26740 2772 27694
rect 2716 26674 2772 26684
rect 2492 26462 2494 26514
rect 2546 26462 2548 26514
rect 2492 26068 2548 26462
rect 2828 26180 2884 29934
rect 2940 29650 2996 35756
rect 3276 31948 3332 40796
rect 3612 38668 3668 43652
rect 3836 42756 3892 42766
rect 3724 42644 3780 42654
rect 3724 42082 3780 42588
rect 3724 42030 3726 42082
rect 3778 42030 3780 42082
rect 3724 41524 3780 42030
rect 3836 41858 3892 42700
rect 3836 41806 3838 41858
rect 3890 41806 3892 41858
rect 3836 41794 3892 41806
rect 3948 41748 4004 41758
rect 3724 41468 3892 41524
rect 3724 41300 3780 41310
rect 3724 41206 3780 41244
rect 3724 41076 3780 41086
rect 3724 40982 3780 41020
rect 3836 39508 3892 41468
rect 3948 41410 4004 41692
rect 3948 41358 3950 41410
rect 4002 41358 4004 41410
rect 3948 41346 4004 41358
rect 4060 39844 4116 55020
rect 4476 54124 4740 54134
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4476 54058 4740 54068
rect 4476 52556 4740 52566
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4476 52490 4740 52500
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 8876 50370 8932 56030
rect 14140 56084 14196 59200
rect 19516 56194 19572 59200
rect 19836 56476 20100 56486
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 19836 56410 20100 56420
rect 19516 56142 19518 56194
rect 19570 56142 19572 56194
rect 19516 56130 19572 56142
rect 25564 56196 25620 59200
rect 25900 56196 25956 56206
rect 25564 56194 25956 56196
rect 25564 56142 25902 56194
rect 25954 56142 25956 56194
rect 25564 56140 25956 56142
rect 25900 56130 25956 56140
rect 29932 56196 29988 56206
rect 14140 56018 14196 56028
rect 14364 56082 14420 56094
rect 14364 56030 14366 56082
rect 14418 56030 14420 56082
rect 10108 55972 10164 55982
rect 8876 50318 8878 50370
rect 8930 50318 8932 50370
rect 8876 50306 8932 50318
rect 9212 50482 9268 50494
rect 9212 50430 9214 50482
rect 9266 50430 9268 50482
rect 9212 49924 9268 50430
rect 9772 49924 9828 49934
rect 9212 49922 9828 49924
rect 9212 49870 9774 49922
rect 9826 49870 9828 49922
rect 9212 49868 9828 49870
rect 9772 49858 9828 49868
rect 9996 49698 10052 49710
rect 9996 49646 9998 49698
rect 10050 49646 10052 49698
rect 9548 49588 9604 49598
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 8764 48244 8820 48254
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 7756 47684 7812 47694
rect 7196 47460 7252 47470
rect 5852 46340 5908 46350
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 5852 45778 5908 46284
rect 6412 46340 6468 46350
rect 6412 46002 6468 46284
rect 6412 45950 6414 46002
rect 6466 45950 6468 46002
rect 6412 45938 6468 45950
rect 5852 45726 5854 45778
rect 5906 45726 5908 45778
rect 5628 45668 5684 45678
rect 5628 45574 5684 45612
rect 5740 45332 5796 45342
rect 5404 45106 5460 45118
rect 5404 45054 5406 45106
rect 5458 45054 5460 45106
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 5068 44100 5124 44110
rect 5068 44006 5124 44044
rect 5404 43540 5460 45054
rect 5404 43474 5460 43484
rect 5740 43762 5796 45276
rect 5852 45106 5908 45726
rect 5852 45054 5854 45106
rect 5906 45054 5908 45106
rect 5852 45042 5908 45054
rect 5964 45778 6020 45790
rect 5964 45726 5966 45778
rect 6018 45726 6020 45778
rect 5964 44546 6020 45726
rect 5964 44494 5966 44546
rect 6018 44494 6020 44546
rect 5964 44482 6020 44494
rect 6076 44212 6132 44222
rect 6636 44212 6692 44222
rect 6076 44210 6692 44212
rect 6076 44158 6078 44210
rect 6130 44158 6638 44210
rect 6690 44158 6692 44210
rect 6076 44156 6692 44158
rect 6076 44146 6132 44156
rect 5740 43710 5742 43762
rect 5794 43710 5796 43762
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4956 42980 5012 42990
rect 4956 42886 5012 42924
rect 5740 42866 5796 43710
rect 5964 44100 6020 44110
rect 5964 43708 6020 44044
rect 6300 43762 6356 44156
rect 6636 44146 6692 44156
rect 6748 44100 6804 44110
rect 6748 44006 6804 44044
rect 6860 44098 6916 44110
rect 6860 44046 6862 44098
rect 6914 44046 6916 44098
rect 6300 43710 6302 43762
rect 6354 43710 6356 43762
rect 5964 43652 6132 43708
rect 6300 43698 6356 43710
rect 6860 43708 6916 44046
rect 5740 42814 5742 42866
rect 5794 42814 5796 42866
rect 5740 42802 5796 42814
rect 4844 42644 4900 42654
rect 4844 42550 4900 42588
rect 5516 42082 5572 42094
rect 5516 42030 5518 42082
rect 5570 42030 5572 42082
rect 5404 41970 5460 41982
rect 5404 41918 5406 41970
rect 5458 41918 5460 41970
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 5404 41300 5460 41918
rect 5516 41748 5572 42030
rect 5740 41970 5796 41982
rect 5740 41918 5742 41970
rect 5794 41918 5796 41970
rect 5740 41860 5796 41918
rect 5964 41972 6020 41982
rect 5964 41878 6020 41916
rect 5740 41794 5796 41804
rect 5516 41682 5572 41692
rect 5404 41244 5572 41300
rect 4956 40852 5012 40862
rect 4956 40626 5012 40796
rect 4956 40574 4958 40626
rect 5010 40574 5012 40626
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4060 39778 4116 39788
rect 4956 39732 5012 40574
rect 4732 39676 5012 39732
rect 5404 40292 5460 40302
rect 4172 39620 4228 39630
rect 4396 39620 4452 39630
rect 4172 39618 4340 39620
rect 4172 39566 4174 39618
rect 4226 39566 4340 39618
rect 4172 39564 4340 39566
rect 4172 39554 4228 39564
rect 3836 39452 4116 39508
rect 4060 39394 4116 39452
rect 4060 39342 4062 39394
rect 4114 39342 4116 39394
rect 4060 39330 4116 39342
rect 3724 39060 3780 39070
rect 3724 38966 3780 39004
rect 3948 38836 4004 38846
rect 4172 38836 4228 38846
rect 4004 38834 4228 38836
rect 4004 38782 4174 38834
rect 4226 38782 4228 38834
rect 4004 38780 4228 38782
rect 3948 38770 4004 38780
rect 4172 38770 4228 38780
rect 4284 38836 4340 39564
rect 4284 38770 4340 38780
rect 4396 38724 4452 39564
rect 4732 39618 4788 39676
rect 4732 39566 4734 39618
rect 4786 39566 4788 39618
rect 4732 39060 4788 39566
rect 4620 38836 4676 38846
rect 4620 38742 4676 38780
rect 4732 38834 4788 39004
rect 4732 38782 4734 38834
rect 4786 38782 4788 38834
rect 4732 38770 4788 38782
rect 4956 39506 5012 39518
rect 4956 39454 4958 39506
rect 5010 39454 5012 39506
rect 3612 38612 3780 38668
rect 4396 38658 4452 38668
rect 3612 38052 3668 38062
rect 3612 37958 3668 37996
rect 3500 34916 3556 34926
rect 3500 34822 3556 34860
rect 3388 32452 3444 32462
rect 3388 32450 3556 32452
rect 3388 32398 3390 32450
rect 3442 32398 3556 32450
rect 3388 32396 3556 32398
rect 3388 32386 3444 32396
rect 3276 31892 3444 31948
rect 3388 31780 3444 31892
rect 3388 31714 3444 31724
rect 3276 31556 3332 31566
rect 2940 29598 2942 29650
rect 2994 29598 2996 29650
rect 2940 28642 2996 29598
rect 2940 28590 2942 28642
rect 2994 28590 2996 28642
rect 2940 28578 2996 28590
rect 3052 31554 3332 31556
rect 3052 31502 3278 31554
rect 3330 31502 3332 31554
rect 3052 31500 3332 31502
rect 2492 25284 2548 26012
rect 2716 26124 2884 26180
rect 2940 26850 2996 26862
rect 2940 26798 2942 26850
rect 2994 26798 2996 26850
rect 2940 26178 2996 26798
rect 2940 26126 2942 26178
rect 2994 26126 2996 26178
rect 2492 25218 2548 25228
rect 2604 25732 2660 25742
rect 2268 24780 2436 24836
rect 2156 24052 2212 24062
rect 2044 23996 2156 24052
rect 2156 23938 2212 23996
rect 2156 23886 2158 23938
rect 2210 23886 2212 23938
rect 2156 23874 2212 23886
rect 2268 23826 2324 24780
rect 2492 24724 2548 24734
rect 2268 23774 2270 23826
rect 2322 23774 2324 23826
rect 2044 23716 2100 23726
rect 1820 23044 1876 23054
rect 1820 22950 1876 22988
rect 1932 22932 1988 22942
rect 1932 22482 1988 22876
rect 1932 22430 1934 22482
rect 1986 22430 1988 22482
rect 1932 22418 1988 22430
rect 2044 21588 2100 23660
rect 2268 23716 2324 23774
rect 2268 23650 2324 23660
rect 2380 24610 2436 24622
rect 2380 24558 2382 24610
rect 2434 24558 2436 24610
rect 2380 23828 2436 24558
rect 2492 23938 2548 24668
rect 2492 23886 2494 23938
rect 2546 23886 2548 23938
rect 2492 23874 2548 23886
rect 2156 23604 2212 23614
rect 2156 21810 2212 23548
rect 2380 23548 2436 23772
rect 2380 23492 2548 23548
rect 2268 23042 2324 23054
rect 2268 22990 2270 23042
rect 2322 22990 2324 23042
rect 2268 22932 2324 22990
rect 2268 22866 2324 22876
rect 2156 21758 2158 21810
rect 2210 21758 2212 21810
rect 2156 21746 2212 21758
rect 2044 21532 2436 21588
rect 2268 21364 2324 21374
rect 1932 20916 1988 20926
rect 1708 20914 1988 20916
rect 1708 20862 1934 20914
rect 1986 20862 1988 20914
rect 1708 20860 1988 20862
rect 1932 20850 1988 20860
rect 2044 20804 2100 20814
rect 1708 20692 1764 20702
rect 1708 18226 1764 20636
rect 1932 20132 1988 20142
rect 1932 19010 1988 20076
rect 1932 18958 1934 19010
rect 1986 18958 1988 19010
rect 1932 18676 1988 18958
rect 1932 18610 1988 18620
rect 1708 18174 1710 18226
rect 1762 18174 1764 18226
rect 1708 18162 1764 18174
rect 1820 18338 1876 18350
rect 1820 18286 1822 18338
rect 1874 18286 1876 18338
rect 1820 18228 1876 18286
rect 1820 17892 1876 18172
rect 1708 17836 1876 17892
rect 1596 17780 1652 17790
rect 1372 12898 1428 12908
rect 1484 13076 1540 13086
rect 1260 10770 1316 10780
rect 1484 8428 1540 13020
rect 1148 6626 1204 6636
rect 1372 8372 1540 8428
rect 1372 5348 1428 8372
rect 1372 5282 1428 5292
rect 1036 4386 1092 4396
rect 1596 2772 1652 17724
rect 1708 15204 1764 17836
rect 2044 17780 2100 20748
rect 2156 20244 2212 20254
rect 2156 20130 2212 20188
rect 2156 20078 2158 20130
rect 2210 20078 2212 20130
rect 2156 20066 2212 20078
rect 2268 18564 2324 21308
rect 2380 20914 2436 21532
rect 2380 20862 2382 20914
rect 2434 20862 2436 20914
rect 2380 20850 2436 20862
rect 2380 19236 2436 19246
rect 2380 19142 2436 19180
rect 1708 15138 1764 15148
rect 1820 17724 2100 17780
rect 2156 18508 2324 18564
rect 1708 14980 1764 14990
rect 1708 8428 1764 14924
rect 1820 14754 1876 17724
rect 2044 17554 2100 17566
rect 2044 17502 2046 17554
rect 2098 17502 2100 17554
rect 2044 16884 2100 17502
rect 2156 17106 2212 18508
rect 2268 18338 2324 18350
rect 2268 18286 2270 18338
rect 2322 18286 2324 18338
rect 2268 17892 2324 18286
rect 2268 17826 2324 17836
rect 2156 17054 2158 17106
rect 2210 17054 2212 17106
rect 2156 17042 2212 17054
rect 2492 17106 2548 23492
rect 2604 20132 2660 25676
rect 2716 25060 2772 26124
rect 2940 25732 2996 26126
rect 2940 25666 2996 25676
rect 2828 25396 2884 25406
rect 2828 25302 2884 25340
rect 2716 23548 2772 25004
rect 2828 25172 2884 25182
rect 2828 24836 2884 25116
rect 2828 24834 2996 24836
rect 2828 24782 2830 24834
rect 2882 24782 2996 24834
rect 2828 24780 2996 24782
rect 2828 24770 2884 24780
rect 2940 24052 2996 24780
rect 3052 24724 3108 31500
rect 3276 31490 3332 31500
rect 3500 31556 3556 32396
rect 3724 31780 3780 38612
rect 3948 38612 4004 38622
rect 3836 32564 3892 32574
rect 3836 32470 3892 32508
rect 3724 31724 3892 31780
rect 3724 31556 3780 31566
rect 3500 31490 3556 31500
rect 3612 31554 3780 31556
rect 3612 31502 3726 31554
rect 3778 31502 3780 31554
rect 3612 31500 3780 31502
rect 3164 30882 3220 30894
rect 3164 30830 3166 30882
rect 3218 30830 3220 30882
rect 3164 30434 3220 30830
rect 3164 30382 3166 30434
rect 3218 30382 3220 30434
rect 3164 30370 3220 30382
rect 3612 30434 3668 31500
rect 3724 31490 3780 31500
rect 3724 31220 3780 31230
rect 3836 31220 3892 31724
rect 3948 31332 4004 38556
rect 4844 38612 4900 38622
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4172 38276 4228 38286
rect 4172 38052 4228 38220
rect 4732 38276 4788 38286
rect 4060 38050 4228 38052
rect 4060 37998 4174 38050
rect 4226 37998 4228 38050
rect 4060 37996 4228 37998
rect 4060 37490 4116 37996
rect 4172 37986 4228 37996
rect 4620 38052 4676 38062
rect 4284 37940 4340 37950
rect 4060 37438 4062 37490
rect 4114 37438 4116 37490
rect 4060 35138 4116 37438
rect 4060 35086 4062 35138
rect 4114 35086 4116 35138
rect 4060 35074 4116 35086
rect 4172 37716 4228 37726
rect 4060 34692 4116 34702
rect 4060 34598 4116 34636
rect 4172 33572 4228 37660
rect 4284 35812 4340 37884
rect 4396 37938 4452 37950
rect 4396 37886 4398 37938
rect 4450 37886 4452 37938
rect 4396 37828 4452 37886
rect 4396 37762 4452 37772
rect 4508 37940 4564 37950
rect 4508 37266 4564 37884
rect 4508 37214 4510 37266
rect 4562 37214 4564 37266
rect 4508 37202 4564 37214
rect 4620 37156 4676 37996
rect 4732 37490 4788 38220
rect 4732 37438 4734 37490
rect 4786 37438 4788 37490
rect 4732 37426 4788 37438
rect 4844 37490 4900 38556
rect 4956 38164 5012 39454
rect 5404 39060 5460 40236
rect 5404 38994 5460 39004
rect 5516 40178 5572 41244
rect 5740 41076 5796 41086
rect 5740 40982 5796 41020
rect 5516 40126 5518 40178
rect 5570 40126 5572 40178
rect 5516 39058 5572 40126
rect 5740 40740 5796 40750
rect 5740 39730 5796 40684
rect 5852 40292 5908 40302
rect 5852 40198 5908 40236
rect 6076 39844 6132 43652
rect 6748 43652 6916 43708
rect 7196 43708 7252 47404
rect 7308 45666 7364 45678
rect 7308 45614 7310 45666
rect 7362 45614 7364 45666
rect 7308 44324 7364 45614
rect 7308 44268 7588 44324
rect 7308 43988 7364 44268
rect 7532 44210 7588 44268
rect 7532 44158 7534 44210
rect 7586 44158 7588 44210
rect 7532 44146 7588 44158
rect 7308 43932 7700 43988
rect 6748 43428 6804 43652
rect 7084 43650 7140 43662
rect 7196 43652 7364 43708
rect 7084 43598 7086 43650
rect 7138 43598 7140 43650
rect 6972 43540 7028 43550
rect 6748 43362 6804 43372
rect 6860 43484 6972 43540
rect 6412 42980 6468 42990
rect 6412 42886 6468 42924
rect 6300 42756 6356 42766
rect 6300 42662 6356 42700
rect 6860 42756 6916 43484
rect 6972 43408 7028 43484
rect 7084 42980 7140 43598
rect 7308 43650 7364 43652
rect 7308 43598 7310 43650
rect 7362 43598 7364 43650
rect 7308 43586 7364 43598
rect 7644 43428 7700 43932
rect 7644 43334 7700 43372
rect 7756 43092 7812 47628
rect 8764 47570 8820 48188
rect 8988 47684 9044 47694
rect 8988 47590 9044 47628
rect 8764 47518 8766 47570
rect 8818 47518 8820 47570
rect 8764 47460 8820 47518
rect 8764 47394 8820 47404
rect 9324 47236 9380 47246
rect 9324 47142 9380 47180
rect 9548 47012 9604 49532
rect 9772 49252 9828 49262
rect 9660 49026 9716 49038
rect 9660 48974 9662 49026
rect 9714 48974 9716 49026
rect 9660 47236 9716 48974
rect 9772 48466 9828 49196
rect 9996 48802 10052 49646
rect 10108 49588 10164 55916
rect 13916 55972 13972 55982
rect 13916 55878 13972 55916
rect 14364 55972 14420 56030
rect 14364 55906 14420 55916
rect 15148 56084 15204 56094
rect 15148 55970 15204 56028
rect 20636 56084 20692 56094
rect 21420 56084 21476 56094
rect 20636 56082 21476 56084
rect 20636 56030 20638 56082
rect 20690 56030 21422 56082
rect 21474 56030 21476 56082
rect 20636 56028 21476 56030
rect 20636 56018 20692 56028
rect 15148 55918 15150 55970
rect 15202 55918 15204 55970
rect 15148 55906 15204 55918
rect 13580 55076 13636 55086
rect 10108 49522 10164 49532
rect 10444 49810 10500 49822
rect 10444 49758 10446 49810
rect 10498 49758 10500 49810
rect 9996 48750 9998 48802
rect 10050 48750 10052 48802
rect 9996 48738 10052 48750
rect 10108 48914 10164 48926
rect 10108 48862 10110 48914
rect 10162 48862 10164 48914
rect 9772 48414 9774 48466
rect 9826 48414 9828 48466
rect 9772 48402 9828 48414
rect 9772 48244 9828 48254
rect 9772 48150 9828 48188
rect 9996 48244 10052 48254
rect 10108 48244 10164 48862
rect 10332 48916 10388 48926
rect 10332 48822 10388 48860
rect 10444 48356 10500 49758
rect 13244 49810 13300 49822
rect 13244 49758 13246 49810
rect 13298 49758 13300 49810
rect 13244 49588 13300 49758
rect 13468 49810 13524 49822
rect 13468 49758 13470 49810
rect 13522 49758 13524 49810
rect 13244 49522 13300 49532
rect 13356 49698 13412 49710
rect 13356 49646 13358 49698
rect 13410 49646 13412 49698
rect 13356 49252 13412 49646
rect 13468 49364 13524 49758
rect 13468 49298 13524 49308
rect 12460 49196 13412 49252
rect 9996 48242 10164 48244
rect 9996 48190 9998 48242
rect 10050 48190 10164 48242
rect 9996 48188 10164 48190
rect 10220 48242 10276 48254
rect 10220 48190 10222 48242
rect 10274 48190 10276 48242
rect 10444 48224 10500 48300
rect 11452 48916 11508 48926
rect 9996 47796 10052 48188
rect 9884 47740 10052 47796
rect 9884 47346 9940 47740
rect 10220 47684 10276 48190
rect 10220 47618 10276 47628
rect 11452 47682 11508 48860
rect 12460 48914 12516 49196
rect 12460 48862 12462 48914
rect 12514 48862 12516 48914
rect 12460 48850 12516 48862
rect 12572 49028 12628 49038
rect 11788 48354 11844 48366
rect 11788 48302 11790 48354
rect 11842 48302 11844 48354
rect 11452 47630 11454 47682
rect 11506 47630 11508 47682
rect 11452 47618 11508 47630
rect 11676 48242 11732 48254
rect 11676 48190 11678 48242
rect 11730 48190 11732 48242
rect 10332 47570 10388 47582
rect 10332 47518 10334 47570
rect 10386 47518 10388 47570
rect 10332 47460 10388 47518
rect 10332 47394 10388 47404
rect 10444 47460 10500 47470
rect 11452 47460 11508 47470
rect 10444 47458 11508 47460
rect 10444 47406 10446 47458
rect 10498 47406 11454 47458
rect 11506 47406 11508 47458
rect 10444 47404 11508 47406
rect 9884 47294 9886 47346
rect 9938 47294 9940 47346
rect 9884 47236 9940 47294
rect 10332 47236 10388 47246
rect 9884 47180 10164 47236
rect 9660 47170 9716 47180
rect 9548 46956 10052 47012
rect 9100 46562 9156 46574
rect 9100 46510 9102 46562
rect 9154 46510 9156 46562
rect 9100 46340 9156 46510
rect 9100 46274 9156 46284
rect 9100 45780 9156 45790
rect 9100 45686 9156 45724
rect 8204 45668 8260 45678
rect 8092 45666 8260 45668
rect 8092 45614 8206 45666
rect 8258 45614 8260 45666
rect 8092 45612 8260 45614
rect 7868 44324 7924 44334
rect 7868 44230 7924 44268
rect 8092 43652 8148 45612
rect 8204 45602 8260 45612
rect 8428 45332 8484 45342
rect 8428 45238 8484 45276
rect 9772 45332 9828 45342
rect 9660 45220 9716 45230
rect 8988 44884 9044 44894
rect 8540 44882 9044 44884
rect 8540 44830 8990 44882
rect 9042 44830 9044 44882
rect 8540 44828 9044 44830
rect 8540 44324 8596 44828
rect 8988 44818 9044 44828
rect 8540 44192 8596 44268
rect 8764 44324 8820 44334
rect 8764 44210 8820 44268
rect 8764 44158 8766 44210
rect 8818 44158 8820 44210
rect 7084 42914 7140 42924
rect 7196 43036 7812 43092
rect 7980 43428 8036 43438
rect 7196 42866 7252 43036
rect 7196 42814 7198 42866
rect 7250 42814 7252 42866
rect 7196 42802 7252 42814
rect 6860 42690 6916 42700
rect 7308 42756 7364 42766
rect 7308 42754 7924 42756
rect 7308 42702 7310 42754
rect 7362 42702 7924 42754
rect 7308 42700 7924 42702
rect 7308 42690 7364 42700
rect 6972 42644 7028 42654
rect 6972 42642 7140 42644
rect 6972 42590 6974 42642
rect 7026 42590 7140 42642
rect 6972 42588 7140 42590
rect 6972 42578 7028 42588
rect 6748 42532 6804 42542
rect 6748 42530 6916 42532
rect 6748 42478 6750 42530
rect 6802 42478 6916 42530
rect 6748 42476 6916 42478
rect 6748 42466 6804 42476
rect 6748 42082 6804 42094
rect 6748 42030 6750 42082
rect 6802 42030 6804 42082
rect 6412 41972 6468 41982
rect 6188 41970 6468 41972
rect 6188 41918 6414 41970
rect 6466 41918 6468 41970
rect 6188 41916 6468 41918
rect 6188 41074 6244 41916
rect 6412 41906 6468 41916
rect 6748 41860 6804 42030
rect 6524 41186 6580 41198
rect 6524 41134 6526 41186
rect 6578 41134 6580 41186
rect 6188 41022 6190 41074
rect 6242 41022 6244 41074
rect 6188 40178 6244 41022
rect 6300 41076 6356 41086
rect 6300 40982 6356 41020
rect 6300 40740 6356 40750
rect 6300 40626 6356 40684
rect 6300 40574 6302 40626
rect 6354 40574 6356 40626
rect 6300 40562 6356 40574
rect 6524 40516 6580 41134
rect 6748 41076 6804 41804
rect 6860 41858 6916 42476
rect 6860 41806 6862 41858
rect 6914 41806 6916 41858
rect 6860 41794 6916 41806
rect 6972 42082 7028 42094
rect 6972 42030 6974 42082
rect 7026 42030 7028 42082
rect 6972 41972 7028 42030
rect 6860 41076 6916 41086
rect 6748 41020 6860 41076
rect 6748 40740 6804 40750
rect 6748 40626 6804 40684
rect 6748 40574 6750 40626
rect 6802 40574 6804 40626
rect 6748 40562 6804 40574
rect 6524 40450 6580 40460
rect 6188 40126 6190 40178
rect 6242 40126 6244 40178
rect 6188 40114 6244 40126
rect 6076 39788 6356 39844
rect 5740 39678 5742 39730
rect 5794 39678 5796 39730
rect 5740 39666 5796 39678
rect 5964 39620 6020 39630
rect 6188 39620 6244 39630
rect 5964 39526 6020 39564
rect 6076 39618 6244 39620
rect 6076 39566 6190 39618
rect 6242 39566 6244 39618
rect 6076 39564 6244 39566
rect 5516 39006 5518 39058
rect 5570 39006 5572 39058
rect 5516 38994 5572 39006
rect 6076 38948 6132 39564
rect 6188 39554 6244 39564
rect 5628 38892 6132 38948
rect 6188 39060 6244 39070
rect 6300 39060 6356 39788
rect 6860 39842 6916 41020
rect 6972 40516 7028 41916
rect 7084 41748 7140 42588
rect 7756 42532 7812 42542
rect 7756 42438 7812 42476
rect 7084 41682 7140 41692
rect 7420 42420 7476 42430
rect 6972 40450 7028 40460
rect 7308 40962 7364 40974
rect 7308 40910 7310 40962
rect 7362 40910 7364 40962
rect 7308 40404 7364 40910
rect 7308 40338 7364 40348
rect 7420 40292 7476 42364
rect 7868 41410 7924 42700
rect 7868 41358 7870 41410
rect 7922 41358 7924 41410
rect 7868 41346 7924 41358
rect 7980 41188 8036 43372
rect 8092 43092 8148 43596
rect 8092 42532 8148 43036
rect 8092 42466 8148 42476
rect 8204 43762 8260 43774
rect 8204 43710 8206 43762
rect 8258 43710 8260 43762
rect 8204 42420 8260 43710
rect 8764 43708 8820 44158
rect 8988 44212 9044 44222
rect 8988 43762 9044 44156
rect 9324 44212 9380 44222
rect 9324 44118 9380 44156
rect 9660 44210 9716 45164
rect 9660 44158 9662 44210
rect 9714 44158 9716 44210
rect 8988 43710 8990 43762
rect 9042 43710 9044 43762
rect 8764 43652 8932 43708
rect 8988 43698 9044 43710
rect 9660 43708 9716 44158
rect 8428 43538 8484 43550
rect 8428 43486 8430 43538
rect 8482 43486 8484 43538
rect 8428 43428 8484 43486
rect 8428 43362 8484 43372
rect 8204 42354 8260 42364
rect 8316 43204 8372 43214
rect 7756 41132 8036 41188
rect 7532 40740 7588 40750
rect 7532 40514 7588 40684
rect 7532 40462 7534 40514
rect 7586 40462 7588 40514
rect 7532 40450 7588 40462
rect 7644 40516 7700 40526
rect 7644 40422 7700 40460
rect 7420 40236 7700 40292
rect 7308 40180 7364 40190
rect 6860 39790 6862 39842
rect 6914 39790 6916 39842
rect 6860 39778 6916 39790
rect 6972 40178 7364 40180
rect 6972 40126 7310 40178
rect 7362 40126 7364 40178
rect 6972 40124 7364 40126
rect 6188 39058 6356 39060
rect 6188 39006 6190 39058
rect 6242 39006 6356 39058
rect 6188 39004 6356 39006
rect 6412 39618 6468 39630
rect 6412 39566 6414 39618
rect 6466 39566 6468 39618
rect 5404 38836 5460 38846
rect 5628 38836 5684 38892
rect 6188 38836 6244 39004
rect 5068 38834 5684 38836
rect 5068 38782 5406 38834
rect 5458 38782 5684 38834
rect 5068 38780 5684 38782
rect 5740 38780 6244 38836
rect 5068 38274 5124 38780
rect 5404 38770 5460 38780
rect 5180 38612 5236 38622
rect 5180 38518 5236 38556
rect 5068 38222 5070 38274
rect 5122 38222 5124 38274
rect 5068 38210 5124 38222
rect 4956 38098 5012 38108
rect 5628 38164 5684 38174
rect 5628 38070 5684 38108
rect 5740 38050 5796 38780
rect 5740 37998 5742 38050
rect 5794 37998 5796 38050
rect 5740 37986 5796 37998
rect 5852 38612 5908 38622
rect 4844 37438 4846 37490
rect 4898 37438 4900 37490
rect 4844 37426 4900 37438
rect 4956 37828 5012 37838
rect 4956 37490 5012 37772
rect 4956 37438 4958 37490
rect 5010 37438 5012 37490
rect 4956 37426 5012 37438
rect 4620 37090 4676 37100
rect 5180 37266 5236 37278
rect 5180 37214 5182 37266
rect 5234 37214 5236 37266
rect 5180 37156 5236 37214
rect 5180 37090 5236 37100
rect 5628 37156 5684 37166
rect 5628 37062 5684 37100
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 5068 36260 5124 36270
rect 5068 36258 5348 36260
rect 5068 36206 5070 36258
rect 5122 36206 5348 36258
rect 5068 36204 5348 36206
rect 5068 36194 5124 36204
rect 4396 35812 4452 35822
rect 4284 35810 4452 35812
rect 4284 35758 4398 35810
rect 4450 35758 4452 35810
rect 4284 35756 4452 35758
rect 4396 35746 4452 35756
rect 4956 35698 5012 35710
rect 4956 35646 4958 35698
rect 5010 35646 5012 35698
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4284 35140 4340 35150
rect 4844 35140 4900 35150
rect 4284 35138 4564 35140
rect 4284 35086 4286 35138
rect 4338 35086 4564 35138
rect 4284 35084 4564 35086
rect 4284 35074 4340 35084
rect 4508 34804 4564 35084
rect 4844 35046 4900 35084
rect 4956 35028 5012 35646
rect 4956 34962 5012 34972
rect 5292 35586 5348 36204
rect 5292 35534 5294 35586
rect 5346 35534 5348 35586
rect 5068 34916 5124 34926
rect 5068 34914 5236 34916
rect 5068 34862 5070 34914
rect 5122 34862 5236 34914
rect 5068 34860 5236 34862
rect 5068 34850 5124 34860
rect 4508 34802 4676 34804
rect 4508 34750 4510 34802
rect 4562 34750 4676 34802
rect 4508 34748 4676 34750
rect 4508 34738 4564 34748
rect 4620 34354 4676 34748
rect 4732 34692 4788 34702
rect 4732 34598 4788 34636
rect 4620 34302 4622 34354
rect 4674 34302 4676 34354
rect 4620 34290 4676 34302
rect 5068 34018 5124 34030
rect 5068 33966 5070 34018
rect 5122 33966 5124 34018
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4396 33572 4452 33582
rect 4172 33570 4452 33572
rect 4172 33518 4398 33570
rect 4450 33518 4452 33570
rect 4172 33516 4452 33518
rect 4396 33506 4452 33516
rect 4508 33460 4564 33470
rect 4508 33346 4564 33404
rect 5068 33460 5124 33966
rect 5068 33394 5124 33404
rect 4508 33294 4510 33346
rect 4562 33294 4564 33346
rect 4508 33282 4564 33294
rect 4732 33346 4788 33358
rect 4732 33294 4734 33346
rect 4786 33294 4788 33346
rect 4732 32786 4788 33294
rect 4732 32734 4734 32786
rect 4786 32734 4788 32786
rect 4732 32722 4788 32734
rect 4284 32452 4340 32462
rect 4284 32358 4340 32396
rect 5180 32452 5236 34860
rect 4844 32338 4900 32350
rect 4844 32286 4846 32338
rect 4898 32286 4900 32338
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4844 32004 4900 32286
rect 5068 32338 5124 32350
rect 5068 32286 5070 32338
rect 5122 32286 5124 32338
rect 5068 32116 5124 32286
rect 5068 32050 5124 32060
rect 4844 31938 4900 31948
rect 4172 31668 4228 31678
rect 4172 31574 4228 31612
rect 4620 31556 4676 31566
rect 4620 31554 5012 31556
rect 4620 31502 4622 31554
rect 4674 31502 5012 31554
rect 4620 31500 5012 31502
rect 4620 31490 4676 31500
rect 3948 31266 4004 31276
rect 3724 31218 3836 31220
rect 3724 31166 3726 31218
rect 3778 31166 3836 31218
rect 3724 31164 3836 31166
rect 3724 31154 3780 31164
rect 3836 31088 3892 31164
rect 4620 31220 4676 31230
rect 4620 31126 4676 31164
rect 4172 30882 4228 30894
rect 4172 30830 4174 30882
rect 4226 30830 4228 30882
rect 4172 30772 4228 30830
rect 4956 30884 5012 31500
rect 5068 31554 5124 31566
rect 5068 31502 5070 31554
rect 5122 31502 5124 31554
rect 5068 31444 5124 31502
rect 5068 31378 5124 31388
rect 5068 31220 5124 31230
rect 5180 31220 5236 32396
rect 5292 32004 5348 35534
rect 5404 34018 5460 34030
rect 5404 33966 5406 34018
rect 5458 33966 5460 34018
rect 5404 33348 5460 33966
rect 5852 33684 5908 38556
rect 6188 38610 6244 38780
rect 6412 38836 6468 39566
rect 6412 38770 6468 38780
rect 6188 38558 6190 38610
rect 6242 38558 6244 38610
rect 6188 38546 6244 38558
rect 6636 38724 6692 38734
rect 6636 38610 6692 38668
rect 6636 38558 6638 38610
rect 6690 38558 6692 38610
rect 6300 38050 6356 38062
rect 6300 37998 6302 38050
rect 6354 37998 6356 38050
rect 5964 37940 6020 37950
rect 5964 37846 6020 37884
rect 6188 37828 6244 37838
rect 6188 37734 6244 37772
rect 6300 37156 6356 37998
rect 6636 37268 6692 38558
rect 6748 38722 6804 38734
rect 6748 38670 6750 38722
rect 6802 38670 6804 38722
rect 6748 38612 6804 38670
rect 6972 38668 7028 40124
rect 7308 40114 7364 40124
rect 7308 39732 7364 39742
rect 7420 39732 7476 40236
rect 7308 39730 7476 39732
rect 7308 39678 7310 39730
rect 7362 39678 7476 39730
rect 7308 39676 7476 39678
rect 7532 40068 7588 40078
rect 7308 39666 7364 39676
rect 6748 38546 6804 38556
rect 6860 38612 7028 38668
rect 7084 38834 7140 38846
rect 7084 38782 7086 38834
rect 7138 38782 7140 38834
rect 6860 37490 6916 38612
rect 7084 37716 7140 38782
rect 7420 38834 7476 38846
rect 7420 38782 7422 38834
rect 7474 38782 7476 38834
rect 7420 38668 7476 38782
rect 6860 37438 6862 37490
rect 6914 37438 6916 37490
rect 6860 37426 6916 37438
rect 6972 37660 7140 37716
rect 7196 38612 7476 38668
rect 6860 37268 6916 37278
rect 6636 37266 6916 37268
rect 6636 37214 6862 37266
rect 6914 37214 6916 37266
rect 6636 37212 6916 37214
rect 6860 37202 6916 37212
rect 6300 37062 6356 37100
rect 6636 36932 6692 36942
rect 6076 36260 6132 36270
rect 6300 36260 6356 36270
rect 6076 36258 6300 36260
rect 6076 36206 6078 36258
rect 6130 36206 6300 36258
rect 6076 36204 6300 36206
rect 6076 36194 6132 36204
rect 6076 35586 6132 35598
rect 6076 35534 6078 35586
rect 6130 35534 6132 35586
rect 6076 35474 6132 35534
rect 6076 35422 6078 35474
rect 6130 35422 6132 35474
rect 6076 34802 6132 35422
rect 6188 35028 6244 35038
rect 6188 34934 6244 34972
rect 6300 34916 6356 36204
rect 6524 36258 6580 36270
rect 6524 36206 6526 36258
rect 6578 36206 6580 36258
rect 6524 35700 6580 36206
rect 6412 35698 6580 35700
rect 6412 35646 6526 35698
rect 6578 35646 6580 35698
rect 6412 35644 6580 35646
rect 6412 35586 6468 35644
rect 6524 35634 6580 35644
rect 6412 35534 6414 35586
rect 6466 35534 6468 35586
rect 6412 35522 6468 35534
rect 6636 35476 6692 36876
rect 6972 36932 7028 37660
rect 6972 36866 7028 36876
rect 7084 37492 7140 37502
rect 7196 37492 7252 38612
rect 7084 37490 7252 37492
rect 7084 37438 7086 37490
rect 7138 37438 7252 37490
rect 7084 37436 7252 37438
rect 7420 38162 7476 38174
rect 7420 38110 7422 38162
rect 7474 38110 7476 38162
rect 6972 36260 7028 36270
rect 6972 36166 7028 36204
rect 7084 35922 7140 37436
rect 7196 37268 7252 37278
rect 7196 36260 7252 37212
rect 7308 37266 7364 37278
rect 7308 37214 7310 37266
rect 7362 37214 7364 37266
rect 7308 36932 7364 37214
rect 7308 36866 7364 36876
rect 7420 37266 7476 38110
rect 7420 37214 7422 37266
rect 7474 37214 7476 37266
rect 7420 36706 7476 37214
rect 7420 36654 7422 36706
rect 7474 36654 7476 36706
rect 7420 36642 7476 36654
rect 7308 36260 7364 36270
rect 7196 36258 7364 36260
rect 7196 36206 7310 36258
rect 7362 36206 7364 36258
rect 7196 36204 7364 36206
rect 7084 35870 7086 35922
rect 7138 35870 7140 35922
rect 7084 35858 7140 35870
rect 7196 36036 7252 36046
rect 7196 35922 7252 35980
rect 7196 35870 7198 35922
rect 7250 35870 7252 35922
rect 7196 35858 7252 35870
rect 6300 34822 6356 34860
rect 6524 35420 6692 35476
rect 6972 35698 7028 35710
rect 6972 35646 6974 35698
rect 7026 35646 7028 35698
rect 6076 34750 6078 34802
rect 6130 34750 6132 34802
rect 5852 33618 5908 33628
rect 5964 34130 6020 34142
rect 5964 34078 5966 34130
rect 6018 34078 6020 34130
rect 5964 33460 6020 34078
rect 6076 34020 6132 34750
rect 6524 34354 6580 35420
rect 6524 34302 6526 34354
rect 6578 34302 6580 34354
rect 6524 34290 6580 34302
rect 6636 34802 6692 34814
rect 6636 34750 6638 34802
rect 6690 34750 6692 34802
rect 6636 34356 6692 34750
rect 6636 34290 6692 34300
rect 6972 34356 7028 35646
rect 7308 35700 7364 36204
rect 7308 35634 7364 35644
rect 6972 34262 7028 34300
rect 7196 35028 7252 35038
rect 6412 34242 6468 34254
rect 6412 34190 6414 34242
rect 6466 34190 6468 34242
rect 6076 33954 6132 33964
rect 6188 34130 6244 34142
rect 6188 34078 6190 34130
rect 6242 34078 6244 34130
rect 5740 33404 6020 33460
rect 5740 33348 5796 33404
rect 5404 33346 5796 33348
rect 5404 33294 5742 33346
rect 5794 33294 5796 33346
rect 5404 33292 5796 33294
rect 5740 33012 5796 33292
rect 5404 32562 5460 32574
rect 5404 32510 5406 32562
rect 5458 32510 5460 32562
rect 5404 32452 5460 32510
rect 5404 32386 5460 32396
rect 5628 32340 5684 32350
rect 5628 32246 5684 32284
rect 5740 32116 5796 32956
rect 5852 33236 5908 33246
rect 6188 33236 6244 34078
rect 6412 34132 6468 34190
rect 7196 34244 7252 34972
rect 6412 34076 6580 34132
rect 5852 33234 6244 33236
rect 5852 33182 5854 33234
rect 5906 33182 6244 33234
rect 5852 33180 6244 33182
rect 6300 33572 6356 33582
rect 5852 32452 5908 33180
rect 5852 32386 5908 32396
rect 6300 32562 6356 33516
rect 6524 32786 6580 34076
rect 7196 34130 7252 34188
rect 7196 34078 7198 34130
rect 7250 34078 7252 34130
rect 7196 34066 7252 34078
rect 7308 33908 7364 33918
rect 7308 33460 7364 33852
rect 6524 32734 6526 32786
rect 6578 32734 6580 32786
rect 6524 32676 6580 32734
rect 6524 32610 6580 32620
rect 6748 33348 6804 33358
rect 6300 32510 6302 32562
rect 6354 32510 6356 32562
rect 6300 32340 6356 32510
rect 6300 32274 6356 32284
rect 5740 32050 5796 32060
rect 6188 32116 6244 32126
rect 5292 31938 5348 31948
rect 6076 32004 6132 32014
rect 6076 31890 6132 31948
rect 6076 31838 6078 31890
rect 6130 31838 6132 31890
rect 6076 31826 6132 31838
rect 5740 31556 5796 31566
rect 5740 31462 5796 31500
rect 6188 31556 6244 32060
rect 6748 32004 6804 33292
rect 7308 33234 7364 33404
rect 7308 33182 7310 33234
rect 7362 33182 7364 33234
rect 7196 33124 7252 33134
rect 7196 33030 7252 33068
rect 7308 32900 7364 33182
rect 6524 31556 6580 31566
rect 6188 31554 6580 31556
rect 6188 31502 6526 31554
rect 6578 31502 6580 31554
rect 6188 31500 6580 31502
rect 5068 31218 5236 31220
rect 5068 31166 5070 31218
rect 5122 31166 5236 31218
rect 5068 31164 5236 31166
rect 5068 31154 5124 31164
rect 5292 30994 5348 31006
rect 5292 30942 5294 30994
rect 5346 30942 5348 30994
rect 4956 30828 5236 30884
rect 4172 30706 4228 30716
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 3612 30382 3614 30434
rect 3666 30382 3668 30434
rect 3612 30370 3668 30382
rect 4284 30434 4340 30446
rect 4284 30382 4286 30434
rect 4338 30382 4340 30434
rect 3724 30100 3780 30110
rect 3724 30006 3780 30044
rect 3276 29986 3332 29998
rect 3276 29934 3278 29986
rect 3330 29934 3332 29986
rect 3164 27972 3220 27982
rect 3164 27878 3220 27916
rect 3276 27634 3332 29934
rect 3836 29988 3892 29998
rect 4172 29988 4228 29998
rect 3276 27582 3278 27634
rect 3330 27582 3332 27634
rect 3276 27570 3332 27582
rect 3388 29652 3444 29662
rect 3164 27188 3220 27198
rect 3388 27188 3444 29596
rect 3500 29314 3556 29326
rect 3500 29262 3502 29314
rect 3554 29262 3556 29314
rect 3500 27412 3556 29262
rect 3724 28868 3780 28878
rect 3724 28754 3780 28812
rect 3724 28702 3726 28754
rect 3778 28702 3780 28754
rect 3724 28690 3780 28702
rect 3724 28084 3780 28094
rect 3612 27746 3668 27758
rect 3612 27694 3614 27746
rect 3666 27694 3668 27746
rect 3612 27636 3668 27694
rect 3612 27570 3668 27580
rect 3500 27356 3668 27412
rect 3500 27188 3556 27198
rect 3388 27132 3500 27188
rect 3164 26964 3220 27132
rect 3500 27122 3556 27132
rect 3500 26964 3556 26974
rect 3164 26962 3556 26964
rect 3164 26910 3502 26962
rect 3554 26910 3556 26962
rect 3164 26908 3556 26910
rect 3500 26898 3556 26908
rect 3612 26964 3668 27356
rect 3724 27188 3780 28028
rect 3836 27524 3892 29932
rect 4060 29986 4228 29988
rect 4060 29934 4174 29986
rect 4226 29934 4228 29986
rect 4060 29932 4228 29934
rect 3948 29314 4004 29326
rect 3948 29262 3950 29314
rect 4002 29262 4004 29314
rect 3948 28308 4004 29262
rect 3948 28242 4004 28252
rect 3948 27860 4004 27870
rect 3948 27766 4004 27804
rect 3836 27468 4004 27524
rect 3836 27188 3892 27198
rect 3724 27132 3836 27188
rect 3500 26628 3556 26638
rect 3500 26514 3556 26572
rect 3500 26462 3502 26514
rect 3554 26462 3556 26514
rect 3500 26450 3556 26462
rect 3612 25732 3668 26908
rect 3836 26850 3892 27132
rect 3836 26798 3838 26850
rect 3890 26798 3892 26850
rect 3836 26786 3892 26798
rect 3836 26516 3892 26526
rect 3836 26422 3892 26460
rect 3500 25730 3668 25732
rect 3500 25678 3614 25730
rect 3666 25678 3668 25730
rect 3500 25676 3668 25678
rect 3276 25284 3332 25294
rect 3276 25190 3332 25228
rect 3052 24668 3332 24724
rect 3052 24498 3108 24510
rect 3052 24446 3054 24498
rect 3106 24446 3108 24498
rect 3052 24276 3108 24446
rect 3052 24210 3108 24220
rect 3164 24164 3220 24202
rect 3164 24098 3220 24108
rect 2940 23996 3108 24052
rect 2940 23882 2996 23894
rect 2940 23830 2942 23882
rect 2994 23830 2996 23882
rect 2940 23716 2996 23830
rect 2940 23650 2996 23660
rect 2716 23492 2884 23548
rect 2828 22596 2884 23492
rect 3052 23154 3108 23996
rect 3052 23102 3054 23154
rect 3106 23102 3108 23154
rect 2828 22540 2996 22596
rect 2828 22372 2884 22382
rect 2828 22278 2884 22316
rect 2828 21700 2884 21710
rect 2828 21606 2884 21644
rect 2604 20066 2660 20076
rect 2716 21588 2772 21598
rect 2604 19906 2660 19918
rect 2604 19854 2606 19906
rect 2658 19854 2660 19906
rect 2604 19796 2660 19854
rect 2604 19730 2660 19740
rect 2716 18564 2772 21532
rect 2828 20916 2884 20926
rect 2940 20916 2996 22540
rect 3052 22260 3108 23102
rect 3052 22194 3108 22204
rect 3164 23940 3220 23950
rect 3164 22036 3220 23884
rect 2828 20914 2996 20916
rect 2828 20862 2830 20914
rect 2882 20862 2996 20914
rect 2828 20860 2996 20862
rect 3052 21980 3220 22036
rect 2828 20850 2884 20860
rect 3052 20692 3108 21980
rect 3052 20626 3108 20636
rect 3164 21700 3220 21710
rect 3052 20356 3108 20366
rect 3052 20242 3108 20300
rect 3052 20190 3054 20242
rect 3106 20190 3108 20242
rect 3052 20178 3108 20190
rect 2940 19348 2996 19358
rect 2828 19010 2884 19022
rect 2828 18958 2830 19010
rect 2882 18958 2884 19010
rect 2828 18788 2884 18958
rect 2828 18722 2884 18732
rect 2492 17054 2494 17106
rect 2546 17054 2548 17106
rect 1932 15874 1988 15886
rect 1932 15822 1934 15874
rect 1986 15822 1988 15874
rect 1932 15428 1988 15822
rect 1932 15362 1988 15372
rect 1820 14702 1822 14754
rect 1874 14702 1876 14754
rect 1820 14690 1876 14702
rect 1932 15092 1988 15102
rect 1932 14642 1988 15036
rect 2044 14980 2100 16828
rect 2492 16772 2548 17054
rect 2492 16706 2548 16716
rect 2604 18508 2772 18564
rect 2156 16658 2212 16670
rect 2156 16606 2158 16658
rect 2210 16606 2212 16658
rect 2156 15538 2212 16606
rect 2604 16548 2660 18508
rect 2716 18338 2772 18350
rect 2716 18286 2718 18338
rect 2770 18286 2772 18338
rect 2716 18226 2772 18286
rect 2716 18174 2718 18226
rect 2770 18174 2772 18226
rect 2716 18162 2772 18174
rect 2156 15486 2158 15538
rect 2210 15486 2212 15538
rect 2156 15474 2212 15486
rect 2268 16492 2660 16548
rect 2268 15316 2324 16492
rect 2604 16324 2660 16492
rect 2604 16258 2660 16268
rect 2940 17106 2996 19292
rect 3052 18450 3108 18462
rect 3052 18398 3054 18450
rect 3106 18398 3108 18450
rect 3052 18340 3108 18398
rect 3052 18274 3108 18284
rect 3052 17780 3108 17790
rect 3052 17686 3108 17724
rect 2940 17054 2942 17106
rect 2994 17054 2996 17106
rect 2940 16658 2996 17054
rect 2940 16606 2942 16658
rect 2994 16606 2996 16658
rect 2380 15876 2436 15886
rect 2380 15874 2548 15876
rect 2380 15822 2382 15874
rect 2434 15822 2548 15874
rect 2380 15820 2548 15822
rect 2380 15810 2436 15820
rect 2044 14914 2100 14924
rect 2156 15260 2324 15316
rect 1932 14590 1934 14642
rect 1986 14590 1988 14642
rect 1932 14578 1988 14590
rect 1820 13972 1876 13982
rect 2156 13972 2212 15260
rect 1820 13970 2212 13972
rect 1820 13918 1822 13970
rect 1874 13918 2212 13970
rect 1820 13916 2212 13918
rect 2268 14754 2324 14766
rect 2268 14702 2270 14754
rect 2322 14702 2324 14754
rect 2268 13970 2324 14702
rect 2268 13918 2270 13970
rect 2322 13918 2324 13970
rect 1820 13906 1876 13916
rect 2268 13522 2324 13918
rect 2380 14306 2436 14318
rect 2380 14254 2382 14306
rect 2434 14254 2436 14306
rect 2380 13636 2436 14254
rect 2492 14196 2548 15820
rect 2828 15874 2884 15886
rect 2828 15822 2830 15874
rect 2882 15822 2884 15874
rect 2716 15764 2772 15774
rect 2604 15652 2660 15662
rect 2604 15538 2660 15596
rect 2604 15486 2606 15538
rect 2658 15486 2660 15538
rect 2604 15474 2660 15486
rect 2716 15316 2772 15708
rect 2716 15250 2772 15260
rect 2828 14532 2884 15822
rect 2940 14644 2996 16606
rect 3052 17220 3108 17230
rect 3052 15540 3108 17164
rect 3164 15876 3220 21644
rect 3276 21698 3332 24668
rect 3388 24500 3444 24510
rect 3388 24406 3444 24444
rect 3500 23940 3556 25676
rect 3612 25666 3668 25676
rect 3724 25282 3780 25294
rect 3724 25230 3726 25282
rect 3778 25230 3780 25282
rect 3276 21646 3278 21698
rect 3330 21646 3332 21698
rect 3276 21588 3332 21646
rect 3276 21522 3332 21532
rect 3388 23884 3556 23940
rect 3612 24948 3668 24958
rect 3612 24276 3668 24892
rect 3276 20580 3332 20590
rect 3276 20486 3332 20524
rect 3388 20468 3444 23884
rect 3500 23716 3556 23726
rect 3500 23622 3556 23660
rect 3500 23156 3556 23166
rect 3500 22036 3556 23100
rect 3612 22596 3668 24220
rect 3724 24164 3780 25230
rect 3948 25060 4004 27468
rect 3724 24098 3780 24108
rect 3836 25004 4004 25060
rect 3836 22596 3892 25004
rect 4060 24948 4116 29932
rect 4172 29922 4228 29932
rect 4172 29316 4228 29326
rect 4172 28754 4228 29260
rect 4172 28702 4174 28754
rect 4226 28702 4228 28754
rect 4172 28690 4228 28702
rect 4172 25284 4228 25294
rect 4172 25190 4228 25228
rect 3948 24892 4116 24948
rect 4284 24948 4340 30382
rect 4620 29986 4676 29998
rect 4620 29934 4622 29986
rect 4674 29934 4676 29986
rect 4620 29652 4676 29934
rect 5068 29988 5124 29998
rect 5068 29894 5124 29932
rect 4620 29586 4676 29596
rect 4844 29540 4900 29550
rect 4396 29316 4452 29326
rect 4396 29222 4452 29260
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4844 28868 4900 29484
rect 4620 28812 4900 28868
rect 5068 29092 5124 29102
rect 4620 28754 4676 28812
rect 4620 28702 4622 28754
rect 4674 28702 4676 28754
rect 4620 28690 4676 28702
rect 5068 28754 5124 29036
rect 5068 28702 5070 28754
rect 5122 28702 5124 28754
rect 5068 28690 5124 28702
rect 4844 28084 4900 28094
rect 4396 27748 4452 27758
rect 4396 27654 4452 27692
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4396 26964 4452 27002
rect 4396 26898 4452 26908
rect 4844 26740 4900 28028
rect 5180 28084 5236 30828
rect 5292 30436 5348 30942
rect 6188 30884 6244 31500
rect 6524 31490 6580 31500
rect 5964 30882 6244 30884
rect 5964 30830 6190 30882
rect 6242 30830 6244 30882
rect 5964 30828 6244 30830
rect 5292 29650 5348 30380
rect 5740 30436 5796 30446
rect 5740 30322 5796 30380
rect 5740 30270 5742 30322
rect 5794 30270 5796 30322
rect 5740 30258 5796 30270
rect 5964 30324 6020 30828
rect 6188 30818 6244 30828
rect 6636 30884 6692 30894
rect 6748 30884 6804 31948
rect 6972 32844 7364 32900
rect 6972 31892 7028 32844
rect 7532 32788 7588 40012
rect 7644 39058 7700 40236
rect 7756 40068 7812 41132
rect 8204 41076 8260 41086
rect 8204 40982 8260 41020
rect 7980 40964 8036 40974
rect 7980 40870 8036 40908
rect 8204 40740 8260 40750
rect 8092 40516 8148 40526
rect 8092 40402 8148 40460
rect 8092 40350 8094 40402
rect 8146 40350 8148 40402
rect 8092 40338 8148 40350
rect 7868 40292 7924 40302
rect 7868 40198 7924 40236
rect 7980 40180 8036 40190
rect 7756 40012 7924 40068
rect 7756 39732 7812 39742
rect 7756 39638 7812 39676
rect 7644 39006 7646 39058
rect 7698 39006 7700 39058
rect 7644 38994 7700 39006
rect 7756 38610 7812 38622
rect 7756 38558 7758 38610
rect 7810 38558 7812 38610
rect 7756 38050 7812 38558
rect 7756 37998 7758 38050
rect 7810 37998 7812 38050
rect 7756 37986 7812 37998
rect 7868 38612 7924 40012
rect 7868 37492 7924 38556
rect 7868 37426 7924 37436
rect 7644 36708 7700 36718
rect 7644 36706 7924 36708
rect 7644 36654 7646 36706
rect 7698 36654 7924 36706
rect 7644 36652 7924 36654
rect 7644 36642 7700 36652
rect 7868 36594 7924 36652
rect 7868 36542 7870 36594
rect 7922 36542 7924 36594
rect 7868 36530 7924 36542
rect 7756 35588 7812 35598
rect 7756 35494 7812 35532
rect 7868 34916 7924 34926
rect 7196 32732 7588 32788
rect 7644 34914 7924 34916
rect 7644 34862 7870 34914
rect 7922 34862 7924 34914
rect 7644 34860 7924 34862
rect 7644 32786 7700 34860
rect 7868 34850 7924 34860
rect 7756 34692 7812 34702
rect 7980 34692 8036 40124
rect 8204 39730 8260 40684
rect 8316 40068 8372 43148
rect 8764 41858 8820 41870
rect 8764 41806 8766 41858
rect 8818 41806 8820 41858
rect 8540 41188 8596 41198
rect 8540 41094 8596 41132
rect 8764 40516 8820 41806
rect 8316 40002 8372 40012
rect 8428 40292 8484 40302
rect 8428 39844 8484 40236
rect 8204 39678 8206 39730
rect 8258 39678 8260 39730
rect 8092 39508 8148 39518
rect 8092 38724 8148 39452
rect 8204 39058 8260 39678
rect 8204 39006 8206 39058
rect 8258 39006 8260 39058
rect 8204 38994 8260 39006
rect 8316 39788 8428 39844
rect 8092 37490 8148 38668
rect 8204 38164 8260 38174
rect 8316 38164 8372 39788
rect 8428 39750 8484 39788
rect 8652 39844 8708 39854
rect 8764 39844 8820 40460
rect 8652 39842 8820 39844
rect 8652 39790 8654 39842
rect 8706 39790 8820 39842
rect 8652 39788 8820 39790
rect 8652 39732 8708 39788
rect 8652 39666 8708 39676
rect 8204 38162 8372 38164
rect 8204 38110 8206 38162
rect 8258 38110 8372 38162
rect 8204 38108 8372 38110
rect 8540 39396 8596 39406
rect 8204 38098 8260 38108
rect 8092 37438 8094 37490
rect 8146 37438 8148 37490
rect 8092 37426 8148 37438
rect 8428 36820 8484 36830
rect 8316 36484 8372 36494
rect 8204 36482 8372 36484
rect 8204 36430 8318 36482
rect 8370 36430 8372 36482
rect 8204 36428 8372 36430
rect 7756 34690 8036 34692
rect 7756 34638 7758 34690
rect 7810 34638 8036 34690
rect 7756 34636 8036 34638
rect 8092 34914 8148 34926
rect 8092 34862 8094 34914
rect 8146 34862 8148 34914
rect 7756 34626 7812 34636
rect 7980 34244 8036 34254
rect 7980 34150 8036 34188
rect 7756 34020 7812 34030
rect 7756 33348 7812 33964
rect 7868 33906 7924 33918
rect 7868 33854 7870 33906
rect 7922 33854 7924 33906
rect 7868 33572 7924 33854
rect 8092 33684 8148 34862
rect 7868 33506 7924 33516
rect 7980 33628 8148 33684
rect 7756 33292 7924 33348
rect 7644 32734 7646 32786
rect 7698 32734 7700 32786
rect 7084 32450 7140 32462
rect 7084 32398 7086 32450
rect 7138 32398 7140 32450
rect 7084 32338 7140 32398
rect 7084 32286 7086 32338
rect 7138 32286 7140 32338
rect 7084 32274 7140 32286
rect 6972 31836 7140 31892
rect 6636 30882 6804 30884
rect 6636 30830 6638 30882
rect 6690 30830 6804 30882
rect 6636 30828 6804 30830
rect 6860 31668 6916 31678
rect 6188 30436 6244 30446
rect 6188 30342 6244 30380
rect 6636 30436 6692 30828
rect 6636 30370 6692 30380
rect 6860 30434 6916 31612
rect 6972 31554 7028 31566
rect 6972 31502 6974 31554
rect 7026 31502 7028 31554
rect 6972 30884 7028 31502
rect 6972 30818 7028 30828
rect 7084 30882 7140 31836
rect 7084 30830 7086 30882
rect 7138 30830 7140 30882
rect 6860 30382 6862 30434
rect 6914 30382 6916 30434
rect 6860 30370 6916 30382
rect 5964 30230 6020 30268
rect 6748 30324 6804 30334
rect 6412 30210 6468 30222
rect 6412 30158 6414 30210
rect 6466 30158 6468 30210
rect 6412 30100 6468 30158
rect 6636 30100 6692 30110
rect 6412 30044 6636 30100
rect 5628 29988 5684 29998
rect 5292 29598 5294 29650
rect 5346 29598 5348 29650
rect 5292 29586 5348 29598
rect 5516 29876 5572 29886
rect 5516 29204 5572 29820
rect 5628 29540 5684 29932
rect 5628 29428 5684 29484
rect 5964 29988 6020 29998
rect 5628 29426 5796 29428
rect 5628 29374 5630 29426
rect 5682 29374 5796 29426
rect 5628 29372 5796 29374
rect 5628 29362 5684 29372
rect 5516 29148 5684 29204
rect 5292 28084 5348 28094
rect 5236 28082 5348 28084
rect 5236 28030 5294 28082
rect 5346 28030 5348 28082
rect 5236 28028 5348 28030
rect 5180 27952 5236 28028
rect 5292 28018 5348 28028
rect 4956 27748 5012 27758
rect 4956 27654 5012 27692
rect 5180 27524 5236 27534
rect 4956 27412 5012 27422
rect 4956 27188 5012 27356
rect 4956 27056 5012 27132
rect 4396 26628 4452 26638
rect 4396 26402 4452 26572
rect 4396 26350 4398 26402
rect 4450 26350 4452 26402
rect 4396 26338 4452 26350
rect 4732 26404 4788 26414
rect 4844 26404 4900 26684
rect 4732 26402 4900 26404
rect 4732 26350 4734 26402
rect 4786 26350 4900 26402
rect 4732 26348 4900 26350
rect 4732 26338 4788 26348
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 3948 23380 4004 24892
rect 4284 24882 4340 24892
rect 4396 25620 4452 25630
rect 4172 24836 4228 24846
rect 4060 24724 4116 24734
rect 4172 24724 4228 24780
rect 4060 24722 4228 24724
rect 4060 24670 4062 24722
rect 4114 24670 4228 24722
rect 4060 24668 4228 24670
rect 4060 24658 4116 24668
rect 3948 23314 4004 23324
rect 4060 23156 4116 23166
rect 4060 23062 4116 23100
rect 3836 22540 4004 22596
rect 3612 22370 3668 22540
rect 3724 22484 3780 22494
rect 3724 22390 3780 22428
rect 3612 22318 3614 22370
rect 3666 22318 3668 22370
rect 3612 22306 3668 22318
rect 3948 22372 4004 22540
rect 3836 22260 3892 22270
rect 3836 22166 3892 22204
rect 3500 21980 3892 22036
rect 3836 21810 3892 21980
rect 3836 21758 3838 21810
rect 3890 21758 3892 21810
rect 3836 21746 3892 21758
rect 3500 21476 3556 21486
rect 3500 21382 3556 21420
rect 3388 20402 3444 20412
rect 3724 20578 3780 20590
rect 3724 20526 3726 20578
rect 3778 20526 3780 20578
rect 3388 20020 3444 20030
rect 3444 19964 3556 20020
rect 3388 19926 3444 19964
rect 3276 19124 3332 19134
rect 3276 19030 3332 19068
rect 3500 18676 3556 19964
rect 3724 19460 3780 20526
rect 3724 19394 3780 19404
rect 3612 19236 3668 19246
rect 3612 18900 3668 19180
rect 3612 18834 3668 18844
rect 3948 19236 4004 22316
rect 4172 22148 4228 24668
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 4396 24500 4452 25564
rect 4732 25620 4788 25630
rect 4844 25620 4900 26348
rect 5180 26066 5236 27468
rect 5404 26404 5460 26414
rect 5404 26310 5460 26348
rect 5180 26014 5182 26066
rect 5234 26014 5236 26066
rect 5180 26002 5236 26014
rect 5180 25844 5236 25854
rect 5180 25730 5236 25788
rect 5180 25678 5182 25730
rect 5234 25678 5236 25730
rect 5180 25666 5236 25678
rect 4788 25564 4900 25620
rect 4956 25620 5012 25630
rect 4732 25554 4788 25564
rect 4956 25526 5012 25564
rect 4620 25284 4676 25294
rect 5068 25284 5124 25294
rect 4620 25282 5012 25284
rect 4620 25230 4622 25282
rect 4674 25230 5012 25282
rect 4620 25228 5012 25230
rect 4620 25218 4676 25228
rect 4284 24444 4452 24500
rect 4844 24724 4900 24734
rect 4284 23940 4340 24444
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4844 24164 4900 24668
rect 4732 24108 4900 24164
rect 4284 23874 4340 23884
rect 4508 24050 4564 24062
rect 4508 23998 4510 24050
rect 4562 23998 4564 24050
rect 4508 23380 4564 23998
rect 4732 23548 4788 24108
rect 4844 23940 4900 23950
rect 4844 23846 4900 23884
rect 4732 23492 4900 23548
rect 4396 23268 4452 23278
rect 4396 23154 4452 23212
rect 4396 23102 4398 23154
rect 4450 23102 4452 23154
rect 4396 23090 4452 23102
rect 4508 22932 4564 23324
rect 4284 22876 4564 22932
rect 4284 22370 4340 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22318 4286 22370
rect 4338 22318 4340 22370
rect 4284 22306 4340 22318
rect 4172 22092 4340 22148
rect 4172 21924 4228 21934
rect 4172 20914 4228 21868
rect 4172 20862 4174 20914
rect 4226 20862 4228 20914
rect 4172 20850 4228 20862
rect 3612 18676 3668 18686
rect 3500 18674 3668 18676
rect 3500 18622 3614 18674
rect 3666 18622 3668 18674
rect 3500 18620 3668 18622
rect 3612 18610 3668 18620
rect 3724 18674 3780 18686
rect 3724 18622 3726 18674
rect 3778 18622 3780 18674
rect 3500 18452 3556 18462
rect 3500 18358 3556 18396
rect 3724 18340 3780 18622
rect 3948 18340 4004 19180
rect 4172 20356 4228 20366
rect 4060 19124 4116 19134
rect 4060 19030 4116 19068
rect 3724 18284 3892 18340
rect 3948 18284 4116 18340
rect 3836 17892 3892 18284
rect 3948 17892 4004 17902
rect 3836 17890 4004 17892
rect 3836 17838 3950 17890
rect 4002 17838 4004 17890
rect 3836 17836 4004 17838
rect 3948 17826 4004 17836
rect 4060 17444 4116 18284
rect 4172 17668 4228 20300
rect 4284 20242 4340 22092
rect 4844 21700 4900 23492
rect 4956 22820 5012 25228
rect 5068 24948 5124 25228
rect 5068 24882 5124 24892
rect 5292 25284 5348 25294
rect 5068 23716 5124 23726
rect 5068 23154 5124 23660
rect 5292 23548 5348 25228
rect 5068 23102 5070 23154
rect 5122 23102 5124 23154
rect 5068 23090 5124 23102
rect 5180 23492 5348 23548
rect 5516 24724 5572 24734
rect 4956 22754 5012 22764
rect 4956 22372 5012 22382
rect 4956 22278 5012 22316
rect 4956 21700 5012 21710
rect 4844 21698 5012 21700
rect 4844 21646 4958 21698
rect 5010 21646 5012 21698
rect 4844 21644 5012 21646
rect 4508 21588 4564 21598
rect 4508 21494 4564 21532
rect 4956 21476 5012 21644
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4284 20190 4286 20242
rect 4338 20190 4340 20242
rect 4284 20178 4340 20190
rect 4396 21028 4452 21038
rect 4396 20020 4452 20972
rect 4620 20692 4676 20702
rect 4620 20598 4676 20636
rect 4956 20356 5012 21420
rect 4956 20290 5012 20300
rect 5068 20578 5124 20590
rect 5068 20526 5070 20578
rect 5122 20526 5124 20578
rect 4732 20132 4788 20142
rect 4172 17602 4228 17612
rect 4284 19964 4452 20020
rect 4508 20020 4564 20030
rect 4172 17444 4228 17454
rect 4060 17442 4228 17444
rect 4060 17390 4174 17442
rect 4226 17390 4228 17442
rect 4060 17388 4228 17390
rect 4172 17378 4228 17388
rect 3500 17220 3556 17230
rect 3276 16996 3332 17006
rect 3276 16210 3332 16940
rect 3388 16884 3444 16894
rect 3500 16884 3556 17164
rect 4284 17220 4340 19964
rect 4508 19926 4564 19964
rect 4732 19906 4788 20076
rect 4956 20020 5012 20030
rect 4732 19854 4734 19906
rect 4786 19854 4788 19906
rect 4732 19842 4788 19854
rect 4844 19964 4956 20020
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4620 19012 4676 19022
rect 4620 18918 4676 18956
rect 4844 18676 4900 19964
rect 4956 19926 5012 19964
rect 4956 19124 5012 19134
rect 4956 19030 5012 19068
rect 4956 18676 5012 18686
rect 4844 18674 5012 18676
rect 4844 18622 4958 18674
rect 5010 18622 5012 18674
rect 4844 18620 5012 18622
rect 4956 18610 5012 18620
rect 4620 18452 4676 18462
rect 4620 18358 4676 18396
rect 4844 18338 4900 18350
rect 4844 18286 4846 18338
rect 4898 18286 4900 18338
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4844 17890 4900 18286
rect 5068 18004 5124 20526
rect 5068 17938 5124 17948
rect 4844 17838 4846 17890
rect 4898 17838 4900 17890
rect 4620 17444 4676 17454
rect 4620 17350 4676 17388
rect 4284 17154 4340 17164
rect 3388 16882 3556 16884
rect 3388 16830 3390 16882
rect 3442 16830 3556 16882
rect 3388 16828 3556 16830
rect 3388 16818 3444 16828
rect 3276 16158 3278 16210
rect 3330 16158 3332 16210
rect 3276 16146 3332 16158
rect 3164 15820 3444 15876
rect 3052 15484 3220 15540
rect 2940 14578 2996 14588
rect 3052 15316 3108 15326
rect 2828 14466 2884 14476
rect 2492 14130 2548 14140
rect 2828 14306 2884 14318
rect 2828 14254 2830 14306
rect 2882 14254 2884 14306
rect 2716 13972 2772 13982
rect 2716 13878 2772 13916
rect 2380 13570 2436 13580
rect 2268 13470 2270 13522
rect 2322 13470 2324 13522
rect 2268 13458 2324 13470
rect 2828 13524 2884 14254
rect 2828 13458 2884 13468
rect 2940 14084 2996 14094
rect 1932 13188 1988 13198
rect 1932 13074 1988 13132
rect 1932 13022 1934 13074
rect 1986 13022 1988 13074
rect 1932 13010 1988 13022
rect 2380 12964 2436 12974
rect 2380 12870 2436 12908
rect 2716 12740 2772 12750
rect 2716 12738 2884 12740
rect 2716 12686 2718 12738
rect 2770 12686 2884 12738
rect 2716 12684 2884 12686
rect 2716 12674 2772 12684
rect 2828 12178 2884 12684
rect 2828 12126 2830 12178
rect 2882 12126 2884 12178
rect 2828 12114 2884 12126
rect 1932 12066 1988 12078
rect 1932 12014 1934 12066
rect 1986 12014 1988 12066
rect 1932 11508 1988 12014
rect 1932 11442 1988 11452
rect 2268 11396 2324 11406
rect 1820 11284 1876 11294
rect 2268 11284 2324 11340
rect 1820 11190 1876 11228
rect 2044 11282 2324 11284
rect 2044 11230 2270 11282
rect 2322 11230 2324 11282
rect 2044 11228 2324 11230
rect 2044 10500 2100 11228
rect 2268 11218 2324 11228
rect 2604 11284 2660 11294
rect 2604 11282 2884 11284
rect 2604 11230 2606 11282
rect 2658 11230 2884 11282
rect 2604 11228 2884 11230
rect 2156 10724 2212 10734
rect 2156 10630 2212 10668
rect 2268 10724 2324 10734
rect 2604 10724 2660 11228
rect 2828 10834 2884 11228
rect 2828 10782 2830 10834
rect 2882 10782 2884 10834
rect 2828 10770 2884 10782
rect 2268 10722 2660 10724
rect 2268 10670 2270 10722
rect 2322 10670 2660 10722
rect 2268 10668 2660 10670
rect 2268 10658 2324 10668
rect 2044 10444 2324 10500
rect 1932 10050 1988 10062
rect 1932 9998 1934 10050
rect 1986 9998 1988 10050
rect 1932 9938 1988 9998
rect 1932 9886 1934 9938
rect 1986 9886 1988 9938
rect 1932 9874 1988 9886
rect 1932 9156 1988 9166
rect 1932 9062 1988 9100
rect 1708 8372 2100 8428
rect 1820 8370 2100 8372
rect 1820 8318 1822 8370
rect 1874 8318 2100 8370
rect 1820 8316 2100 8318
rect 1820 8306 1876 8316
rect 2044 7588 2100 7598
rect 2044 7494 2100 7532
rect 1932 6916 1988 6926
rect 1932 6690 1988 6860
rect 2268 6916 2324 10444
rect 2380 9940 2436 9950
rect 2380 9846 2436 9884
rect 2828 9602 2884 9614
rect 2828 9550 2830 9602
rect 2882 9550 2884 9602
rect 2716 9492 2772 9502
rect 2380 8930 2436 8942
rect 2380 8878 2382 8930
rect 2434 8878 2436 8930
rect 2380 8260 2436 8878
rect 2716 8428 2772 9436
rect 2828 9044 2884 9550
rect 2828 8950 2884 8988
rect 2940 8818 2996 14028
rect 3052 13748 3108 15260
rect 3164 13970 3220 15484
rect 3388 15538 3444 15820
rect 3388 15486 3390 15538
rect 3442 15486 3444 15538
rect 3388 15474 3444 15486
rect 3164 13918 3166 13970
rect 3218 13918 3220 13970
rect 3164 13906 3220 13918
rect 3276 14306 3332 14318
rect 3276 14254 3278 14306
rect 3330 14254 3332 14306
rect 3052 13692 3220 13748
rect 2940 8766 2942 8818
rect 2994 8766 2996 8818
rect 2940 8754 2996 8766
rect 3052 13522 3108 13534
rect 3052 13470 3054 13522
rect 3106 13470 3108 13522
rect 2716 8372 2996 8428
rect 2828 8370 2996 8372
rect 2828 8318 2830 8370
rect 2882 8318 2996 8370
rect 2828 8316 2996 8318
rect 2828 8306 2884 8316
rect 2380 8204 2772 8260
rect 2380 8034 2436 8046
rect 2380 7982 2382 8034
rect 2434 7982 2436 8034
rect 2380 7924 2436 7982
rect 2380 7858 2436 7868
rect 2492 8036 2548 8046
rect 2492 7698 2548 7980
rect 2492 7646 2494 7698
rect 2546 7646 2548 7698
rect 2492 7634 2548 7646
rect 2268 6850 2324 6860
rect 1932 6638 1934 6690
rect 1986 6638 1988 6690
rect 1932 6626 1988 6638
rect 2604 6692 2660 6702
rect 2604 6598 2660 6636
rect 2380 6466 2436 6478
rect 2380 6414 2382 6466
rect 2434 6414 2436 6466
rect 2380 5908 2436 6414
rect 2716 6244 2772 8204
rect 2940 7700 2996 7710
rect 2940 7606 2996 7644
rect 2716 6178 2772 6188
rect 2828 5908 2884 5918
rect 2380 5906 2884 5908
rect 2380 5854 2830 5906
rect 2882 5854 2884 5906
rect 2380 5852 2884 5854
rect 2828 5842 2884 5852
rect 1932 5794 1988 5806
rect 1932 5742 1934 5794
rect 1986 5742 1988 5794
rect 1932 5460 1988 5742
rect 1932 5394 1988 5404
rect 2156 5236 2212 5246
rect 2156 5142 2212 5180
rect 2604 5124 2660 5134
rect 2604 4788 2660 5068
rect 2604 4732 2996 4788
rect 2380 4450 2436 4462
rect 2380 4398 2382 4450
rect 2434 4398 2436 4450
rect 2380 3556 2436 4398
rect 2716 4452 2772 4462
rect 2716 4358 2772 4396
rect 2828 3556 2884 3566
rect 2380 3554 2884 3556
rect 2380 3502 2830 3554
rect 2882 3502 2884 3554
rect 2380 3500 2884 3502
rect 2828 3490 2884 3500
rect 1596 2706 1652 2716
rect 1932 3442 1988 3454
rect 1932 3390 1934 3442
rect 1986 3390 1988 3442
rect 28 1876 84 1886
rect 28 800 84 1820
rect 1932 1876 1988 3390
rect 2940 2996 2996 4732
rect 2940 2930 2996 2940
rect 1932 1810 1988 1820
rect 3052 1316 3108 13470
rect 3164 11508 3220 13692
rect 3276 12964 3332 14254
rect 3500 13972 3556 16828
rect 4396 16994 4452 17006
rect 4396 16942 4398 16994
rect 4450 16942 4452 16994
rect 4396 16884 4452 16942
rect 4396 16818 4452 16828
rect 4620 16882 4676 16894
rect 4620 16830 4622 16882
rect 4674 16830 4676 16882
rect 3948 16772 4004 16782
rect 3836 16770 4004 16772
rect 3836 16718 3950 16770
rect 4002 16718 4004 16770
rect 3836 16716 4004 16718
rect 3612 16660 3668 16670
rect 3612 16210 3668 16604
rect 3612 16158 3614 16210
rect 3666 16158 3668 16210
rect 3612 15876 3668 16158
rect 3612 15810 3668 15820
rect 3836 15092 3892 16716
rect 3948 16706 4004 16716
rect 4060 16772 4116 16782
rect 3948 15540 4004 15550
rect 3948 15446 4004 15484
rect 3836 15026 3892 15036
rect 3612 14644 3668 14654
rect 4060 14644 4116 16716
rect 4620 16660 4676 16830
rect 4284 16604 4676 16660
rect 4172 16100 4228 16110
rect 4172 16006 4228 16044
rect 4284 15988 4340 16604
rect 4844 16548 4900 17838
rect 4956 17442 5012 17454
rect 5180 17444 5236 23492
rect 5516 21810 5572 24668
rect 5628 23380 5684 29148
rect 5740 28868 5796 29372
rect 5852 29316 5908 29326
rect 5852 29222 5908 29260
rect 5852 28868 5908 28878
rect 5740 28866 5908 28868
rect 5740 28814 5854 28866
rect 5906 28814 5908 28866
rect 5740 28812 5908 28814
rect 5852 28802 5908 28812
rect 5964 28754 6020 29932
rect 6188 29428 6244 29438
rect 5964 28702 5966 28754
rect 6018 28702 6020 28754
rect 5964 28690 6020 28702
rect 6076 29316 6132 29326
rect 6076 28420 6132 29260
rect 6076 28326 6132 28364
rect 5852 27748 5908 27758
rect 5852 27654 5908 27692
rect 6076 27188 6132 27198
rect 5740 27074 5796 27086
rect 5740 27022 5742 27074
rect 5794 27022 5796 27074
rect 5740 26964 5796 27022
rect 6076 27074 6132 27132
rect 6188 27186 6244 29372
rect 6524 29316 6580 29326
rect 6524 29222 6580 29260
rect 6300 28308 6356 28318
rect 6300 27860 6356 28252
rect 6524 28084 6580 28094
rect 6524 27990 6580 28028
rect 6636 27860 6692 30044
rect 6748 29204 6804 30268
rect 7084 30100 7140 30830
rect 7084 30034 7140 30044
rect 7084 29540 7140 29550
rect 6972 29428 7028 29438
rect 6972 29334 7028 29372
rect 6748 29148 7028 29204
rect 6300 27804 6468 27860
rect 6300 27636 6356 27646
rect 6300 27542 6356 27580
rect 6188 27134 6190 27186
rect 6242 27134 6244 27186
rect 6188 27122 6244 27134
rect 6076 27022 6078 27074
rect 6130 27022 6132 27074
rect 6076 27010 6132 27022
rect 6300 27076 6356 27086
rect 6412 27076 6468 27804
rect 6300 27074 6468 27076
rect 6300 27022 6302 27074
rect 6354 27022 6468 27074
rect 6300 27020 6468 27022
rect 6524 27804 6692 27860
rect 6860 27860 6916 27870
rect 5740 26898 5796 26908
rect 6300 26516 6356 27020
rect 6300 26450 6356 26460
rect 5740 26292 5796 26302
rect 5740 25284 5796 26236
rect 5852 26178 5908 26190
rect 5852 26126 5854 26178
rect 5906 26126 5908 26178
rect 5852 26066 5908 26126
rect 5852 26014 5854 26066
rect 5906 26014 5908 26066
rect 5852 26002 5908 26014
rect 6300 26178 6356 26190
rect 6300 26126 6302 26178
rect 6354 26126 6356 26178
rect 5740 25190 5796 25228
rect 6076 25620 6132 25630
rect 6076 25282 6132 25564
rect 6076 25230 6078 25282
rect 6130 25230 6132 25282
rect 6076 25060 6132 25230
rect 6076 24994 6132 25004
rect 5852 24722 5908 24734
rect 5852 24670 5854 24722
rect 5906 24670 5908 24722
rect 5740 23380 5796 23390
rect 5628 23378 5796 23380
rect 5628 23326 5742 23378
rect 5794 23326 5796 23378
rect 5628 23324 5796 23326
rect 5740 23314 5796 23324
rect 5852 22484 5908 24670
rect 5964 24612 6020 24622
rect 5964 24388 6020 24556
rect 6300 24612 6356 26126
rect 6300 24546 6356 24556
rect 6412 25172 6468 25182
rect 5964 24050 6020 24332
rect 5964 23998 5966 24050
rect 6018 23998 6020 24050
rect 5964 23986 6020 23998
rect 6188 24500 6244 24510
rect 6188 23828 6244 24444
rect 6188 23762 6244 23772
rect 6300 24164 6356 24174
rect 6188 23604 6244 23614
rect 5852 22418 5908 22428
rect 6076 23380 6132 23390
rect 5852 22260 5908 22270
rect 5852 22166 5908 22204
rect 5516 21758 5518 21810
rect 5570 21758 5572 21810
rect 5516 21746 5572 21758
rect 5852 21924 5908 21934
rect 5404 21586 5460 21598
rect 5404 21534 5406 21586
rect 5458 21534 5460 21586
rect 5404 21028 5460 21534
rect 5404 20962 5460 20972
rect 4956 17390 4958 17442
rect 5010 17390 5012 17442
rect 4956 17220 5012 17390
rect 4956 17154 5012 17164
rect 5068 17388 5236 17444
rect 5404 20244 5460 20254
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4620 16212 4676 16222
rect 4620 16118 4676 16156
rect 4172 15314 4228 15326
rect 4172 15262 4174 15314
rect 4226 15262 4228 15314
rect 4172 15204 4228 15262
rect 4172 15138 4228 15148
rect 4172 14980 4228 14990
rect 4172 14754 4228 14924
rect 4172 14702 4174 14754
rect 4226 14702 4228 14754
rect 4172 14690 4228 14702
rect 3612 14550 3668 14588
rect 3724 14642 4116 14644
rect 3724 14590 4062 14642
rect 4114 14590 4116 14642
rect 3724 14588 4116 14590
rect 3500 13906 3556 13916
rect 3612 13972 3668 13982
rect 3724 13972 3780 14588
rect 4060 14578 4116 14588
rect 3612 13970 3780 13972
rect 3612 13918 3614 13970
rect 3666 13918 3780 13970
rect 3612 13916 3780 13918
rect 3836 14308 3892 14318
rect 3612 13906 3668 13916
rect 3276 12898 3332 12908
rect 3612 12852 3668 12862
rect 3668 12796 3780 12852
rect 3612 12758 3668 12796
rect 3612 12066 3668 12078
rect 3612 12014 3614 12066
rect 3666 12014 3668 12066
rect 3164 11442 3220 11452
rect 3388 11508 3444 11518
rect 3164 11170 3220 11182
rect 3164 11118 3166 11170
rect 3218 11118 3220 11170
rect 3164 10724 3220 11118
rect 3164 10630 3220 10668
rect 3388 11172 3444 11452
rect 3500 11172 3556 11182
rect 3388 11170 3556 11172
rect 3388 11118 3502 11170
rect 3554 11118 3556 11170
rect 3388 11116 3556 11118
rect 3164 10500 3220 10510
rect 3164 10050 3220 10444
rect 3164 9998 3166 10050
rect 3218 9998 3220 10050
rect 3164 9986 3220 9998
rect 3276 10388 3332 10398
rect 3164 9602 3220 9614
rect 3164 9550 3166 9602
rect 3218 9550 3220 9602
rect 3164 9492 3220 9550
rect 3164 9426 3220 9436
rect 3276 9156 3332 10332
rect 3164 9100 3332 9156
rect 3164 8428 3220 9100
rect 3276 8930 3332 8942
rect 3276 8878 3278 8930
rect 3330 8878 3332 8930
rect 3276 8818 3332 8878
rect 3276 8766 3278 8818
rect 3330 8766 3332 8818
rect 3276 8754 3332 8766
rect 3164 8372 3332 8428
rect 3164 8034 3220 8046
rect 3164 7982 3166 8034
rect 3218 7982 3220 8034
rect 3164 7588 3220 7982
rect 3164 7522 3220 7532
rect 3164 6692 3220 6702
rect 3164 4564 3220 6636
rect 3276 6690 3332 8372
rect 3388 7700 3444 11116
rect 3500 11106 3556 11116
rect 3612 11060 3668 12014
rect 3612 10994 3668 11004
rect 3388 7634 3444 7644
rect 3500 9940 3556 9950
rect 3388 7362 3444 7374
rect 3388 7310 3390 7362
rect 3442 7310 3444 7362
rect 3388 7250 3444 7310
rect 3388 7198 3390 7250
rect 3442 7198 3444 7250
rect 3388 7186 3444 7198
rect 3276 6638 3278 6690
rect 3330 6638 3332 6690
rect 3276 6626 3332 6638
rect 3500 6020 3556 9884
rect 3724 9828 3780 12796
rect 3836 10834 3892 14252
rect 4172 13748 4228 13758
rect 4060 13636 4116 13646
rect 4172 13636 4228 13692
rect 4060 13634 4228 13636
rect 4060 13582 4062 13634
rect 4114 13582 4228 13634
rect 4060 13580 4228 13582
rect 4060 13570 4116 13580
rect 3948 12740 4004 12750
rect 3948 12738 4116 12740
rect 3948 12686 3950 12738
rect 4002 12686 4116 12738
rect 3948 12684 4116 12686
rect 3948 12674 4004 12684
rect 3836 10782 3838 10834
rect 3890 10782 3892 10834
rect 3836 10770 3892 10782
rect 3948 12516 4004 12526
rect 3724 9772 3892 9828
rect 3724 9604 3780 9642
rect 3724 9538 3780 9548
rect 3724 9380 3780 9390
rect 3724 9266 3780 9324
rect 3724 9214 3726 9266
rect 3778 9214 3780 9266
rect 3724 9202 3780 9214
rect 3836 8708 3892 9772
rect 3948 9716 4004 12460
rect 4060 12290 4116 12684
rect 4060 12238 4062 12290
rect 4114 12238 4116 12290
rect 4060 11396 4116 12238
rect 4060 11330 4116 11340
rect 4060 9940 4116 9950
rect 4060 9846 4116 9884
rect 3948 9268 4004 9660
rect 4060 9268 4116 9278
rect 3948 9266 4116 9268
rect 3948 9214 4062 9266
rect 4114 9214 4116 9266
rect 3948 9212 4116 9214
rect 3948 9044 4004 9212
rect 4060 9202 4116 9212
rect 3948 8978 4004 8988
rect 3612 8652 4116 8708
rect 3612 8370 3668 8652
rect 3612 8318 3614 8370
rect 3666 8318 3668 8370
rect 3612 8036 3668 8318
rect 3612 7970 3668 7980
rect 4060 8370 4116 8652
rect 4060 8318 4062 8370
rect 4114 8318 4116 8370
rect 3836 7364 3892 7374
rect 3836 7270 3892 7308
rect 3836 6916 3892 6926
rect 3724 6466 3780 6478
rect 3724 6414 3726 6466
rect 3778 6414 3780 6466
rect 3724 6356 3780 6414
rect 3724 6290 3780 6300
rect 3500 5964 3668 6020
rect 3500 5796 3556 5806
rect 3388 5236 3444 5246
rect 3500 5236 3556 5740
rect 3388 5234 3556 5236
rect 3388 5182 3390 5234
rect 3442 5182 3556 5234
rect 3388 5180 3556 5182
rect 3388 5170 3444 5180
rect 3612 5012 3668 5964
rect 3724 5236 3780 5246
rect 3836 5236 3892 6860
rect 4060 6244 4116 8318
rect 4172 7700 4228 13580
rect 4284 11396 4340 15932
rect 4844 15540 4900 16492
rect 5068 16324 5124 17388
rect 4844 15474 4900 15484
rect 4956 16268 5124 16324
rect 5180 16884 5236 16894
rect 4732 15428 4788 15438
rect 4732 15316 4788 15372
rect 4844 15316 4900 15326
rect 4732 15314 4900 15316
rect 4732 15262 4846 15314
rect 4898 15262 4900 15314
rect 4732 15260 4900 15262
rect 4844 15250 4900 15260
rect 4956 15148 5012 16268
rect 5068 16100 5124 16110
rect 5068 16006 5124 16044
rect 4844 15092 5012 15148
rect 5180 15428 5236 16828
rect 5404 16660 5460 20188
rect 5740 19908 5796 19918
rect 5740 19814 5796 19852
rect 5740 19460 5796 19470
rect 5852 19460 5908 21868
rect 6076 20914 6132 23324
rect 6188 23266 6244 23548
rect 6300 23548 6356 24108
rect 6412 23940 6468 25116
rect 6524 24388 6580 27804
rect 6860 27748 6916 27804
rect 6636 27692 6916 27748
rect 6636 27634 6692 27692
rect 6636 27582 6638 27634
rect 6690 27582 6692 27634
rect 6636 27570 6692 27582
rect 6860 26852 6916 26862
rect 6860 26516 6916 26796
rect 6860 26450 6916 26460
rect 6748 26292 6804 26302
rect 6748 26198 6804 26236
rect 6860 26178 6916 26190
rect 6860 26126 6862 26178
rect 6914 26126 6916 26178
rect 6636 25620 6692 25630
rect 6636 24610 6692 25564
rect 6860 25506 6916 26126
rect 6972 25732 7028 29148
rect 7084 28642 7140 29484
rect 7196 29316 7252 32732
rect 7644 32722 7700 32734
rect 7756 32674 7812 32686
rect 7756 32622 7758 32674
rect 7810 32622 7812 32674
rect 7308 32340 7364 32350
rect 7532 32340 7588 32350
rect 7756 32340 7812 32622
rect 7308 32338 7588 32340
rect 7308 32286 7310 32338
rect 7362 32286 7534 32338
rect 7586 32286 7588 32338
rect 7308 32284 7588 32286
rect 7308 32274 7364 32284
rect 7420 30324 7476 32284
rect 7532 32274 7588 32284
rect 7644 32284 7812 32340
rect 7532 31668 7588 31678
rect 7532 31108 7588 31612
rect 7532 31042 7588 31052
rect 7532 30884 7588 30922
rect 7644 30884 7700 32284
rect 7588 30828 7700 30884
rect 7756 31444 7812 31454
rect 7532 30818 7588 30828
rect 7420 30258 7476 30268
rect 7532 30660 7588 30670
rect 7532 29764 7588 30604
rect 7644 29988 7700 29998
rect 7644 29894 7700 29932
rect 7532 29708 7700 29764
rect 7644 29650 7700 29708
rect 7644 29598 7646 29650
rect 7698 29598 7700 29650
rect 7644 29586 7700 29598
rect 7532 29540 7588 29578
rect 7532 29474 7588 29484
rect 7196 29250 7252 29260
rect 7308 29426 7364 29438
rect 7308 29374 7310 29426
rect 7362 29374 7364 29426
rect 7308 29092 7364 29374
rect 7084 28590 7086 28642
rect 7138 28590 7140 28642
rect 7084 27300 7140 28590
rect 7196 29036 7364 29092
rect 7196 28532 7252 29036
rect 7756 28866 7812 31388
rect 7756 28814 7758 28866
rect 7810 28814 7812 28866
rect 7756 28802 7812 28814
rect 7308 28756 7364 28766
rect 7308 28642 7364 28700
rect 7868 28644 7924 33292
rect 7980 33346 8036 33628
rect 8204 33348 8260 36428
rect 8316 36418 8372 36428
rect 8316 35924 8372 35934
rect 8428 35924 8484 36764
rect 8316 35922 8484 35924
rect 8316 35870 8318 35922
rect 8370 35870 8484 35922
rect 8316 35868 8484 35870
rect 8316 35858 8372 35868
rect 8428 34802 8484 34814
rect 8428 34750 8430 34802
rect 8482 34750 8484 34802
rect 8428 34356 8484 34750
rect 8540 34468 8596 39340
rect 8652 38834 8708 38846
rect 8652 38782 8654 38834
rect 8706 38782 8708 38834
rect 8652 38612 8708 38782
rect 8652 38546 8708 38556
rect 8764 38164 8820 38174
rect 8876 38164 8932 43652
rect 9324 43652 9716 43708
rect 9772 45218 9828 45276
rect 9772 45166 9774 45218
rect 9826 45166 9828 45218
rect 8988 41972 9044 41982
rect 8988 41410 9044 41916
rect 8988 41358 8990 41410
rect 9042 41358 9044 41410
rect 8988 41300 9044 41358
rect 8988 41234 9044 41244
rect 8988 41076 9044 41086
rect 8988 39844 9044 41020
rect 9100 40292 9156 40302
rect 9100 40290 9268 40292
rect 9100 40238 9102 40290
rect 9154 40238 9268 40290
rect 9100 40236 9268 40238
rect 9100 40226 9156 40236
rect 9100 39844 9156 39854
rect 8988 39842 9156 39844
rect 8988 39790 9102 39842
rect 9154 39790 9156 39842
rect 8988 39788 9156 39790
rect 9100 39778 9156 39788
rect 8988 38948 9044 38958
rect 9212 38948 9268 40236
rect 8988 38946 9268 38948
rect 8988 38894 8990 38946
rect 9042 38894 9268 38946
rect 8988 38892 9268 38894
rect 8988 38724 9044 38892
rect 8988 38658 9044 38668
rect 8764 38162 8932 38164
rect 8764 38110 8766 38162
rect 8818 38110 8932 38162
rect 8764 38108 8932 38110
rect 8764 38098 8820 38108
rect 8876 38052 8932 38108
rect 8876 37986 8932 37996
rect 9100 37826 9156 37838
rect 9100 37774 9102 37826
rect 9154 37774 9156 37826
rect 9100 37716 9156 37774
rect 9100 37650 9156 37660
rect 8652 36932 8708 36942
rect 8652 35922 8708 36876
rect 9324 36820 9380 43652
rect 9660 43428 9716 43438
rect 9772 43428 9828 45166
rect 9660 43426 9828 43428
rect 9660 43374 9662 43426
rect 9714 43374 9828 43426
rect 9660 43372 9828 43374
rect 9660 43362 9716 43372
rect 9772 42980 9828 43372
rect 9772 42914 9828 42924
rect 9772 41972 9828 41982
rect 9772 41878 9828 41916
rect 9996 41970 10052 46956
rect 10108 46674 10164 47180
rect 10108 46622 10110 46674
rect 10162 46622 10164 46674
rect 10108 46610 10164 46622
rect 10332 46562 10388 47180
rect 10332 46510 10334 46562
rect 10386 46510 10388 46562
rect 10332 46498 10388 46510
rect 10108 46002 10164 46014
rect 10108 45950 10110 46002
rect 10162 45950 10164 46002
rect 10108 45108 10164 45950
rect 10108 45014 10164 45052
rect 10444 44434 10500 47404
rect 11452 47394 11508 47404
rect 11676 47460 11732 48190
rect 11788 47572 11844 48302
rect 12460 48356 12516 48366
rect 12460 48262 12516 48300
rect 12012 48244 12068 48254
rect 12012 48150 12068 48188
rect 11788 47506 11844 47516
rect 12460 47572 12516 47582
rect 11676 47394 11732 47404
rect 12236 47460 12292 47470
rect 12236 47366 12292 47404
rect 11788 47348 11844 47358
rect 10780 46562 10836 46574
rect 10780 46510 10782 46562
rect 10834 46510 10836 46562
rect 10780 46228 10836 46510
rect 10780 46162 10836 46172
rect 11788 46116 11844 47292
rect 12348 46116 12404 46126
rect 12460 46116 12516 47516
rect 12572 47234 12628 48972
rect 12796 49028 12852 49038
rect 12796 48934 12852 48972
rect 12684 48916 12740 48926
rect 12684 48822 12740 48860
rect 12908 48804 12964 48814
rect 12908 48710 12964 48748
rect 13132 48242 13188 48254
rect 13132 48190 13134 48242
rect 13186 48190 13188 48242
rect 13132 48020 13188 48190
rect 12908 47964 13132 48020
rect 12684 47572 12740 47582
rect 12684 47458 12740 47516
rect 12684 47406 12686 47458
rect 12738 47406 12740 47458
rect 12684 47394 12740 47406
rect 12908 47458 12964 47964
rect 13132 47954 13188 47964
rect 12908 47406 12910 47458
rect 12962 47406 12964 47458
rect 12572 47182 12574 47234
rect 12626 47182 12628 47234
rect 12572 47170 12628 47182
rect 12796 46900 12852 46910
rect 12908 46900 12964 47406
rect 12796 46898 12964 46900
rect 12796 46846 12798 46898
rect 12850 46846 12964 46898
rect 12796 46844 12964 46846
rect 13020 47348 13076 47358
rect 12796 46834 12852 46844
rect 11788 46060 12292 46116
rect 11116 45780 11172 45790
rect 10556 45666 10612 45678
rect 10556 45614 10558 45666
rect 10610 45614 10612 45666
rect 10556 45108 10612 45614
rect 11116 45668 11172 45724
rect 11116 45666 11284 45668
rect 11116 45614 11118 45666
rect 11170 45614 11284 45666
rect 11116 45612 11284 45614
rect 11116 45602 11172 45612
rect 10556 45042 10612 45052
rect 10444 44382 10446 44434
rect 10498 44382 10500 44434
rect 10444 44370 10500 44382
rect 10668 44996 10724 45006
rect 10556 44210 10612 44222
rect 10556 44158 10558 44210
rect 10610 44158 10612 44210
rect 10332 44098 10388 44110
rect 10332 44046 10334 44098
rect 10386 44046 10388 44098
rect 10220 43540 10276 43550
rect 10220 43446 10276 43484
rect 10332 42756 10388 44046
rect 10556 43652 10612 44158
rect 10556 43586 10612 43596
rect 10332 42690 10388 42700
rect 9996 41918 9998 41970
rect 10050 41918 10052 41970
rect 9996 41906 10052 41918
rect 9996 41748 10052 41758
rect 9436 41188 9492 41198
rect 9436 41094 9492 41132
rect 9884 41188 9940 41198
rect 9548 41076 9604 41086
rect 9548 40982 9604 41020
rect 9660 41074 9716 41086
rect 9660 41022 9662 41074
rect 9714 41022 9716 41074
rect 9660 40964 9716 41022
rect 9660 39620 9716 40908
rect 9884 40626 9940 41132
rect 9884 40574 9886 40626
rect 9938 40574 9940 40626
rect 9884 40562 9940 40574
rect 9996 40852 10052 41692
rect 10108 41748 10164 41758
rect 10108 41746 10500 41748
rect 10108 41694 10110 41746
rect 10162 41694 10500 41746
rect 10108 41692 10500 41694
rect 10108 41682 10164 41692
rect 10444 41298 10500 41692
rect 10668 41300 10724 44940
rect 10892 44994 10948 45006
rect 10892 44942 10894 44994
rect 10946 44942 10948 44994
rect 10892 44212 10948 44942
rect 11116 44212 11172 44222
rect 10892 44156 11116 44212
rect 11116 44118 11172 44156
rect 10892 43538 10948 43550
rect 10892 43486 10894 43538
rect 10946 43486 10948 43538
rect 10892 42532 10948 43486
rect 11116 43540 11172 43550
rect 11116 43446 11172 43484
rect 11116 43092 11172 43102
rect 11004 42756 11060 42794
rect 11004 42690 11060 42700
rect 11116 42754 11172 43036
rect 11116 42702 11118 42754
rect 11170 42702 11172 42754
rect 11004 42532 11060 42542
rect 10892 42530 11060 42532
rect 10892 42478 11006 42530
rect 11058 42478 11060 42530
rect 10892 42476 11060 42478
rect 11004 42466 11060 42476
rect 10780 41860 10836 41870
rect 10780 41766 10836 41804
rect 11116 41300 11172 42702
rect 10444 41246 10446 41298
rect 10498 41246 10500 41298
rect 10444 41234 10500 41246
rect 10556 41244 10724 41300
rect 11004 41244 11172 41300
rect 10220 41188 10276 41198
rect 10220 41094 10276 41132
rect 9996 40626 10052 40796
rect 9996 40574 9998 40626
rect 10050 40574 10052 40626
rect 9996 40562 10052 40574
rect 10220 40516 10276 40526
rect 9772 40402 9828 40414
rect 9772 40350 9774 40402
rect 9826 40350 9828 40402
rect 9772 39844 9828 40350
rect 9772 39778 9828 39788
rect 9548 39564 9716 39620
rect 9548 36932 9604 39564
rect 9884 39394 9940 39406
rect 9884 39342 9886 39394
rect 9938 39342 9940 39394
rect 9548 36866 9604 36876
rect 9660 38052 9716 38062
rect 9324 36754 9380 36764
rect 8764 36596 8820 36606
rect 9548 36596 9604 36606
rect 8764 36594 9604 36596
rect 8764 36542 8766 36594
rect 8818 36542 9550 36594
rect 9602 36542 9604 36594
rect 8764 36540 9604 36542
rect 8764 36530 8820 36540
rect 9548 36530 9604 36540
rect 8652 35870 8654 35922
rect 8706 35870 8708 35922
rect 8652 35858 8708 35870
rect 9436 36370 9492 36382
rect 9436 36318 9438 36370
rect 9490 36318 9492 36370
rect 9436 36260 9492 36318
rect 8876 35810 8932 35822
rect 8876 35758 8878 35810
rect 8930 35758 8932 35810
rect 8652 35700 8708 35710
rect 8652 35138 8708 35644
rect 8652 35086 8654 35138
rect 8706 35086 8708 35138
rect 8652 35074 8708 35086
rect 8876 35140 8932 35758
rect 8876 35074 8932 35084
rect 8988 35698 9044 35710
rect 8988 35646 8990 35698
rect 9042 35646 9044 35698
rect 8540 34412 8708 34468
rect 8316 33460 8372 33498
rect 8316 33394 8372 33404
rect 7980 33294 7982 33346
rect 8034 33294 8036 33346
rect 7980 33124 8036 33294
rect 7980 33058 8036 33068
rect 8092 33292 8260 33348
rect 8092 31220 8148 33292
rect 8316 33234 8372 33246
rect 8316 33182 8318 33234
rect 8370 33182 8372 33234
rect 8204 33124 8260 33134
rect 8204 33030 8260 33068
rect 8316 31444 8372 33182
rect 8428 33124 8484 34300
rect 8540 34018 8596 34030
rect 8540 33966 8542 34018
rect 8594 33966 8596 34018
rect 8540 33908 8596 33966
rect 8540 33842 8596 33852
rect 8428 33058 8484 33068
rect 8540 33234 8596 33246
rect 8540 33182 8542 33234
rect 8594 33182 8596 33234
rect 8428 32562 8484 32574
rect 8428 32510 8430 32562
rect 8482 32510 8484 32562
rect 8428 31668 8484 32510
rect 8540 31892 8596 33182
rect 8652 32786 8708 34412
rect 8988 34356 9044 35646
rect 9324 35588 9380 35598
rect 9436 35588 9492 36204
rect 9380 35532 9492 35588
rect 9548 36036 9604 36046
rect 9100 35028 9156 35038
rect 9100 34934 9156 34972
rect 8988 34290 9044 34300
rect 9100 34244 9156 34254
rect 9100 34150 9156 34188
rect 8652 32734 8654 32786
rect 8706 32734 8708 32786
rect 8652 32722 8708 32734
rect 8988 33796 9044 33806
rect 8764 32676 8820 32714
rect 8764 32610 8820 32620
rect 8876 32562 8932 32574
rect 8876 32510 8878 32562
rect 8930 32510 8932 32562
rect 8876 31948 8932 32510
rect 8540 31826 8596 31836
rect 8652 31892 8932 31948
rect 8428 31602 8484 31612
rect 8652 31778 8708 31892
rect 8988 31890 9044 33740
rect 8988 31838 8990 31890
rect 9042 31838 9044 31890
rect 8988 31826 9044 31838
rect 9100 33572 9156 33582
rect 8652 31726 8654 31778
rect 8706 31726 8708 31778
rect 8316 31378 8372 31388
rect 8092 31164 8260 31220
rect 8092 30996 8148 31006
rect 8092 30902 8148 30940
rect 7308 28590 7310 28642
rect 7362 28590 7364 28642
rect 7308 28578 7364 28590
rect 7756 28588 7924 28644
rect 8092 30772 8148 30782
rect 8092 30098 8148 30716
rect 8092 30046 8094 30098
rect 8146 30046 8148 30098
rect 7196 28438 7252 28476
rect 7196 27860 7252 27870
rect 7196 27766 7252 27804
rect 7420 27860 7476 27898
rect 7420 27794 7476 27804
rect 7644 27858 7700 27870
rect 7644 27806 7646 27858
rect 7698 27806 7700 27858
rect 7420 27636 7476 27646
rect 7196 27300 7252 27310
rect 7084 27298 7252 27300
rect 7084 27246 7198 27298
rect 7250 27246 7252 27298
rect 7084 27244 7252 27246
rect 7196 27234 7252 27244
rect 7308 27076 7364 27114
rect 7308 27010 7364 27020
rect 7420 26908 7476 27580
rect 7196 26852 7252 26862
rect 7196 26758 7252 26796
rect 7308 26852 7476 26908
rect 7084 26740 7140 26750
rect 7084 26402 7140 26684
rect 7084 26350 7086 26402
rect 7138 26350 7140 26402
rect 7084 26338 7140 26350
rect 7196 26628 7252 26638
rect 7196 26290 7252 26572
rect 7196 26238 7198 26290
rect 7250 26238 7252 26290
rect 7196 26226 7252 26238
rect 7196 25732 7252 25742
rect 6972 25730 7252 25732
rect 6972 25678 7198 25730
rect 7250 25678 7252 25730
rect 6972 25676 7252 25678
rect 7196 25666 7252 25676
rect 7308 25620 7364 26852
rect 7532 26516 7588 26526
rect 6860 25454 6862 25506
rect 6914 25454 6916 25506
rect 6860 25442 6916 25454
rect 7196 25506 7252 25518
rect 7196 25454 7198 25506
rect 7250 25454 7252 25506
rect 7308 25488 7364 25564
rect 7420 26180 7476 26190
rect 7420 25732 7476 26124
rect 7196 25396 7252 25454
rect 7196 25330 7252 25340
rect 7420 25396 7476 25676
rect 7532 25620 7588 26460
rect 7532 25554 7588 25564
rect 7420 25330 7476 25340
rect 6748 25284 6804 25294
rect 6748 25172 6804 25228
rect 6748 25116 7476 25172
rect 7308 24836 7364 24846
rect 6972 24724 7028 24734
rect 6972 24630 7028 24668
rect 7196 24724 7252 24734
rect 6636 24558 6638 24610
rect 6690 24558 6692 24610
rect 6636 24546 6692 24558
rect 7196 24500 7252 24668
rect 6972 24444 7252 24500
rect 6524 24332 6692 24388
rect 6524 23940 6580 23950
rect 6412 23938 6580 23940
rect 6412 23886 6526 23938
rect 6578 23886 6580 23938
rect 6412 23884 6580 23886
rect 6524 23874 6580 23884
rect 6300 23492 6468 23548
rect 6188 23214 6190 23266
rect 6242 23214 6244 23266
rect 6188 23202 6244 23214
rect 6300 22372 6356 22382
rect 6300 22278 6356 22316
rect 6412 22260 6468 23492
rect 6636 23156 6692 24332
rect 6972 24050 7028 24444
rect 6972 23998 6974 24050
rect 7026 23998 7028 24050
rect 6972 23986 7028 23998
rect 6748 23940 6804 23978
rect 6748 23874 6804 23884
rect 7196 23940 7252 23950
rect 7308 23940 7364 24780
rect 7196 23938 7364 23940
rect 7196 23886 7198 23938
rect 7250 23886 7364 23938
rect 7196 23884 7364 23886
rect 7420 23938 7476 25116
rect 7644 24836 7700 27806
rect 7756 27746 7812 28588
rect 7868 27860 7924 27870
rect 7868 27766 7924 27804
rect 7756 27694 7758 27746
rect 7810 27694 7812 27746
rect 7756 27682 7812 27694
rect 8092 27524 8148 30046
rect 8204 29988 8260 31164
rect 8316 31108 8372 31118
rect 8316 31014 8372 31052
rect 8540 30994 8596 31006
rect 8540 30942 8542 30994
rect 8594 30942 8596 30994
rect 8428 30884 8484 30894
rect 8428 30790 8484 30828
rect 8540 30660 8596 30942
rect 8540 30594 8596 30604
rect 8652 30996 8708 31726
rect 8876 31778 8932 31790
rect 8876 31726 8878 31778
rect 8930 31726 8932 31778
rect 8652 30434 8708 30940
rect 8652 30382 8654 30434
rect 8706 30382 8708 30434
rect 8652 30370 8708 30382
rect 8764 30994 8820 31006
rect 8764 30942 8766 30994
rect 8818 30942 8820 30994
rect 8764 30436 8820 30942
rect 8876 30660 8932 31726
rect 9100 31778 9156 33516
rect 9212 33348 9268 33358
rect 9212 33254 9268 33292
rect 9100 31726 9102 31778
rect 9154 31726 9156 31778
rect 9100 31714 9156 31726
rect 8876 30594 8932 30604
rect 8876 30436 8932 30446
rect 8764 30434 8932 30436
rect 8764 30382 8878 30434
rect 8930 30382 8932 30434
rect 8764 30380 8932 30382
rect 8876 30370 8932 30380
rect 8316 30324 8372 30334
rect 8316 30230 8372 30268
rect 9100 30324 9156 30334
rect 9100 30210 9156 30268
rect 9100 30158 9102 30210
rect 9154 30158 9156 30210
rect 9100 30146 9156 30158
rect 8204 29932 8596 29988
rect 8428 29652 8484 29662
rect 7644 24770 7700 24780
rect 7756 27468 8148 27524
rect 8204 29596 8428 29652
rect 7756 24724 7812 27468
rect 8092 27298 8148 27310
rect 8092 27246 8094 27298
rect 8146 27246 8148 27298
rect 8092 27186 8148 27246
rect 8092 27134 8094 27186
rect 8146 27134 8148 27186
rect 8092 27122 8148 27134
rect 7868 26628 7924 26638
rect 7868 26514 7924 26572
rect 7868 26462 7870 26514
rect 7922 26462 7924 26514
rect 7868 26450 7924 26462
rect 7980 26292 8036 26302
rect 7980 25508 8036 26236
rect 8204 25732 8260 29596
rect 8428 29558 8484 29596
rect 8540 29650 8596 29932
rect 8540 29598 8542 29650
rect 8594 29598 8596 29650
rect 8540 29586 8596 29598
rect 8652 29764 8708 29774
rect 8652 29650 8708 29708
rect 8652 29598 8654 29650
rect 8706 29598 8708 29650
rect 8652 29586 8708 29598
rect 9100 29426 9156 29438
rect 9100 29374 9102 29426
rect 9154 29374 9156 29426
rect 9100 28756 9156 29374
rect 9100 28690 9156 28700
rect 8428 28644 8484 28654
rect 8428 28082 8484 28588
rect 8652 28644 8708 28654
rect 8652 28550 8708 28588
rect 9324 28642 9380 35532
rect 9548 35026 9604 35980
rect 9548 34974 9550 35026
rect 9602 34974 9604 35026
rect 9548 34962 9604 34974
rect 9660 35812 9716 37996
rect 9884 37716 9940 39342
rect 9996 38724 10052 38734
rect 9996 38630 10052 38668
rect 10220 38500 10276 40460
rect 10332 39506 10388 39518
rect 10332 39454 10334 39506
rect 10386 39454 10388 39506
rect 10332 38724 10388 39454
rect 10556 38948 10612 41244
rect 10780 41186 10836 41198
rect 10780 41134 10782 41186
rect 10834 41134 10836 41186
rect 10668 41076 10724 41086
rect 10668 40982 10724 41020
rect 10780 40964 10836 41134
rect 10780 40898 10836 40908
rect 10668 39508 10724 39518
rect 10668 39414 10724 39452
rect 10332 38658 10388 38668
rect 10444 38892 10612 38948
rect 10220 38434 10276 38444
rect 10220 38276 10276 38286
rect 10220 38162 10276 38220
rect 10220 38110 10222 38162
rect 10274 38110 10276 38162
rect 10220 38098 10276 38110
rect 9884 37650 9940 37660
rect 10332 36820 10388 36830
rect 9772 36484 9828 36494
rect 9772 36390 9828 36428
rect 10220 36260 10276 36270
rect 10220 36166 10276 36204
rect 9996 36036 10052 36046
rect 9996 35922 10052 35980
rect 9996 35870 9998 35922
rect 10050 35870 10052 35922
rect 9996 35858 10052 35870
rect 9660 34244 9716 35756
rect 10220 35698 10276 35710
rect 10220 35646 10222 35698
rect 10274 35646 10276 35698
rect 10108 35586 10164 35598
rect 10108 35534 10110 35586
rect 10162 35534 10164 35586
rect 9884 35476 9940 35486
rect 9884 34468 9940 35420
rect 9996 35140 10052 35150
rect 10108 35140 10164 35534
rect 10220 35364 10276 35646
rect 10332 35698 10388 36764
rect 10444 36260 10500 38892
rect 10780 38834 10836 38846
rect 10780 38782 10782 38834
rect 10834 38782 10836 38834
rect 10556 38724 10612 38734
rect 10556 38164 10612 38668
rect 10556 37490 10612 38108
rect 10780 37828 10836 38782
rect 10892 38834 10948 38846
rect 10892 38782 10894 38834
rect 10946 38782 10948 38834
rect 10892 38052 10948 38782
rect 11004 38162 11060 41244
rect 11116 40290 11172 40302
rect 11116 40238 11118 40290
rect 11170 40238 11172 40290
rect 11116 40068 11172 40238
rect 11116 39396 11172 40012
rect 11116 39302 11172 39340
rect 11228 38500 11284 45612
rect 11788 45666 11844 45678
rect 11788 45614 11790 45666
rect 11842 45614 11844 45666
rect 11564 44996 11620 45006
rect 11788 44996 11844 45614
rect 12012 45220 12068 45230
rect 12012 45126 12068 45164
rect 11620 44940 11844 44996
rect 11564 44902 11620 44940
rect 11452 44100 11508 44110
rect 11340 42980 11396 42990
rect 11452 42980 11508 44044
rect 11900 44100 11956 44110
rect 11788 43652 11844 43662
rect 11788 43558 11844 43596
rect 11340 42978 11508 42980
rect 11340 42926 11342 42978
rect 11394 42926 11508 42978
rect 11340 42924 11508 42926
rect 11900 43538 11956 44044
rect 11900 43486 11902 43538
rect 11954 43486 11956 43538
rect 11900 42978 11956 43486
rect 12012 44098 12068 44110
rect 12012 44046 12014 44098
rect 12066 44046 12068 44098
rect 12012 43540 12068 44046
rect 12012 43474 12068 43484
rect 12124 43314 12180 43326
rect 12124 43262 12126 43314
rect 12178 43262 12180 43314
rect 12124 43092 12180 43262
rect 12124 43026 12180 43036
rect 11900 42926 11902 42978
rect 11954 42926 11956 42978
rect 11340 42914 11396 42924
rect 11900 42868 11956 42926
rect 12012 42868 12068 42878
rect 11900 42866 12068 42868
rect 11900 42814 12014 42866
rect 12066 42814 12068 42866
rect 11900 42812 12068 42814
rect 12012 42802 12068 42812
rect 11452 42756 11508 42766
rect 11340 41858 11396 41870
rect 11340 41806 11342 41858
rect 11394 41806 11396 41858
rect 11340 40516 11396 41806
rect 11340 40450 11396 40460
rect 11452 39060 11508 42700
rect 12236 42084 12292 46060
rect 12348 46114 12516 46116
rect 12348 46062 12350 46114
rect 12402 46062 12516 46114
rect 12348 46060 12516 46062
rect 12348 46050 12404 46060
rect 12684 45890 12740 45902
rect 12684 45838 12686 45890
rect 12738 45838 12740 45890
rect 12684 45332 12740 45838
rect 12908 45780 12964 45790
rect 12684 45266 12740 45276
rect 12796 45778 12964 45780
rect 12796 45726 12910 45778
rect 12962 45726 12964 45778
rect 12796 45724 12964 45726
rect 12572 45220 12628 45230
rect 12572 45126 12628 45164
rect 12796 45106 12852 45724
rect 12908 45714 12964 45724
rect 13020 45330 13076 47292
rect 13244 46562 13300 46574
rect 13244 46510 13246 46562
rect 13298 46510 13300 46562
rect 13020 45278 13022 45330
rect 13074 45278 13076 45330
rect 13020 45266 13076 45278
rect 13132 45332 13188 45342
rect 13244 45332 13300 46510
rect 13580 45892 13636 55020
rect 19836 54908 20100 54918
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 19836 54842 20100 54852
rect 19836 53340 20100 53350
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 19836 53274 20100 53284
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 13916 49812 13972 49822
rect 13916 49810 14084 49812
rect 13916 49758 13918 49810
rect 13970 49758 14084 49810
rect 13916 49756 14084 49758
rect 13916 49746 13972 49756
rect 13692 49588 13748 49598
rect 13692 49140 13748 49532
rect 13916 49364 13972 49374
rect 13916 49250 13972 49308
rect 13916 49198 13918 49250
rect 13970 49198 13972 49250
rect 13916 49186 13972 49198
rect 13692 49026 13748 49084
rect 13692 48974 13694 49026
rect 13746 48974 13748 49026
rect 13692 48962 13748 48974
rect 14028 49028 14084 49756
rect 20636 49810 20692 49822
rect 20636 49758 20638 49810
rect 20690 49758 20692 49810
rect 17612 49700 17668 49710
rect 14476 49364 14532 49374
rect 14140 49028 14196 49038
rect 14028 49026 14196 49028
rect 14028 48974 14142 49026
rect 14194 48974 14196 49026
rect 14028 48972 14196 48974
rect 13804 48804 13860 48814
rect 13804 48710 13860 48748
rect 14140 48354 14196 48972
rect 14140 48302 14142 48354
rect 14194 48302 14196 48354
rect 13804 48244 13860 48254
rect 13804 48150 13860 48188
rect 14028 48020 14084 48030
rect 13804 47460 13860 47470
rect 13804 47366 13860 47404
rect 14028 47460 14084 47964
rect 14028 47366 14084 47404
rect 13916 47348 13972 47358
rect 13916 47254 13972 47292
rect 14028 46676 14084 46686
rect 14028 46582 14084 46620
rect 13804 46562 13860 46574
rect 13804 46510 13806 46562
rect 13858 46510 13860 46562
rect 13692 46116 13748 46126
rect 13804 46116 13860 46510
rect 13692 46114 13860 46116
rect 13692 46062 13694 46114
rect 13746 46062 13860 46114
rect 13692 46060 13860 46062
rect 13692 46050 13748 46060
rect 13580 45836 13748 45892
rect 13188 45276 13300 45332
rect 13580 45332 13636 45342
rect 13132 45218 13188 45276
rect 13580 45238 13636 45276
rect 13132 45166 13134 45218
rect 13186 45166 13188 45218
rect 13132 45154 13188 45166
rect 12796 45054 12798 45106
rect 12850 45054 12852 45106
rect 12796 44996 12852 45054
rect 12796 44930 12852 44940
rect 13132 44212 13188 44222
rect 12908 44098 12964 44110
rect 12908 44046 12910 44098
rect 12962 44046 12964 44098
rect 12908 43708 12964 44046
rect 12796 43652 12964 43708
rect 13132 43708 13188 44156
rect 13580 43876 13636 43886
rect 13580 43708 13636 43820
rect 13132 43652 13636 43708
rect 12572 43540 12628 43550
rect 12796 43540 12852 43652
rect 13132 43650 13188 43652
rect 13132 43598 13134 43650
rect 13186 43598 13188 43650
rect 13132 43586 13188 43598
rect 13580 43650 13636 43652
rect 13580 43598 13582 43650
rect 13634 43598 13636 43650
rect 13580 43586 13636 43598
rect 12628 43484 12852 43540
rect 12572 43408 12628 43484
rect 12348 43314 12404 43326
rect 12348 43262 12350 43314
rect 12402 43262 12404 43314
rect 12348 42756 12404 43262
rect 12460 42978 12516 42990
rect 12460 42926 12462 42978
rect 12514 42926 12516 42978
rect 12460 42866 12516 42926
rect 12460 42814 12462 42866
rect 12514 42814 12516 42866
rect 12460 42802 12516 42814
rect 12684 42980 12740 42990
rect 12348 42690 12404 42700
rect 12348 42084 12404 42094
rect 12236 42082 12404 42084
rect 12236 42030 12350 42082
rect 12402 42030 12404 42082
rect 12236 42028 12404 42030
rect 12348 42018 12404 42028
rect 11676 40964 11732 40974
rect 11564 40962 11732 40964
rect 11564 40910 11678 40962
rect 11730 40910 11732 40962
rect 11564 40908 11732 40910
rect 11564 40402 11620 40908
rect 11676 40898 11732 40908
rect 12572 40962 12628 40974
rect 12572 40910 12574 40962
rect 12626 40910 12628 40962
rect 11564 40350 11566 40402
rect 11618 40350 11620 40402
rect 11564 40180 11620 40350
rect 11564 40114 11620 40124
rect 12124 40404 12180 40414
rect 12572 40404 12628 40910
rect 12124 40402 12628 40404
rect 12124 40350 12126 40402
rect 12178 40350 12628 40402
rect 12124 40348 12628 40350
rect 12124 40068 12180 40348
rect 12348 40180 12404 40190
rect 12348 40086 12404 40124
rect 12572 40178 12628 40190
rect 12572 40126 12574 40178
rect 12626 40126 12628 40178
rect 12124 40002 12180 40012
rect 12572 39956 12628 40126
rect 12572 39890 12628 39900
rect 11676 39394 11732 39406
rect 11676 39342 11678 39394
rect 11730 39342 11732 39394
rect 11564 39060 11620 39070
rect 11452 39058 11620 39060
rect 11452 39006 11566 39058
rect 11618 39006 11620 39058
rect 11452 39004 11620 39006
rect 11564 38994 11620 39004
rect 11340 38834 11396 38846
rect 11340 38782 11342 38834
rect 11394 38782 11396 38834
rect 11340 38724 11396 38782
rect 11396 38668 11508 38724
rect 11340 38658 11396 38668
rect 11228 38444 11396 38500
rect 11004 38110 11006 38162
rect 11058 38110 11060 38162
rect 11004 38098 11060 38110
rect 10892 37986 10948 37996
rect 11116 38052 11172 38062
rect 11004 37940 11060 37950
rect 11116 37940 11172 37996
rect 11004 37938 11172 37940
rect 11004 37886 11006 37938
rect 11058 37886 11172 37938
rect 11004 37884 11172 37886
rect 11228 37940 11284 37950
rect 11004 37874 11060 37884
rect 11228 37846 11284 37884
rect 10892 37828 10948 37838
rect 10780 37826 10948 37828
rect 10780 37774 10894 37826
rect 10946 37774 10948 37826
rect 10780 37772 10948 37774
rect 10892 37716 10948 37772
rect 10892 37650 10948 37660
rect 10556 37438 10558 37490
rect 10610 37438 10612 37490
rect 10556 37426 10612 37438
rect 11116 37604 11172 37614
rect 11004 37156 11060 37166
rect 11116 37156 11172 37548
rect 11004 37154 11172 37156
rect 11004 37102 11006 37154
rect 11058 37102 11172 37154
rect 11004 37100 11172 37102
rect 11004 37090 11060 37100
rect 10668 36260 10724 36270
rect 10444 36204 10612 36260
rect 10332 35646 10334 35698
rect 10386 35646 10388 35698
rect 10332 35634 10388 35646
rect 10220 35298 10276 35308
rect 10332 35140 10388 35150
rect 10108 35138 10388 35140
rect 10108 35086 10334 35138
rect 10386 35086 10388 35138
rect 10108 35084 10388 35086
rect 9996 34916 10052 35084
rect 10332 35074 10388 35084
rect 10108 34916 10164 34926
rect 9996 34914 10164 34916
rect 9996 34862 10110 34914
rect 10162 34862 10164 34914
rect 9996 34860 10164 34862
rect 10108 34850 10164 34860
rect 9884 34402 9940 34412
rect 10556 34354 10612 36204
rect 10668 35698 10724 36204
rect 10668 35646 10670 35698
rect 10722 35646 10724 35698
rect 10668 35634 10724 35646
rect 11004 36258 11060 36270
rect 11004 36206 11006 36258
rect 11058 36206 11060 36258
rect 11004 35364 11060 36206
rect 11004 35298 11060 35308
rect 10668 34916 10724 34926
rect 10668 34822 10724 34860
rect 10556 34302 10558 34354
rect 10610 34302 10612 34354
rect 10556 34290 10612 34302
rect 11004 34356 11060 34366
rect 11004 34262 11060 34300
rect 9660 34132 9716 34188
rect 9772 34132 9828 34142
rect 9660 34130 9828 34132
rect 9660 34078 9774 34130
rect 9826 34078 9828 34130
rect 9660 34076 9828 34078
rect 9772 34066 9828 34076
rect 9996 34130 10052 34142
rect 9996 34078 9998 34130
rect 10050 34078 10052 34130
rect 9660 33122 9716 33134
rect 9660 33070 9662 33122
rect 9714 33070 9716 33122
rect 9660 33012 9716 33070
rect 9660 32946 9716 32956
rect 9772 32676 9828 32686
rect 9660 32452 9716 32462
rect 9324 28590 9326 28642
rect 9378 28590 9380 28642
rect 8428 28030 8430 28082
rect 8482 28030 8484 28082
rect 8428 28018 8484 28030
rect 9100 28420 9156 28430
rect 8764 27860 8820 27870
rect 8764 27766 8820 27804
rect 8988 27748 9044 27758
rect 9100 27748 9156 28364
rect 9324 28308 9380 28590
rect 9324 28242 9380 28252
rect 9436 32450 9716 32452
rect 9436 32398 9662 32450
rect 9714 32398 9716 32450
rect 9436 32396 9716 32398
rect 8988 27746 9156 27748
rect 8988 27694 8990 27746
rect 9042 27694 9156 27746
rect 8988 27692 9156 27694
rect 8988 27682 9044 27692
rect 8428 27412 8484 27422
rect 8316 27300 8372 27338
rect 8316 27234 8372 27244
rect 8428 27186 8484 27356
rect 8428 27134 8430 27186
rect 8482 27134 8484 27186
rect 8316 27076 8372 27086
rect 8316 26516 8372 27020
rect 8428 26740 8484 27134
rect 9100 26964 9156 27692
rect 9436 27636 9492 32396
rect 9660 32386 9716 32396
rect 9772 31778 9828 32620
rect 9996 32564 10052 34078
rect 10108 34130 10164 34142
rect 10108 34078 10110 34130
rect 10162 34078 10164 34130
rect 10108 33460 10164 34078
rect 11116 34020 11172 37100
rect 11340 36932 11396 38444
rect 11452 38050 11508 38668
rect 11676 38668 11732 39342
rect 12124 39394 12180 39406
rect 12124 39342 12126 39394
rect 12178 39342 12180 39394
rect 12124 38948 12180 39342
rect 12572 39394 12628 39406
rect 12572 39342 12574 39394
rect 12626 39342 12628 39394
rect 12460 38948 12516 38958
rect 12180 38892 12292 38948
rect 12124 38882 12180 38892
rect 12124 38722 12180 38734
rect 12124 38670 12126 38722
rect 12178 38670 12180 38722
rect 11676 38612 12068 38668
rect 11452 37998 11454 38050
rect 11506 37998 11508 38050
rect 11452 37986 11508 37998
rect 11676 38500 11732 38510
rect 11676 37940 11732 38444
rect 11676 37884 11844 37940
rect 11788 37604 11844 37884
rect 11676 37548 11844 37604
rect 11676 37492 11732 37548
rect 11676 37426 11732 37436
rect 12012 37492 12068 38612
rect 12124 37716 12180 38670
rect 12236 38050 12292 38892
rect 12460 38854 12516 38892
rect 12572 38610 12628 39342
rect 12572 38558 12574 38610
rect 12626 38558 12628 38610
rect 12572 38546 12628 38558
rect 12684 38276 12740 42924
rect 12796 42196 12852 43484
rect 13692 42980 13748 45836
rect 14028 45890 14084 45902
rect 14028 45838 14030 45890
rect 14082 45838 14084 45890
rect 14028 45332 14084 45838
rect 14028 45266 14084 45276
rect 14028 44996 14084 45006
rect 14028 44902 14084 44940
rect 14140 43708 14196 48302
rect 14476 47682 14532 49308
rect 15820 49252 15876 49262
rect 15820 49138 15876 49196
rect 15820 49086 15822 49138
rect 15874 49086 15876 49138
rect 15820 49074 15876 49086
rect 17052 49252 17108 49262
rect 16044 49028 16100 49038
rect 16044 48934 16100 48972
rect 16940 49028 16996 49038
rect 16940 48934 16996 48972
rect 17052 48914 17108 49196
rect 17052 48862 17054 48914
rect 17106 48862 17108 48914
rect 17052 48850 17108 48862
rect 16380 48804 16436 48814
rect 16268 48802 16436 48804
rect 16268 48750 16382 48802
rect 16434 48750 16436 48802
rect 16268 48748 16436 48750
rect 16268 48468 16324 48748
rect 16380 48738 16436 48748
rect 17276 48802 17332 48814
rect 17276 48750 17278 48802
rect 17330 48750 17332 48802
rect 14476 47630 14478 47682
rect 14530 47630 14532 47682
rect 14364 46900 14420 46910
rect 14364 46806 14420 46844
rect 14476 46676 14532 47630
rect 15148 48130 15204 48142
rect 15148 48078 15150 48130
rect 15202 48078 15204 48130
rect 15148 47460 15204 48078
rect 15932 48132 15988 48142
rect 15932 48038 15988 48076
rect 16268 48130 16324 48412
rect 17276 48356 17332 48750
rect 17276 48290 17332 48300
rect 16268 48078 16270 48130
rect 16322 48078 16324 48130
rect 16268 48066 16324 48078
rect 16604 48244 16660 48254
rect 16604 47682 16660 48188
rect 16604 47630 16606 47682
rect 16658 47630 16660 47682
rect 16604 47618 16660 47630
rect 16716 47570 16772 47582
rect 16716 47518 16718 47570
rect 16770 47518 16772 47570
rect 14924 47234 14980 47246
rect 14924 47182 14926 47234
rect 14978 47182 14980 47234
rect 14924 47124 14980 47182
rect 14924 47058 14980 47068
rect 15148 47124 15204 47404
rect 15148 47058 15204 47068
rect 16268 47458 16324 47470
rect 16268 47406 16270 47458
rect 16322 47406 16324 47458
rect 16268 46900 16324 47406
rect 16268 46834 16324 46844
rect 14476 46610 14532 46620
rect 16716 46786 16772 47518
rect 17052 47236 17108 47246
rect 16828 46900 16884 46910
rect 16828 46806 16884 46844
rect 17052 46898 17108 47180
rect 17052 46846 17054 46898
rect 17106 46846 17108 46898
rect 17052 46834 17108 46846
rect 16716 46734 16718 46786
rect 16770 46734 16772 46786
rect 14252 45890 14308 45902
rect 14252 45838 14254 45890
rect 14306 45838 14308 45890
rect 14252 44996 14308 45838
rect 14700 45666 14756 45678
rect 14700 45614 14702 45666
rect 14754 45614 14756 45666
rect 14700 45332 14756 45614
rect 14252 44930 14308 44940
rect 14588 45108 14644 45118
rect 14252 44324 14308 44334
rect 14252 44230 14308 44268
rect 14364 43764 14420 43774
rect 13692 42914 13748 42924
rect 14028 43652 14196 43708
rect 14252 43652 14420 43708
rect 12796 42130 12852 42140
rect 12908 42868 12964 42878
rect 12908 41970 12964 42812
rect 13804 42868 13860 42878
rect 13804 42774 13860 42812
rect 13580 42756 13636 42766
rect 13244 42754 13636 42756
rect 13244 42702 13582 42754
rect 13634 42702 13636 42754
rect 13244 42700 13636 42702
rect 13020 42532 13076 42542
rect 13020 42530 13188 42532
rect 13020 42478 13022 42530
rect 13074 42478 13188 42530
rect 13020 42476 13188 42478
rect 13020 42466 13076 42476
rect 12908 41918 12910 41970
rect 12962 41918 12964 41970
rect 12908 41906 12964 41918
rect 13132 42084 13188 42476
rect 13132 41858 13188 42028
rect 13132 41806 13134 41858
rect 13186 41806 13188 41858
rect 13132 41794 13188 41806
rect 13020 40962 13076 40974
rect 13020 40910 13022 40962
rect 13074 40910 13076 40962
rect 13020 40292 13076 40910
rect 13244 40626 13300 42700
rect 13580 42690 13636 42700
rect 13692 42644 13748 42654
rect 13244 40574 13246 40626
rect 13298 40574 13300 40626
rect 13244 40562 13300 40574
rect 13356 42196 13412 42206
rect 13020 40226 13076 40236
rect 12796 40180 12852 40190
rect 12796 40086 12852 40124
rect 13020 39394 13076 39406
rect 13020 39342 13022 39394
rect 13074 39342 13076 39394
rect 13020 39284 13076 39342
rect 13020 39218 13076 39228
rect 13020 38836 13076 38846
rect 12236 37998 12238 38050
rect 12290 37998 12292 38050
rect 12236 37986 12292 37998
rect 12572 38220 12740 38276
rect 12796 38610 12852 38622
rect 12796 38558 12798 38610
rect 12850 38558 12852 38610
rect 12348 37828 12404 37838
rect 12348 37734 12404 37772
rect 12460 37826 12516 37838
rect 12460 37774 12462 37826
rect 12514 37774 12516 37826
rect 12236 37716 12292 37726
rect 12124 37660 12236 37716
rect 11452 37380 11508 37390
rect 11452 37286 11508 37324
rect 11900 37266 11956 37278
rect 11900 37214 11902 37266
rect 11954 37214 11956 37266
rect 11340 36876 11732 36932
rect 11564 36372 11620 36382
rect 11228 35812 11284 35822
rect 11228 35718 11284 35756
rect 11340 35474 11396 35486
rect 11340 35422 11342 35474
rect 11394 35422 11396 35474
rect 11340 35364 11396 35422
rect 11340 35298 11396 35308
rect 11564 35140 11620 36316
rect 11452 35084 11620 35140
rect 11340 34916 11396 34926
rect 11228 34244 11284 34254
rect 11228 34150 11284 34188
rect 11340 34242 11396 34860
rect 11340 34190 11342 34242
rect 11394 34190 11396 34242
rect 11340 34178 11396 34190
rect 11228 34020 11284 34030
rect 11116 33964 11228 34020
rect 10108 33394 10164 33404
rect 9772 31726 9774 31778
rect 9826 31726 9828 31778
rect 9660 30882 9716 30894
rect 9660 30830 9662 30882
rect 9714 30830 9716 30882
rect 9660 30772 9716 30830
rect 9660 30706 9716 30716
rect 9772 30434 9828 31726
rect 9884 32508 10052 32564
rect 10108 32564 10164 32574
rect 9884 30884 9940 32508
rect 10108 31444 10164 32508
rect 10220 32450 10276 32462
rect 10220 32398 10222 32450
rect 10274 32398 10276 32450
rect 10220 32004 10276 32398
rect 10892 32452 10948 32462
rect 10892 32358 10948 32396
rect 10220 31938 10276 31948
rect 10332 31892 10388 31902
rect 10332 31798 10388 31836
rect 10668 31892 10724 31902
rect 10332 31668 10388 31678
rect 10108 31378 10164 31388
rect 10220 31554 10276 31566
rect 10220 31502 10222 31554
rect 10274 31502 10276 31554
rect 9884 30818 9940 30828
rect 10220 30772 10276 31502
rect 10220 30706 10276 30716
rect 9772 30382 9774 30434
rect 9826 30382 9828 30434
rect 9772 30370 9828 30382
rect 9548 29988 9604 29998
rect 9548 29652 9604 29932
rect 10108 29986 10164 29998
rect 10108 29934 10110 29986
rect 10162 29934 10164 29986
rect 9548 29586 9604 29596
rect 9884 29764 9940 29774
rect 9436 27570 9492 27580
rect 9548 29204 9604 29214
rect 9324 26964 9380 26974
rect 9100 26962 9380 26964
rect 9100 26910 9326 26962
rect 9378 26910 9380 26962
rect 9100 26908 9380 26910
rect 8988 26852 9044 26862
rect 8988 26850 9156 26852
rect 8988 26798 8990 26850
rect 9042 26798 9156 26850
rect 8988 26796 9156 26798
rect 8988 26786 9044 26796
rect 8428 26674 8484 26684
rect 8316 26450 8372 26460
rect 8540 26516 8596 26526
rect 8428 26292 8484 26302
rect 8428 26198 8484 26236
rect 8204 25676 8372 25732
rect 7980 25376 8036 25452
rect 7756 24658 7812 24668
rect 7868 25172 7924 25182
rect 7868 24050 7924 25116
rect 7980 24164 8036 24174
rect 7980 24070 8036 24108
rect 7868 23998 7870 24050
rect 7922 23998 7924 24050
rect 7868 23986 7924 23998
rect 7420 23886 7422 23938
rect 7474 23886 7476 23938
rect 7196 23874 7252 23884
rect 7420 23874 7476 23886
rect 8204 23940 8260 23950
rect 7420 23714 7476 23726
rect 7420 23662 7422 23714
rect 7474 23662 7476 23714
rect 6636 23090 6692 23100
rect 6748 23604 6804 23614
rect 6748 22484 6804 23548
rect 6748 22418 6804 22428
rect 6860 23492 6916 23502
rect 6636 22372 6692 22382
rect 6636 22278 6692 22316
rect 6412 22258 6580 22260
rect 6412 22206 6414 22258
rect 6466 22206 6580 22258
rect 6412 22204 6580 22206
rect 6412 22194 6468 22204
rect 6524 21812 6580 22204
rect 6748 22148 6804 22158
rect 6636 21812 6692 21822
rect 6524 21810 6692 21812
rect 6524 21758 6638 21810
rect 6690 21758 6692 21810
rect 6524 21756 6692 21758
rect 6636 21746 6692 21756
rect 6076 20862 6078 20914
rect 6130 20862 6132 20914
rect 6076 20850 6132 20862
rect 6412 21700 6468 21710
rect 6412 21586 6468 21644
rect 6412 21534 6414 21586
rect 6466 21534 6468 21586
rect 6300 20804 6356 20814
rect 6300 20710 6356 20748
rect 6300 20580 6356 20590
rect 6076 19908 6132 19918
rect 6076 19906 6244 19908
rect 6076 19854 6078 19906
rect 6130 19854 6244 19906
rect 6076 19852 6244 19854
rect 6076 19842 6132 19852
rect 5740 19458 5908 19460
rect 5740 19406 5742 19458
rect 5794 19406 5908 19458
rect 5740 19404 5908 19406
rect 6076 19684 6132 19694
rect 5516 18564 5572 18574
rect 5516 18450 5572 18508
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 5516 18386 5572 18398
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4508 14532 4564 14542
rect 4508 14438 4564 14476
rect 4508 13972 4564 13982
rect 4508 13878 4564 13916
rect 4844 13860 4900 15092
rect 4956 14980 5012 14990
rect 4956 14754 5012 14924
rect 4956 14702 4958 14754
rect 5010 14702 5012 14754
rect 4956 14690 5012 14702
rect 4956 14308 5012 14318
rect 4956 14214 5012 14252
rect 5068 13860 5124 13870
rect 4844 13804 5012 13860
rect 4844 13634 4900 13646
rect 4844 13582 4846 13634
rect 4898 13582 4900 13634
rect 4844 13524 4900 13582
rect 4844 13458 4900 13468
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4620 13188 4676 13198
rect 4620 13074 4676 13132
rect 4620 13022 4622 13074
rect 4674 13022 4676 13074
rect 4620 12964 4676 13022
rect 4620 12898 4676 12908
rect 4396 12516 4452 12526
rect 4396 12402 4452 12460
rect 4396 12350 4398 12402
rect 4450 12350 4452 12402
rect 4396 12338 4452 12350
rect 4476 11788 4740 11798
rect 4956 11788 5012 13804
rect 5068 13524 5124 13804
rect 5180 13748 5236 15372
rect 5292 16604 5460 16660
rect 5516 18004 5572 18014
rect 5292 13972 5348 16604
rect 5516 16324 5572 17948
rect 5628 17556 5684 17566
rect 5628 17106 5684 17500
rect 5628 17054 5630 17106
rect 5682 17054 5684 17106
rect 5628 17042 5684 17054
rect 5740 16996 5796 19404
rect 5740 16864 5796 16940
rect 5852 19010 5908 19022
rect 5852 18958 5854 19010
rect 5906 18958 5908 19010
rect 5852 16772 5908 18958
rect 5964 19012 6020 19022
rect 5964 18674 6020 18956
rect 5964 18622 5966 18674
rect 6018 18622 6020 18674
rect 5964 18610 6020 18622
rect 6076 18674 6132 19628
rect 6076 18622 6078 18674
rect 6130 18622 6132 18674
rect 6076 18610 6132 18622
rect 6188 18564 6244 19852
rect 6188 18470 6244 18508
rect 6300 18228 6356 20524
rect 6412 20244 6468 21534
rect 6636 20804 6692 20814
rect 6636 20710 6692 20748
rect 6748 20580 6804 22092
rect 6748 20514 6804 20524
rect 6860 20244 6916 23436
rect 7196 23492 7252 23502
rect 7196 23044 7252 23436
rect 7084 22484 7140 22494
rect 6972 22372 7028 22382
rect 6972 22278 7028 22316
rect 6412 20178 6468 20188
rect 6748 20188 6916 20244
rect 6972 21476 7028 21486
rect 6636 19908 6692 19918
rect 6076 18172 6356 18228
rect 6524 19236 6580 19246
rect 6524 19124 6580 19180
rect 6636 19124 6692 19852
rect 6524 19122 6692 19124
rect 6524 19070 6638 19122
rect 6690 19070 6692 19122
rect 6524 19068 6692 19070
rect 5964 17444 6020 17454
rect 5964 17350 6020 17388
rect 6076 17220 6132 18172
rect 6524 17778 6580 19068
rect 6636 19058 6692 19068
rect 6524 17726 6526 17778
rect 6578 17726 6580 17778
rect 6524 17714 6580 17726
rect 6636 18004 6692 18014
rect 5852 16706 5908 16716
rect 5964 17164 6132 17220
rect 6412 17444 6468 17454
rect 5516 16268 5908 16324
rect 5740 15988 5796 15998
rect 5740 15894 5796 15932
rect 5404 15540 5460 15550
rect 5404 15446 5460 15484
rect 5740 15314 5796 15326
rect 5740 15262 5742 15314
rect 5794 15262 5796 15314
rect 5740 14420 5796 15262
rect 5852 14642 5908 16268
rect 5852 14590 5854 14642
rect 5906 14590 5908 14642
rect 5852 14578 5908 14590
rect 5740 14354 5796 14364
rect 5292 13906 5348 13916
rect 5740 13972 5796 13982
rect 5180 13682 5236 13692
rect 5740 13860 5796 13916
rect 5852 13860 5908 13870
rect 5740 13858 5908 13860
rect 5740 13806 5854 13858
rect 5906 13806 5908 13858
rect 5740 13804 5908 13806
rect 5292 13634 5348 13646
rect 5292 13582 5294 13634
rect 5346 13582 5348 13634
rect 5292 13524 5348 13582
rect 5068 13468 5236 13524
rect 5068 12738 5124 12750
rect 5068 12686 5070 12738
rect 5122 12686 5124 12738
rect 5068 12628 5124 12686
rect 5068 12562 5124 12572
rect 5068 12404 5124 12414
rect 5068 12290 5124 12348
rect 5068 12238 5070 12290
rect 5122 12238 5124 12290
rect 5068 12226 5124 12238
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11732 5012 11788
rect 5180 12178 5236 13468
rect 5292 12292 5348 13468
rect 5628 13300 5684 13310
rect 5292 12226 5348 12236
rect 5404 13188 5460 13198
rect 5180 12126 5182 12178
rect 5234 12126 5236 12178
rect 4844 11506 4900 11732
rect 4844 11454 4846 11506
rect 4898 11454 4900 11506
rect 4844 11442 4900 11454
rect 5068 11620 5124 11630
rect 4284 11330 4340 11340
rect 4956 11396 5012 11406
rect 4396 11172 4452 11182
rect 4284 10836 4340 10846
rect 4284 10742 4340 10780
rect 4396 10612 4452 11116
rect 4508 11170 4564 11182
rect 4508 11118 4510 11170
rect 4562 11118 4564 11170
rect 4508 10724 4564 11118
rect 4732 11170 4788 11182
rect 4732 11118 4734 11170
rect 4786 11118 4788 11170
rect 4620 11060 4676 11070
rect 4620 10834 4676 11004
rect 4620 10782 4622 10834
rect 4674 10782 4676 10834
rect 4620 10770 4676 10782
rect 4508 10658 4564 10668
rect 4284 10556 4452 10612
rect 4284 8932 4340 10556
rect 4732 10388 4788 11118
rect 4732 10322 4788 10332
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4956 10052 5012 11340
rect 4844 9996 5012 10052
rect 4620 9716 4676 9726
rect 4620 9622 4676 9660
rect 4508 8932 4564 8942
rect 4284 8930 4564 8932
rect 4284 8878 4510 8930
rect 4562 8878 4564 8930
rect 4284 8876 4564 8878
rect 4284 8484 4340 8876
rect 4508 8866 4564 8876
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4508 8484 4564 8494
rect 4284 8428 4452 8484
rect 4284 7700 4340 7710
rect 4172 7698 4340 7700
rect 4172 7646 4286 7698
rect 4338 7646 4340 7698
rect 4172 7644 4340 7646
rect 4284 7634 4340 7644
rect 4172 7252 4228 7262
rect 4172 6690 4228 7196
rect 4396 7252 4452 8428
rect 4396 7186 4452 7196
rect 4508 8370 4564 8428
rect 4508 8318 4510 8370
rect 4562 8318 4564 8370
rect 4508 7250 4564 8318
rect 4620 7700 4676 7710
rect 4844 7700 4900 9996
rect 4956 9828 5012 9838
rect 4956 9734 5012 9772
rect 5068 9266 5124 11564
rect 5180 10948 5236 12126
rect 5180 10892 5348 10948
rect 5180 10722 5236 10734
rect 5180 10670 5182 10722
rect 5234 10670 5236 10722
rect 5180 10612 5236 10670
rect 5180 10546 5236 10556
rect 5068 9214 5070 9266
rect 5122 9214 5124 9266
rect 5068 9202 5124 9214
rect 5068 9044 5124 9054
rect 5068 8370 5124 8988
rect 5068 8318 5070 8370
rect 5122 8318 5124 8370
rect 5068 8306 5124 8318
rect 5180 7700 5236 7710
rect 4620 7698 5236 7700
rect 4620 7646 4622 7698
rect 4674 7646 5182 7698
rect 5234 7646 5236 7698
rect 4620 7644 5236 7646
rect 4620 7588 4676 7644
rect 4620 7522 4676 7532
rect 4508 7198 4510 7250
rect 4562 7198 4564 7250
rect 4508 7186 4564 7198
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 5180 6804 5236 7644
rect 5180 6738 5236 6748
rect 4172 6638 4174 6690
rect 4226 6638 4228 6690
rect 4172 6626 4228 6638
rect 4508 6580 4564 6590
rect 4508 6486 4564 6524
rect 4956 6468 5012 6478
rect 4060 6188 4228 6244
rect 3948 6132 4004 6142
rect 3948 6038 4004 6076
rect 3724 5234 4116 5236
rect 3724 5182 3726 5234
rect 3778 5182 4116 5234
rect 3724 5180 4116 5182
rect 3724 5170 3780 5180
rect 3612 4956 3892 5012
rect 3276 4564 3332 4574
rect 3164 4562 3332 4564
rect 3164 4510 3278 4562
rect 3330 4510 3332 4562
rect 3164 4508 3332 4510
rect 3276 4498 3332 4508
rect 3612 4452 3668 4462
rect 3612 4358 3668 4396
rect 3836 3108 3892 4956
rect 4060 4562 4116 5180
rect 4060 4510 4062 4562
rect 4114 4510 4116 4562
rect 4060 4498 4116 4510
rect 3836 3042 3892 3052
rect 4172 2548 4228 6188
rect 4508 6132 4564 6142
rect 4508 6038 4564 6076
rect 4956 6130 5012 6412
rect 4956 6078 4958 6130
rect 5010 6078 5012 6130
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4508 5236 4564 5246
rect 4508 5142 4564 5180
rect 4956 5236 5012 6078
rect 4956 5104 5012 5180
rect 5068 6466 5124 6478
rect 5068 6414 5070 6466
rect 5122 6414 5124 6466
rect 4956 4676 5012 4686
rect 4620 4564 4676 4574
rect 4620 4470 4676 4508
rect 4956 4562 5012 4620
rect 4956 4510 4958 4562
rect 5010 4510 5012 4562
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 4956 3668 5012 4510
rect 5068 4340 5124 6414
rect 5292 6132 5348 10892
rect 5404 9716 5460 13132
rect 5628 12516 5684 13244
rect 5516 10610 5572 10622
rect 5516 10558 5518 10610
rect 5570 10558 5572 10610
rect 5516 10276 5572 10558
rect 5516 10210 5572 10220
rect 5404 9650 5460 9660
rect 5516 8930 5572 8942
rect 5516 8878 5518 8930
rect 5570 8878 5572 8930
rect 5516 8820 5572 8878
rect 5628 8932 5684 12460
rect 5740 11172 5796 13804
rect 5852 13794 5908 13804
rect 5964 13524 6020 17164
rect 6076 16994 6132 17006
rect 6076 16942 6078 16994
rect 6130 16942 6132 16994
rect 6076 15874 6132 16942
rect 6412 16884 6468 17388
rect 6412 16212 6468 16828
rect 6636 17220 6692 17948
rect 6524 16212 6580 16222
rect 6412 16210 6580 16212
rect 6412 16158 6526 16210
rect 6578 16158 6580 16210
rect 6412 16156 6580 16158
rect 6524 16146 6580 16156
rect 6076 15822 6078 15874
rect 6130 15822 6132 15874
rect 6076 15148 6132 15822
rect 6636 15988 6692 17164
rect 6636 15148 6692 15932
rect 6748 15538 6804 20188
rect 6860 19234 6916 19246
rect 6860 19182 6862 19234
rect 6914 19182 6916 19234
rect 6860 16548 6916 19182
rect 6972 18562 7028 21420
rect 6972 18510 6974 18562
rect 7026 18510 7028 18562
rect 6972 17668 7028 18510
rect 6972 17602 7028 17612
rect 7084 17556 7140 22428
rect 7196 21588 7252 22988
rect 7196 21522 7252 21532
rect 7308 23156 7364 23166
rect 7196 21362 7252 21374
rect 7196 21310 7198 21362
rect 7250 21310 7252 21362
rect 7196 20132 7252 21310
rect 7308 20244 7364 23100
rect 7420 22372 7476 23662
rect 7644 23716 7700 23726
rect 7532 23604 7588 23614
rect 7532 23380 7588 23548
rect 7532 23154 7588 23324
rect 7532 23102 7534 23154
rect 7586 23102 7588 23154
rect 7532 23090 7588 23102
rect 7532 22484 7588 22494
rect 7644 22484 7700 23660
rect 7756 23716 7812 23726
rect 7756 23714 7924 23716
rect 7756 23662 7758 23714
rect 7810 23662 7924 23714
rect 7756 23660 7924 23662
rect 7756 23650 7812 23660
rect 7868 23604 7924 23660
rect 7868 23538 7924 23548
rect 7532 22482 7700 22484
rect 7532 22430 7534 22482
rect 7586 22430 7700 22482
rect 7532 22428 7700 22430
rect 8204 23378 8260 23884
rect 8204 23326 8206 23378
rect 8258 23326 8260 23378
rect 7532 22418 7588 22428
rect 7420 22278 7476 22316
rect 7644 22148 7700 22158
rect 7644 22054 7700 22092
rect 8092 22146 8148 22158
rect 8092 22094 8094 22146
rect 8146 22094 8148 22146
rect 8092 21924 8148 22094
rect 8092 21858 8148 21868
rect 7980 21812 8036 21822
rect 7980 21718 8036 21756
rect 7868 21588 7924 21598
rect 7868 21494 7924 21532
rect 8092 21586 8148 21598
rect 8092 21534 8094 21586
rect 8146 21534 8148 21586
rect 7644 21476 7700 21486
rect 7644 21382 7700 21420
rect 7980 21476 8036 21486
rect 7308 20178 7364 20188
rect 7420 21362 7476 21374
rect 7420 21310 7422 21362
rect 7474 21310 7476 21362
rect 7196 19906 7252 20076
rect 7196 19854 7198 19906
rect 7250 19854 7252 19906
rect 7308 20020 7364 20030
rect 7420 20020 7476 21310
rect 7644 20802 7700 20814
rect 7644 20750 7646 20802
rect 7698 20750 7700 20802
rect 7364 19964 7476 20020
rect 7532 20690 7588 20702
rect 7532 20638 7534 20690
rect 7586 20638 7588 20690
rect 7532 20580 7588 20638
rect 7308 19888 7364 19964
rect 7196 19842 7252 19854
rect 7308 18452 7364 18462
rect 7532 18452 7588 20524
rect 7644 19906 7700 20750
rect 7980 20580 8036 21420
rect 8092 21364 8148 21534
rect 8092 21298 8148 21308
rect 7980 20514 8036 20524
rect 7644 19854 7646 19906
rect 7698 19854 7700 19906
rect 7644 19842 7700 19854
rect 7980 20244 8036 20254
rect 7756 19460 7812 19470
rect 7756 19346 7812 19404
rect 7756 19294 7758 19346
rect 7810 19294 7812 19346
rect 7756 19282 7812 19294
rect 7868 18564 7924 18574
rect 7868 18470 7924 18508
rect 7308 18450 7476 18452
rect 7308 18398 7310 18450
rect 7362 18398 7476 18450
rect 7308 18396 7476 18398
rect 7308 18386 7364 18396
rect 6860 16482 6916 16492
rect 6972 16996 7028 17006
rect 7084 16996 7140 17500
rect 6972 16994 7140 16996
rect 6972 16942 6974 16994
rect 7026 16942 7140 16994
rect 6972 16940 7140 16942
rect 7308 16996 7364 17006
rect 6748 15486 6750 15538
rect 6802 15486 6804 15538
rect 6748 15474 6804 15486
rect 6972 15428 7028 16940
rect 7308 16902 7364 16940
rect 7196 16884 7252 16894
rect 7196 16790 7252 16828
rect 7420 16772 7476 18396
rect 7532 18386 7588 18396
rect 7532 18116 7588 18126
rect 7532 17890 7588 18060
rect 7532 17838 7534 17890
rect 7586 17838 7588 17890
rect 7532 17826 7588 17838
rect 7644 17668 7700 17678
rect 7644 17574 7700 17612
rect 7532 17554 7588 17566
rect 7532 17502 7534 17554
rect 7586 17502 7588 17554
rect 7532 17444 7588 17502
rect 7868 17556 7924 17566
rect 7532 17388 7700 17444
rect 7308 16548 7364 16558
rect 7084 16212 7140 16222
rect 7084 15874 7140 16156
rect 7308 15986 7364 16492
rect 7420 16436 7476 16716
rect 7532 17108 7588 17118
rect 7532 16770 7588 17052
rect 7532 16718 7534 16770
rect 7586 16718 7588 16770
rect 7532 16706 7588 16718
rect 7420 16380 7588 16436
rect 7308 15934 7310 15986
rect 7362 15934 7364 15986
rect 7308 15922 7364 15934
rect 7420 15988 7476 15998
rect 7420 15894 7476 15932
rect 7532 15986 7588 16380
rect 7532 15934 7534 15986
rect 7586 15934 7588 15986
rect 7532 15922 7588 15934
rect 7084 15822 7086 15874
rect 7138 15822 7140 15874
rect 7084 15764 7140 15822
rect 7084 15708 7364 15764
rect 6972 15362 7028 15372
rect 7196 15428 7252 15438
rect 6076 15092 6356 15148
rect 6188 13860 6244 13870
rect 6188 13766 6244 13804
rect 5964 13458 6020 13468
rect 6076 12962 6132 12974
rect 6076 12910 6078 12962
rect 6130 12910 6132 12962
rect 5852 12852 5908 12862
rect 5852 12178 5908 12796
rect 6076 12402 6132 12910
rect 6076 12350 6078 12402
rect 6130 12350 6132 12402
rect 6076 12338 6132 12350
rect 6188 12964 6244 12974
rect 6188 12402 6244 12908
rect 6188 12350 6190 12402
rect 6242 12350 6244 12402
rect 5852 12126 5854 12178
rect 5906 12126 5908 12178
rect 5852 12114 5908 12126
rect 5964 12180 6020 12190
rect 5740 11170 5908 11172
rect 5740 11118 5742 11170
rect 5794 11118 5908 11170
rect 5740 11116 5908 11118
rect 5740 11106 5796 11116
rect 5852 9828 5908 11116
rect 5964 10050 6020 12124
rect 6188 11172 6244 12350
rect 6300 11732 6356 15092
rect 6524 15092 6692 15148
rect 6860 15314 6916 15326
rect 6860 15262 6862 15314
rect 6914 15262 6916 15314
rect 6860 15204 6916 15262
rect 7196 15314 7252 15372
rect 7196 15262 7198 15314
rect 7250 15262 7252 15314
rect 7196 15250 7252 15262
rect 6860 15138 6916 15148
rect 7308 15202 7364 15708
rect 7644 15540 7700 17388
rect 7756 16660 7812 16670
rect 7756 16566 7812 16604
rect 7868 16210 7924 17500
rect 7980 17332 8036 20188
rect 8092 20020 8148 20030
rect 8092 19348 8148 19964
rect 8092 19282 8148 19292
rect 8092 19012 8148 19022
rect 8092 18918 8148 18956
rect 8092 18562 8148 18574
rect 8092 18510 8094 18562
rect 8146 18510 8148 18562
rect 8092 17556 8148 18510
rect 8204 18116 8260 23326
rect 8316 20914 8372 25676
rect 8428 25506 8484 25518
rect 8428 25454 8430 25506
rect 8482 25454 8484 25506
rect 8428 25396 8484 25454
rect 8428 25330 8484 25340
rect 8428 24724 8484 24734
rect 8428 24630 8484 24668
rect 8540 24388 8596 26460
rect 8652 26066 8708 26078
rect 8652 26014 8654 26066
rect 8706 26014 8708 26066
rect 8652 25956 8708 26014
rect 8988 26068 9044 26078
rect 8988 25974 9044 26012
rect 8652 25890 8708 25900
rect 9100 25284 9156 26796
rect 9212 26516 9268 26908
rect 9324 26898 9380 26908
rect 9212 26450 9268 26460
rect 9324 26740 9380 26750
rect 9100 25218 9156 25228
rect 9324 25956 9380 26684
rect 9212 24724 9268 24734
rect 8540 23716 8596 24332
rect 9100 24610 9156 24622
rect 9100 24558 9102 24610
rect 9154 24558 9156 24610
rect 9100 24388 9156 24558
rect 9100 24322 9156 24332
rect 9100 24164 9156 24174
rect 8876 24052 8932 24062
rect 8876 23958 8932 23996
rect 8540 23378 8596 23660
rect 8540 23326 8542 23378
rect 8594 23326 8596 23378
rect 8540 23314 8596 23326
rect 8988 23044 9044 23054
rect 9100 23044 9156 24108
rect 8988 23042 9156 23044
rect 8988 22990 8990 23042
rect 9042 22990 9156 23042
rect 8988 22988 9156 22990
rect 8540 22596 8596 22606
rect 8540 22482 8596 22540
rect 8540 22430 8542 22482
rect 8594 22430 8596 22482
rect 8540 22418 8596 22430
rect 8316 20862 8318 20914
rect 8370 20862 8372 20914
rect 8316 20850 8372 20862
rect 8428 22372 8484 22382
rect 8428 20018 8484 22316
rect 8988 22036 9044 22988
rect 9100 22820 9156 22830
rect 9100 22260 9156 22764
rect 9212 22594 9268 24668
rect 9212 22542 9214 22594
rect 9266 22542 9268 22594
rect 9212 22530 9268 22542
rect 9324 22370 9380 25900
rect 9436 25282 9492 25294
rect 9436 25230 9438 25282
rect 9490 25230 9492 25282
rect 9436 24164 9492 25230
rect 9436 24098 9492 24108
rect 9324 22318 9326 22370
rect 9378 22318 9380 22370
rect 9324 22306 9380 22318
rect 9212 22260 9268 22270
rect 9100 22258 9268 22260
rect 9100 22206 9214 22258
rect 9266 22206 9268 22258
rect 9100 22204 9268 22206
rect 8988 21970 9044 21980
rect 9212 21924 9268 22204
rect 9212 21858 9268 21868
rect 8876 21588 8932 21598
rect 8428 19966 8430 20018
rect 8482 19966 8484 20018
rect 8428 19236 8484 19966
rect 8428 19170 8484 19180
rect 8540 20580 8596 20590
rect 8428 18676 8484 18686
rect 8204 18050 8260 18060
rect 8316 18450 8372 18462
rect 8316 18398 8318 18450
rect 8370 18398 8372 18450
rect 8204 17780 8260 17790
rect 8204 17686 8260 17724
rect 8092 17490 8148 17500
rect 8316 17554 8372 18398
rect 8316 17502 8318 17554
rect 8370 17502 8372 17554
rect 7980 17276 8260 17332
rect 7868 16158 7870 16210
rect 7922 16158 7924 16210
rect 7868 16146 7924 16158
rect 7644 15474 7700 15484
rect 7980 15988 8036 15998
rect 7308 15150 7310 15202
rect 7362 15150 7364 15202
rect 7308 15138 7364 15150
rect 7644 15204 7700 15214
rect 6748 15092 6804 15102
rect 6412 14420 6468 14430
rect 6412 12180 6468 14364
rect 6412 12114 6468 12124
rect 6300 11676 6468 11732
rect 6188 11106 6244 11116
rect 6300 10724 6356 10734
rect 6300 10630 6356 10668
rect 6412 10612 6468 11676
rect 6412 10480 6468 10556
rect 5964 9998 5966 10050
rect 6018 9998 6020 10050
rect 5964 9986 6020 9998
rect 6412 10276 6468 10286
rect 6412 9938 6468 10220
rect 6412 9886 6414 9938
rect 6466 9886 6468 9938
rect 6188 9828 6244 9838
rect 5852 9772 6020 9828
rect 5628 8866 5684 8876
rect 5516 8754 5572 8764
rect 5292 6038 5348 6076
rect 5404 7588 5460 7598
rect 5404 4676 5460 7532
rect 5516 7476 5572 7486
rect 5516 7382 5572 7420
rect 5740 6804 5796 6814
rect 5740 6710 5796 6748
rect 5516 6580 5572 6590
rect 5516 5908 5572 6524
rect 5740 6244 5796 6254
rect 5740 6130 5796 6188
rect 5740 6078 5742 6130
rect 5794 6078 5796 6130
rect 5740 6066 5796 6078
rect 5964 6132 6020 9772
rect 6076 7812 6132 7822
rect 6076 7474 6132 7756
rect 6076 7422 6078 7474
rect 6130 7422 6132 7474
rect 6076 6916 6132 7422
rect 6188 7476 6244 9772
rect 6300 9492 6356 9502
rect 6300 9266 6356 9436
rect 6300 9214 6302 9266
rect 6354 9214 6356 9266
rect 6300 9202 6356 9214
rect 6412 9268 6468 9886
rect 6524 9940 6580 15092
rect 6636 14418 6692 14430
rect 6636 14366 6638 14418
rect 6690 14366 6692 14418
rect 6636 13076 6692 14366
rect 6748 13970 6804 15036
rect 7644 14868 7700 15148
rect 7644 14812 7924 14868
rect 7420 14644 7476 14654
rect 6860 14532 6916 14542
rect 6860 14438 6916 14476
rect 7196 14532 7252 14542
rect 6972 14420 7028 14430
rect 7196 14420 7252 14476
rect 6972 14418 7252 14420
rect 6972 14366 6974 14418
rect 7026 14366 7252 14418
rect 6972 14364 7252 14366
rect 6972 14354 7028 14364
rect 6748 13918 6750 13970
rect 6802 13918 6804 13970
rect 6748 13906 6804 13918
rect 6860 14084 6916 14094
rect 6636 13010 6692 13020
rect 6524 9874 6580 9884
rect 6636 11396 6692 11406
rect 6412 9212 6580 9268
rect 6524 9156 6580 9212
rect 6524 9062 6580 9100
rect 6412 9044 6468 9054
rect 6412 8950 6468 8988
rect 6636 8428 6692 11340
rect 6748 10836 6804 10846
rect 6748 10500 6804 10780
rect 6748 10434 6804 10444
rect 6860 8596 6916 14028
rect 7420 14084 7476 14588
rect 7644 14644 7700 14654
rect 7644 14550 7700 14588
rect 7756 14530 7812 14542
rect 7756 14478 7758 14530
rect 7810 14478 7812 14530
rect 7532 14420 7588 14430
rect 7532 14326 7588 14364
rect 7420 14018 7476 14028
rect 7756 13972 7812 14478
rect 7756 13906 7812 13916
rect 7868 13858 7924 14812
rect 7868 13806 7870 13858
rect 7922 13806 7924 13858
rect 7756 13748 7812 13758
rect 7756 13654 7812 13692
rect 7308 13634 7364 13646
rect 7308 13582 7310 13634
rect 7362 13582 7364 13634
rect 7196 12964 7252 12974
rect 6972 12180 7028 12190
rect 6972 12086 7028 12124
rect 6972 11508 7028 11518
rect 7196 11508 7252 12908
rect 7308 12516 7364 13582
rect 7868 13300 7924 13806
rect 7868 13234 7924 13244
rect 7756 13076 7812 13086
rect 7756 12982 7812 13020
rect 7980 12516 8036 15932
rect 8092 15316 8148 15354
rect 8092 15250 8148 15260
rect 8092 14418 8148 14430
rect 8092 14366 8094 14418
rect 8146 14366 8148 14418
rect 8092 13972 8148 14366
rect 8092 13906 8148 13916
rect 8092 13746 8148 13758
rect 8092 13694 8094 13746
rect 8146 13694 8148 13746
rect 8092 12740 8148 13694
rect 8092 12674 8148 12684
rect 7308 12450 7364 12460
rect 7532 12460 8036 12516
rect 6972 11506 7252 11508
rect 6972 11454 6974 11506
rect 7026 11454 7252 11506
rect 6972 11452 7252 11454
rect 6972 9044 7028 11452
rect 7420 11396 7476 11406
rect 7420 11302 7476 11340
rect 7084 10612 7140 10622
rect 7084 9826 7140 10556
rect 7532 10052 7588 12460
rect 8092 12290 8148 12302
rect 8092 12238 8094 12290
rect 8146 12238 8148 12290
rect 7084 9774 7086 9826
rect 7138 9774 7140 9826
rect 7084 9762 7140 9774
rect 7196 9996 7588 10052
rect 7644 12180 7700 12190
rect 7196 9380 7252 9996
rect 7196 9266 7252 9324
rect 7196 9214 7198 9266
rect 7250 9214 7252 9266
rect 7196 9202 7252 9214
rect 7308 9828 7364 9838
rect 7308 9714 7364 9772
rect 7308 9662 7310 9714
rect 7362 9662 7364 9714
rect 6972 8988 7252 9044
rect 6860 8540 7028 8596
rect 6636 8372 6916 8428
rect 6860 8370 6916 8372
rect 6860 8318 6862 8370
rect 6914 8318 6916 8370
rect 6860 8306 6916 8318
rect 6412 8258 6468 8270
rect 6412 8206 6414 8258
rect 6466 8206 6468 8258
rect 6412 7700 6468 8206
rect 6748 8258 6804 8270
rect 6748 8206 6750 8258
rect 6802 8206 6804 8258
rect 6524 7700 6580 7710
rect 6412 7698 6580 7700
rect 6412 7646 6526 7698
rect 6578 7646 6580 7698
rect 6412 7644 6580 7646
rect 6524 7634 6580 7644
rect 6748 7700 6804 8206
rect 6748 7634 6804 7644
rect 6636 7588 6692 7598
rect 6636 7494 6692 7532
rect 6412 7476 6468 7486
rect 6188 7474 6468 7476
rect 6188 7422 6414 7474
rect 6466 7422 6468 7474
rect 6188 7420 6468 7422
rect 6412 7410 6468 7420
rect 6748 7476 6804 7486
rect 6076 6850 6132 6860
rect 6748 6914 6804 7420
rect 6748 6862 6750 6914
rect 6802 6862 6804 6914
rect 6748 6850 6804 6862
rect 6412 6690 6468 6702
rect 6412 6638 6414 6690
rect 6466 6638 6468 6690
rect 6300 6132 6356 6142
rect 5964 6130 6356 6132
rect 5964 6078 6302 6130
rect 6354 6078 6356 6130
rect 5964 6076 6356 6078
rect 6300 6066 6356 6076
rect 6412 6020 6468 6638
rect 6412 5954 6468 5964
rect 6524 6356 6580 6366
rect 5516 5852 5908 5908
rect 5404 4610 5460 4620
rect 5516 5236 5572 5246
rect 5516 4562 5572 5180
rect 5852 5236 5908 5852
rect 6524 5796 6580 6300
rect 6748 6132 6804 6142
rect 6972 6132 7028 8540
rect 7084 7476 7140 7486
rect 7084 7382 7140 7420
rect 6748 6130 7028 6132
rect 6748 6078 6750 6130
rect 6802 6078 7028 6130
rect 6748 6076 7028 6078
rect 7084 6692 7140 6702
rect 6748 6066 6804 6076
rect 6300 5740 6580 5796
rect 6636 6020 6692 6030
rect 5852 5104 5908 5180
rect 6188 5348 6244 5358
rect 5964 5124 6020 5134
rect 5516 4510 5518 4562
rect 5570 4510 5572 4562
rect 5516 4498 5572 4510
rect 5964 4562 6020 5068
rect 5964 4510 5966 4562
rect 6018 4510 6020 4562
rect 5964 4498 6020 4510
rect 5068 4274 5124 4284
rect 5068 3668 5124 3678
rect 4956 3666 5124 3668
rect 4956 3614 5070 3666
rect 5122 3614 5124 3666
rect 4956 3612 5124 3614
rect 5068 3602 5124 3612
rect 4620 3444 4676 3482
rect 4620 3378 4676 3388
rect 5404 3444 5460 3454
rect 4172 2482 4228 2492
rect 3052 1250 3108 1260
rect 5404 800 5460 3388
rect 5852 3444 5908 3482
rect 5852 3378 5908 3388
rect 6188 1540 6244 5292
rect 6300 5234 6356 5740
rect 6300 5182 6302 5234
rect 6354 5182 6356 5234
rect 6300 4564 6356 5182
rect 6636 4676 6692 5964
rect 7084 5796 7140 6636
rect 6860 5124 6916 5134
rect 6860 5030 6916 5068
rect 7084 4900 7140 5740
rect 7084 4834 7140 4844
rect 6636 4620 6916 4676
rect 6412 4564 6468 4574
rect 6300 4562 6468 4564
rect 6300 4510 6414 4562
rect 6466 4510 6468 4562
rect 6300 4508 6468 4510
rect 6412 4498 6468 4508
rect 6636 4564 6692 4620
rect 6636 4498 6692 4508
rect 6860 4562 6916 4620
rect 6860 4510 6862 4562
rect 6914 4510 6916 4562
rect 6860 4498 6916 4510
rect 7196 4228 7252 8988
rect 7308 8148 7364 9662
rect 7420 9714 7476 9726
rect 7420 9662 7422 9714
rect 7474 9662 7476 9714
rect 7420 9044 7476 9662
rect 7476 8988 7588 9044
rect 7420 8978 7476 8988
rect 7532 8260 7588 8988
rect 7644 8932 7700 12124
rect 7980 12066 8036 12078
rect 7980 12014 7982 12066
rect 8034 12014 8036 12066
rect 7980 11508 8036 12014
rect 7980 11442 8036 11452
rect 8092 12068 8148 12238
rect 8092 11060 8148 12012
rect 8204 11788 8260 17276
rect 8316 17220 8372 17502
rect 8316 17154 8372 17164
rect 8316 16996 8372 17006
rect 8316 13524 8372 16940
rect 8428 16436 8484 18620
rect 8540 18674 8596 20524
rect 8652 19236 8708 19246
rect 8652 19122 8708 19180
rect 8652 19070 8654 19122
rect 8706 19070 8708 19122
rect 8652 19058 8708 19070
rect 8540 18622 8542 18674
rect 8594 18622 8596 18674
rect 8540 18610 8596 18622
rect 8764 18564 8820 18574
rect 8540 18452 8596 18462
rect 8540 18358 8596 18396
rect 8652 18340 8708 18350
rect 8652 17892 8708 18284
rect 8652 17826 8708 17836
rect 8764 17666 8820 18508
rect 8764 17614 8766 17666
rect 8818 17614 8820 17666
rect 8540 17556 8596 17566
rect 8540 17462 8596 17500
rect 8764 17108 8820 17614
rect 8428 16370 8484 16380
rect 8540 17052 8820 17108
rect 8428 16212 8484 16222
rect 8428 16118 8484 16156
rect 8540 15148 8596 17052
rect 8652 16884 8708 16894
rect 8876 16884 8932 21532
rect 9100 21474 9156 21486
rect 9100 21422 9102 21474
rect 9154 21422 9156 21474
rect 8988 20804 9044 20814
rect 8988 20710 9044 20748
rect 9100 20468 9156 21422
rect 9100 20402 9156 20412
rect 8988 19906 9044 19918
rect 8988 19854 8990 19906
rect 9042 19854 9044 19906
rect 8988 19572 9044 19854
rect 9044 19516 9156 19572
rect 8988 19506 9044 19516
rect 8988 19236 9044 19246
rect 8988 19142 9044 19180
rect 8988 18788 9044 18798
rect 8988 18450 9044 18732
rect 9100 18676 9156 19516
rect 9100 18610 9156 18620
rect 8988 18398 8990 18450
rect 9042 18398 9044 18450
rect 8988 18386 9044 18398
rect 9100 18452 9156 18462
rect 9100 17106 9156 18396
rect 9212 18116 9268 18126
rect 9212 17890 9268 18060
rect 9548 18004 9604 29148
rect 9772 28308 9828 28318
rect 9772 28082 9828 28252
rect 9772 28030 9774 28082
rect 9826 28030 9828 28082
rect 9660 27636 9716 27646
rect 9660 26514 9716 27580
rect 9660 26462 9662 26514
rect 9714 26462 9716 26514
rect 9660 26450 9716 26462
rect 9772 25284 9828 28030
rect 9884 27412 9940 29708
rect 9996 29314 10052 29326
rect 9996 29262 9998 29314
rect 10050 29262 10052 29314
rect 9996 29204 10052 29262
rect 9996 29138 10052 29148
rect 9996 28756 10052 28766
rect 9996 28530 10052 28700
rect 9996 28478 9998 28530
rect 10050 28478 10052 28530
rect 9996 28466 10052 28478
rect 10108 28420 10164 29934
rect 10108 28354 10164 28364
rect 10220 28644 10276 28654
rect 10220 28084 10276 28588
rect 10220 27952 10276 28028
rect 9884 27074 9940 27356
rect 10332 27186 10388 31612
rect 10444 31556 10500 31566
rect 10444 31462 10500 31500
rect 10556 30884 10612 30894
rect 10556 30790 10612 30828
rect 10444 29986 10500 29998
rect 10444 29934 10446 29986
rect 10498 29934 10500 29986
rect 10444 29876 10500 29934
rect 10444 29810 10500 29820
rect 10668 29652 10724 31836
rect 10556 29596 10724 29652
rect 10780 31556 10836 31566
rect 10892 31556 10948 31566
rect 10836 31554 10948 31556
rect 10836 31502 10894 31554
rect 10946 31502 10948 31554
rect 10836 31500 10948 31502
rect 10780 30324 10836 31500
rect 10892 31490 10948 31500
rect 10892 31220 10948 31230
rect 10892 30660 10948 31164
rect 10892 30594 10948 30604
rect 11116 31108 11172 31118
rect 11116 30324 11172 31052
rect 10444 29428 10500 29438
rect 10444 29334 10500 29372
rect 10332 27134 10334 27186
rect 10386 27134 10388 27186
rect 10332 27122 10388 27134
rect 10444 29092 10500 29102
rect 10444 27860 10500 29036
rect 9884 27022 9886 27074
rect 9938 27022 9940 27074
rect 9884 27010 9940 27022
rect 10444 27074 10500 27804
rect 10444 27022 10446 27074
rect 10498 27022 10500 27074
rect 10444 27010 10500 27022
rect 10332 26964 10388 27002
rect 10332 26898 10388 26908
rect 10108 26850 10164 26862
rect 10108 26798 10110 26850
rect 10162 26798 10164 26850
rect 9884 26402 9940 26414
rect 9884 26350 9886 26402
rect 9938 26350 9940 26402
rect 9884 26068 9940 26350
rect 9884 26002 9940 26012
rect 9996 26290 10052 26302
rect 9996 26238 9998 26290
rect 10050 26238 10052 26290
rect 9996 25956 10052 26238
rect 9996 25890 10052 25900
rect 10108 25618 10164 26798
rect 10108 25566 10110 25618
rect 10162 25566 10164 25618
rect 10108 25554 10164 25566
rect 10444 26628 10500 26638
rect 10444 25508 10500 26572
rect 10556 26402 10612 29596
rect 10780 29540 10836 30268
rect 10668 29484 10836 29540
rect 10892 30268 11172 30324
rect 10892 29988 10948 30268
rect 10668 28980 10724 29484
rect 10780 29204 10836 29214
rect 10780 29110 10836 29148
rect 10668 28924 10836 28980
rect 10780 28532 10836 28924
rect 10892 28754 10948 29932
rect 11004 30098 11060 30110
rect 11004 30046 11006 30098
rect 11058 30046 11060 30098
rect 11004 29540 11060 30046
rect 11116 30100 11172 30110
rect 11116 30006 11172 30044
rect 11228 29876 11284 33964
rect 11452 31890 11508 35084
rect 11452 31838 11454 31890
rect 11506 31838 11508 31890
rect 11452 31826 11508 31838
rect 11564 34916 11620 34926
rect 11452 30882 11508 30894
rect 11452 30830 11454 30882
rect 11506 30830 11508 30882
rect 11452 30772 11508 30830
rect 11452 30706 11508 30716
rect 11004 29474 11060 29484
rect 11116 29820 11284 29876
rect 11340 29986 11396 29998
rect 11340 29934 11342 29986
rect 11394 29934 11396 29986
rect 11004 29316 11060 29326
rect 11004 29222 11060 29260
rect 10892 28702 10894 28754
rect 10946 28702 10948 28754
rect 10892 28690 10948 28702
rect 10780 28476 10948 28532
rect 10780 28196 10836 28206
rect 10668 28084 10724 28094
rect 10668 27990 10724 28028
rect 10556 26350 10558 26402
rect 10610 26350 10612 26402
rect 10556 26292 10612 26350
rect 10556 26226 10612 26236
rect 10780 26964 10836 28140
rect 10444 25452 10612 25508
rect 9996 25396 10052 25406
rect 9996 25302 10052 25340
rect 9772 25218 9828 25228
rect 10220 25284 10276 25294
rect 10220 25282 10388 25284
rect 10220 25230 10222 25282
rect 10274 25230 10388 25282
rect 10220 25228 10388 25230
rect 10220 25218 10276 25228
rect 9772 25060 9828 25070
rect 9660 23938 9716 23950
rect 9660 23886 9662 23938
rect 9714 23886 9716 23938
rect 9660 20018 9716 23886
rect 9772 23940 9828 25004
rect 10108 25060 10164 25070
rect 9884 24836 9940 24846
rect 9884 24742 9940 24780
rect 10108 24612 10164 25004
rect 10108 24518 10164 24556
rect 9772 23826 9828 23884
rect 10220 23938 10276 23950
rect 10220 23886 10222 23938
rect 10274 23886 10276 23938
rect 9772 23774 9774 23826
rect 9826 23774 9828 23826
rect 9772 23762 9828 23774
rect 9996 23828 10052 23838
rect 9660 19966 9662 20018
rect 9714 19966 9716 20018
rect 9660 19122 9716 19966
rect 9660 19070 9662 19122
rect 9714 19070 9716 19122
rect 9660 19058 9716 19070
rect 9772 21924 9828 21934
rect 9548 17938 9604 17948
rect 9772 18450 9828 21868
rect 9996 21476 10052 23772
rect 10220 23716 10276 23886
rect 10220 23650 10276 23660
rect 10220 22596 10276 22606
rect 10108 22370 10164 22382
rect 10108 22318 10110 22370
rect 10162 22318 10164 22370
rect 10108 22148 10164 22318
rect 10108 22082 10164 22092
rect 10108 21700 10164 21710
rect 10220 21700 10276 22540
rect 10332 22372 10388 25228
rect 10444 25282 10500 25294
rect 10444 25230 10446 25282
rect 10498 25230 10500 25282
rect 10444 25172 10500 25230
rect 10444 25106 10500 25116
rect 10444 24724 10500 24762
rect 10444 24658 10500 24668
rect 10556 24612 10612 25452
rect 10780 24722 10836 26908
rect 10892 26514 10948 28476
rect 11116 28420 11172 29820
rect 11228 29652 11284 29662
rect 11228 28866 11284 29596
rect 11228 28814 11230 28866
rect 11282 28814 11284 28866
rect 11228 28802 11284 28814
rect 11340 28756 11396 29934
rect 11564 29652 11620 34860
rect 11676 32788 11732 36876
rect 11900 36484 11956 37214
rect 11900 36418 11956 36428
rect 12012 36260 12068 37436
rect 12236 37490 12292 37660
rect 12460 37604 12516 37774
rect 12460 37538 12516 37548
rect 12236 37438 12238 37490
rect 12290 37438 12292 37490
rect 12236 37426 12292 37438
rect 12460 36260 12516 36270
rect 12012 36258 12516 36260
rect 12012 36206 12014 36258
rect 12066 36206 12462 36258
rect 12514 36206 12516 36258
rect 12012 36204 12516 36206
rect 11788 35812 11844 35822
rect 11788 35718 11844 35756
rect 11788 34914 11844 34926
rect 11788 34862 11790 34914
rect 11842 34862 11844 34914
rect 11788 34244 11844 34862
rect 12012 34916 12068 36204
rect 12460 36194 12516 36204
rect 12572 36036 12628 38220
rect 12684 38052 12740 38062
rect 12796 38052 12852 38558
rect 12684 38050 12852 38052
rect 12684 37998 12686 38050
rect 12738 37998 12852 38050
rect 12684 37996 12852 37998
rect 12908 38050 12964 38062
rect 12908 37998 12910 38050
rect 12962 37998 12964 38050
rect 12684 36260 12740 37996
rect 12908 37716 12964 37998
rect 12908 37650 12964 37660
rect 12908 37154 12964 37166
rect 12908 37102 12910 37154
rect 12962 37102 12964 37154
rect 12908 37044 12964 37102
rect 12908 36978 12964 36988
rect 12908 36260 12964 36270
rect 12684 36204 12908 36260
rect 12908 36166 12964 36204
rect 12236 35980 12628 36036
rect 12236 35026 12292 35980
rect 12460 35812 12516 35822
rect 12908 35812 12964 35822
rect 13020 35812 13076 38780
rect 13356 38668 13412 42140
rect 13692 41298 13748 42588
rect 13916 42532 13972 42542
rect 13804 42530 13972 42532
rect 13804 42478 13918 42530
rect 13970 42478 13972 42530
rect 13804 42476 13972 42478
rect 13804 41412 13860 42476
rect 13916 42466 13972 42476
rect 14028 42194 14084 43652
rect 14252 43650 14308 43652
rect 14252 43598 14254 43650
rect 14306 43598 14308 43650
rect 14252 43586 14308 43598
rect 14252 43428 14308 43438
rect 14140 43314 14196 43326
rect 14140 43262 14142 43314
rect 14194 43262 14196 43314
rect 14140 42644 14196 43262
rect 14252 43092 14308 43372
rect 14252 43026 14308 43036
rect 14140 42550 14196 42588
rect 14028 42142 14030 42194
rect 14082 42142 14084 42194
rect 14028 42130 14084 42142
rect 13916 42084 13972 42094
rect 13916 41990 13972 42028
rect 14252 41970 14308 41982
rect 14252 41918 14254 41970
rect 14306 41918 14308 41970
rect 13916 41412 13972 41422
rect 13804 41410 14084 41412
rect 13804 41358 13918 41410
rect 13970 41358 14084 41410
rect 13804 41356 14084 41358
rect 13916 41346 13972 41356
rect 13692 41246 13694 41298
rect 13746 41246 13748 41298
rect 13692 41234 13748 41246
rect 13692 40292 13748 40302
rect 13692 39620 13748 40236
rect 13804 40180 13860 40190
rect 13804 40086 13860 40124
rect 13916 40178 13972 40190
rect 13916 40126 13918 40178
rect 13970 40126 13972 40178
rect 13916 39956 13972 40126
rect 13916 39890 13972 39900
rect 13916 39732 13972 39742
rect 14028 39732 14084 41356
rect 14252 41410 14308 41918
rect 14252 41358 14254 41410
rect 14306 41358 14308 41410
rect 14252 41346 14308 41358
rect 14476 41970 14532 41982
rect 14476 41918 14478 41970
rect 14530 41918 14532 41970
rect 14476 40514 14532 41918
rect 14476 40462 14478 40514
rect 14530 40462 14532 40514
rect 14476 40450 14532 40462
rect 14140 40292 14196 40302
rect 14140 40198 14196 40236
rect 14364 40178 14420 40190
rect 14364 40126 14366 40178
rect 14418 40126 14420 40178
rect 13916 39730 14084 39732
rect 13916 39678 13918 39730
rect 13970 39678 14084 39730
rect 13916 39676 14084 39678
rect 14140 39956 14196 39966
rect 13916 39666 13972 39676
rect 13804 39620 13860 39630
rect 13692 39618 13860 39620
rect 13692 39566 13806 39618
rect 13858 39566 13860 39618
rect 13692 39564 13860 39566
rect 13804 39554 13860 39564
rect 14140 39618 14196 39900
rect 14140 39566 14142 39618
rect 14194 39566 14196 39618
rect 14028 39396 14084 39406
rect 14028 39302 14084 39340
rect 14028 38834 14084 38846
rect 14028 38782 14030 38834
rect 14082 38782 14084 38834
rect 13244 38612 13412 38668
rect 13468 38722 13524 38734
rect 13468 38670 13470 38722
rect 13522 38670 13524 38722
rect 13132 37268 13188 37278
rect 13132 35922 13188 37212
rect 13244 36932 13300 38612
rect 13244 36866 13300 36876
rect 13356 37266 13412 37278
rect 13356 37214 13358 37266
rect 13410 37214 13412 37266
rect 13356 37044 13412 37214
rect 13468 37268 13524 38670
rect 13916 38724 13972 38734
rect 13916 38630 13972 38668
rect 14028 38388 14084 38782
rect 14028 38322 14084 38332
rect 14028 38050 14084 38062
rect 14028 37998 14030 38050
rect 14082 37998 14084 38050
rect 13916 37492 13972 37502
rect 14028 37492 14084 37998
rect 13916 37490 14084 37492
rect 13916 37438 13918 37490
rect 13970 37438 14084 37490
rect 13916 37436 14084 37438
rect 13916 37426 13972 37436
rect 13804 37380 13860 37390
rect 13804 37286 13860 37324
rect 13580 37268 13636 37278
rect 13468 37266 13636 37268
rect 13468 37214 13582 37266
rect 13634 37214 13636 37266
rect 13468 37212 13636 37214
rect 13132 35870 13134 35922
rect 13186 35870 13188 35922
rect 13132 35858 13188 35870
rect 12460 35810 13076 35812
rect 12460 35758 12462 35810
rect 12514 35758 12910 35810
rect 12962 35758 13076 35810
rect 12460 35756 13076 35758
rect 12460 35746 12516 35756
rect 12908 35746 12964 35756
rect 13244 35588 13300 35598
rect 13244 35494 13300 35532
rect 12236 34974 12238 35026
rect 12290 34974 12292 35026
rect 12236 34962 12292 34974
rect 12012 34850 12068 34860
rect 12796 34916 12852 34926
rect 12012 34468 12068 34478
rect 11900 34244 11956 34254
rect 11788 34188 11900 34244
rect 11676 32722 11732 32732
rect 11788 33684 11844 33694
rect 11788 32674 11844 33628
rect 11788 32622 11790 32674
rect 11842 32622 11844 32674
rect 11788 32610 11844 32622
rect 11900 33236 11956 34188
rect 12012 33684 12068 34412
rect 12796 34020 12852 34860
rect 13244 34804 13300 34814
rect 12012 33618 12068 33628
rect 12572 34018 12852 34020
rect 12572 33966 12798 34018
rect 12850 33966 12852 34018
rect 12572 33964 12852 33966
rect 11900 31218 11956 33180
rect 12460 33236 12516 33246
rect 12460 33142 12516 33180
rect 12124 33122 12180 33134
rect 12124 33070 12126 33122
rect 12178 33070 12180 33122
rect 12124 31778 12180 33070
rect 12348 33124 12404 33134
rect 12348 33030 12404 33068
rect 12460 32564 12516 32574
rect 12460 32470 12516 32508
rect 12348 31892 12404 31902
rect 12348 31798 12404 31836
rect 12124 31726 12126 31778
rect 12178 31726 12180 31778
rect 12124 31714 12180 31726
rect 11900 31166 11902 31218
rect 11954 31166 11956 31218
rect 11900 31154 11956 31166
rect 12236 30996 12292 31006
rect 12236 30902 12292 30940
rect 11788 30884 11844 30894
rect 11564 29586 11620 29596
rect 11676 30212 11732 30222
rect 11788 30212 11844 30828
rect 11676 30210 11844 30212
rect 11676 30158 11678 30210
rect 11730 30158 11844 30210
rect 11676 30156 11844 30158
rect 12012 30660 12068 30670
rect 11676 30100 11732 30156
rect 11676 29538 11732 30044
rect 11676 29486 11678 29538
rect 11730 29486 11732 29538
rect 11676 29474 11732 29486
rect 11900 29764 11956 29774
rect 11564 29428 11620 29438
rect 11564 29334 11620 29372
rect 11340 28690 11396 28700
rect 11228 28644 11284 28654
rect 11228 28550 11284 28588
rect 11676 28532 11732 28542
rect 11116 28364 11396 28420
rect 11228 27300 11284 27310
rect 11116 26964 11172 27002
rect 11116 26898 11172 26908
rect 11228 26740 11284 27244
rect 11228 26674 11284 26684
rect 10892 26462 10894 26514
rect 10946 26462 10948 26514
rect 10892 26450 10948 26462
rect 10892 26290 10948 26302
rect 11116 26292 11172 26302
rect 10892 26238 10894 26290
rect 10946 26238 10948 26290
rect 10892 26068 10948 26238
rect 10892 26002 10948 26012
rect 11004 26290 11172 26292
rect 11004 26238 11118 26290
rect 11170 26238 11172 26290
rect 11004 26236 11172 26238
rect 10780 24670 10782 24722
rect 10834 24670 10836 24722
rect 10556 24556 10724 24612
rect 10444 23716 10500 23726
rect 10444 23622 10500 23660
rect 10556 23714 10612 23726
rect 10556 23662 10558 23714
rect 10610 23662 10612 23714
rect 10556 23604 10612 23662
rect 10556 23538 10612 23548
rect 10668 23266 10724 24556
rect 10668 23214 10670 23266
rect 10722 23214 10724 23266
rect 10668 23202 10724 23214
rect 10444 23156 10500 23166
rect 10444 23154 10612 23156
rect 10444 23102 10446 23154
rect 10498 23102 10612 23154
rect 10444 23100 10612 23102
rect 10444 23090 10500 23100
rect 10332 21924 10388 22316
rect 10444 22148 10500 22158
rect 10444 22054 10500 22092
rect 10556 22036 10612 23100
rect 10780 23044 10836 24670
rect 10668 22988 10836 23044
rect 10892 24724 10948 24734
rect 10668 22258 10724 22988
rect 10780 22820 10836 22830
rect 10780 22594 10836 22764
rect 10780 22542 10782 22594
rect 10834 22542 10836 22594
rect 10780 22530 10836 22542
rect 10668 22206 10670 22258
rect 10722 22206 10724 22258
rect 10668 22194 10724 22206
rect 10556 21980 10724 22036
rect 10332 21868 10612 21924
rect 10556 21810 10612 21868
rect 10556 21758 10558 21810
rect 10610 21758 10612 21810
rect 10556 21746 10612 21758
rect 10108 21698 10276 21700
rect 10108 21646 10110 21698
rect 10162 21646 10276 21698
rect 10108 21644 10276 21646
rect 10108 21634 10164 21644
rect 10332 21588 10388 21598
rect 9996 21410 10052 21420
rect 10220 21586 10388 21588
rect 10220 21534 10334 21586
rect 10386 21534 10388 21586
rect 10220 21532 10388 21534
rect 10220 20132 10276 21532
rect 10332 21522 10388 21532
rect 10556 21474 10612 21486
rect 10556 21422 10558 21474
rect 10610 21422 10612 21474
rect 10332 21028 10388 21038
rect 10332 20802 10388 20972
rect 10332 20750 10334 20802
rect 10386 20750 10388 20802
rect 10332 20738 10388 20750
rect 10556 20804 10612 21422
rect 10556 20738 10612 20748
rect 9996 20076 10276 20132
rect 10668 20130 10724 21980
rect 10668 20078 10670 20130
rect 10722 20078 10724 20130
rect 9996 18788 10052 20076
rect 10668 20066 10724 20078
rect 10780 21924 10836 21934
rect 10444 20020 10500 20030
rect 10500 19964 10612 20020
rect 10444 19926 10500 19964
rect 10332 19906 10388 19918
rect 10332 19854 10334 19906
rect 10386 19854 10388 19906
rect 10332 19684 10388 19854
rect 10332 19618 10388 19628
rect 9996 18722 10052 18732
rect 10108 19572 10164 19582
rect 9772 18398 9774 18450
rect 9826 18398 9828 18450
rect 9772 18340 9828 18398
rect 9212 17838 9214 17890
rect 9266 17838 9268 17890
rect 9212 17826 9268 17838
rect 9772 17892 9828 18284
rect 10108 17892 10164 19516
rect 10332 19348 10388 19358
rect 10332 19254 10388 19292
rect 10220 19234 10276 19246
rect 10220 19182 10222 19234
rect 10274 19182 10276 19234
rect 10220 19124 10276 19182
rect 10220 19058 10276 19068
rect 10444 19236 10500 19246
rect 10220 18788 10276 18798
rect 10220 18116 10276 18732
rect 10332 18340 10388 18350
rect 10444 18340 10500 19180
rect 10332 18338 10500 18340
rect 10332 18286 10334 18338
rect 10386 18286 10500 18338
rect 10332 18284 10500 18286
rect 10556 18564 10612 19964
rect 10780 19572 10836 21868
rect 10892 19908 10948 24668
rect 10892 19842 10948 19852
rect 10780 19506 10836 19516
rect 10892 19236 10948 19246
rect 10892 19142 10948 19180
rect 10332 18274 10388 18284
rect 10220 18060 10388 18116
rect 10220 17892 10276 17902
rect 10108 17890 10276 17892
rect 10108 17838 10222 17890
rect 10274 17838 10276 17890
rect 10108 17836 10276 17838
rect 9772 17826 9828 17836
rect 10220 17826 10276 17836
rect 9324 17780 9380 17790
rect 9324 17668 9380 17724
rect 9660 17780 9716 17790
rect 9660 17686 9716 17724
rect 9100 17054 9102 17106
rect 9154 17054 9156 17106
rect 9100 17042 9156 17054
rect 9212 17612 9380 17668
rect 9884 17666 9940 17678
rect 9884 17614 9886 17666
rect 9938 17614 9940 17666
rect 8652 16882 8932 16884
rect 8652 16830 8654 16882
rect 8706 16830 8932 16882
rect 8652 16828 8932 16830
rect 8652 16818 8708 16828
rect 8764 16548 8820 16558
rect 8652 15540 8708 15550
rect 8652 15446 8708 15484
rect 8316 13458 8372 13468
rect 8428 15092 8596 15148
rect 8428 12180 8484 15092
rect 8652 14532 8708 14542
rect 8652 14438 8708 14476
rect 8428 12114 8484 12124
rect 8540 14420 8596 14430
rect 8540 13746 8596 14364
rect 8764 14308 8820 16492
rect 9100 16212 9156 16222
rect 8876 15874 8932 15886
rect 8876 15822 8878 15874
rect 8930 15822 8932 15874
rect 8876 15764 8932 15822
rect 8876 15698 8932 15708
rect 8988 15876 9044 15886
rect 8540 13694 8542 13746
rect 8594 13694 8596 13746
rect 8204 11732 8372 11788
rect 8316 11506 8372 11732
rect 8316 11454 8318 11506
rect 8370 11454 8372 11506
rect 8316 11442 8372 11454
rect 7980 11004 8092 11060
rect 7868 10724 7924 10734
rect 7868 10630 7924 10668
rect 7756 10612 7812 10622
rect 7756 10518 7812 10556
rect 7756 8932 7812 8942
rect 7644 8876 7756 8932
rect 7756 8838 7812 8876
rect 7420 8148 7476 8158
rect 7308 8146 7476 8148
rect 7308 8094 7422 8146
rect 7474 8094 7476 8146
rect 7308 8092 7476 8094
rect 7420 8082 7476 8092
rect 7420 7924 7476 7934
rect 7308 7700 7364 7710
rect 7308 7606 7364 7644
rect 7308 6132 7364 6142
rect 7420 6132 7476 7868
rect 7532 7586 7588 8204
rect 7532 7534 7534 7586
rect 7586 7534 7588 7586
rect 7532 7522 7588 7534
rect 7644 8258 7700 8270
rect 7644 8206 7646 8258
rect 7698 8206 7700 8258
rect 7644 6804 7700 8206
rect 7980 8036 8036 11004
rect 8092 10994 8148 11004
rect 8316 10724 8372 10734
rect 8204 10612 8260 10622
rect 8092 9940 8148 9950
rect 8092 9846 8148 9884
rect 8204 9492 8260 10556
rect 7868 7980 8036 8036
rect 8092 9436 8260 9492
rect 7756 7700 7812 7710
rect 7756 7586 7812 7644
rect 7756 7534 7758 7586
rect 7810 7534 7812 7586
rect 7756 7522 7812 7534
rect 7644 6738 7700 6748
rect 7868 6692 7924 7980
rect 7308 6130 7476 6132
rect 7308 6078 7310 6130
rect 7362 6078 7476 6130
rect 7308 6076 7476 6078
rect 7756 6636 7924 6692
rect 7980 7812 8036 7822
rect 7308 6066 7364 6076
rect 7644 5796 7700 5806
rect 7644 5702 7700 5740
rect 7308 5348 7364 5358
rect 7308 5234 7364 5292
rect 7308 5182 7310 5234
rect 7362 5182 7364 5234
rect 7308 5170 7364 5182
rect 7756 5012 7812 6636
rect 7868 6466 7924 6478
rect 7868 6414 7870 6466
rect 7922 6414 7924 6466
rect 7868 5796 7924 6414
rect 7868 5730 7924 5740
rect 7308 4956 7812 5012
rect 7868 5122 7924 5134
rect 7868 5070 7870 5122
rect 7922 5070 7924 5122
rect 7868 5012 7924 5070
rect 7308 4562 7364 4956
rect 7868 4946 7924 4956
rect 7308 4510 7310 4562
rect 7362 4510 7364 4562
rect 7308 4498 7364 4510
rect 7196 4162 7252 4172
rect 7756 4226 7812 4238
rect 7756 4174 7758 4226
rect 7810 4174 7812 4226
rect 7756 4114 7812 4174
rect 7756 4062 7758 4114
rect 7810 4062 7812 4114
rect 7756 4050 7812 4062
rect 7196 3666 7252 3678
rect 7196 3614 7198 3666
rect 7250 3614 7252 3666
rect 7196 2324 7252 3614
rect 7756 3668 7812 3678
rect 7980 3668 8036 7756
rect 8092 6580 8148 9436
rect 8204 9268 8260 9278
rect 8204 9174 8260 9212
rect 8316 8708 8372 10668
rect 8540 9940 8596 13694
rect 8652 14252 8820 14308
rect 8988 15204 9044 15820
rect 9100 15764 9156 16156
rect 9100 15698 9156 15708
rect 8652 12402 8708 14252
rect 8876 13860 8932 13870
rect 8876 13766 8932 13804
rect 8764 13524 8820 13534
rect 8764 12850 8820 13468
rect 8764 12798 8766 12850
rect 8818 12798 8820 12850
rect 8764 12786 8820 12798
rect 8652 12350 8654 12402
rect 8706 12350 8708 12402
rect 8652 12338 8708 12350
rect 8988 12404 9044 15148
rect 9100 14530 9156 14542
rect 9100 14478 9102 14530
rect 9154 14478 9156 14530
rect 9100 13188 9156 14478
rect 9212 13636 9268 17612
rect 9884 17332 9940 17614
rect 10332 17444 10388 18060
rect 10556 17892 10612 18508
rect 10780 19012 10836 19022
rect 10780 18450 10836 18956
rect 10780 18398 10782 18450
rect 10834 18398 10836 18450
rect 10780 18228 10836 18398
rect 10836 18172 10948 18228
rect 10780 18162 10836 18172
rect 10556 17836 10836 17892
rect 10780 17666 10836 17836
rect 10780 17614 10782 17666
rect 10834 17614 10836 17666
rect 10780 17602 10836 17614
rect 10332 17378 10388 17388
rect 9884 17266 9940 17276
rect 10108 17108 10164 17118
rect 10108 17014 10164 17052
rect 10332 17108 10388 17118
rect 9772 16882 9828 16894
rect 9772 16830 9774 16882
rect 9826 16830 9828 16882
rect 9772 16772 9828 16830
rect 9324 16436 9380 16446
rect 9324 15986 9380 16380
rect 9660 16324 9716 16334
rect 9324 15934 9326 15986
rect 9378 15934 9380 15986
rect 9324 15922 9380 15934
rect 9548 16098 9604 16110
rect 9548 16046 9550 16098
rect 9602 16046 9604 16098
rect 9548 15148 9604 16046
rect 9660 15538 9716 16268
rect 9660 15486 9662 15538
rect 9714 15486 9716 15538
rect 9660 15474 9716 15486
rect 9436 15092 9604 15148
rect 9772 15148 9828 16716
rect 10332 16210 10388 17052
rect 10892 17108 10948 18172
rect 11004 17666 11060 26236
rect 11116 26226 11172 26236
rect 11228 25282 11284 25294
rect 11228 25230 11230 25282
rect 11282 25230 11284 25282
rect 11228 25172 11284 25230
rect 11228 25106 11284 25116
rect 11340 23378 11396 28364
rect 11452 28196 11508 28206
rect 11452 27970 11508 28140
rect 11452 27918 11454 27970
rect 11506 27918 11508 27970
rect 11452 26962 11508 27918
rect 11676 27858 11732 28476
rect 11676 27806 11678 27858
rect 11730 27806 11732 27858
rect 11676 27300 11732 27806
rect 11676 27234 11732 27244
rect 11452 26910 11454 26962
rect 11506 26910 11508 26962
rect 11452 26740 11508 26910
rect 11452 25732 11508 26684
rect 11788 26180 11844 26190
rect 11788 26086 11844 26124
rect 11452 25666 11508 25676
rect 11564 25956 11620 25966
rect 11452 25508 11508 25518
rect 11452 25414 11508 25452
rect 11564 25506 11620 25900
rect 11564 25454 11566 25506
rect 11618 25454 11620 25506
rect 11564 25442 11620 25454
rect 11676 25284 11732 25294
rect 11676 25282 11844 25284
rect 11676 25230 11678 25282
rect 11730 25230 11844 25282
rect 11676 25228 11844 25230
rect 11676 25218 11732 25228
rect 11452 24948 11508 24958
rect 11452 24164 11508 24892
rect 11564 24612 11620 24622
rect 11564 24610 11732 24612
rect 11564 24558 11566 24610
rect 11618 24558 11732 24610
rect 11564 24556 11732 24558
rect 11564 24546 11620 24556
rect 11564 24164 11620 24174
rect 11452 24162 11620 24164
rect 11452 24110 11566 24162
rect 11618 24110 11620 24162
rect 11452 24108 11620 24110
rect 11564 23940 11620 24108
rect 11564 23874 11620 23884
rect 11340 23326 11342 23378
rect 11394 23326 11396 23378
rect 11340 23314 11396 23326
rect 11116 22372 11172 22382
rect 11116 22036 11172 22316
rect 11116 21586 11172 21980
rect 11116 21534 11118 21586
rect 11170 21534 11172 21586
rect 11116 21522 11172 21534
rect 11228 22148 11284 22158
rect 11004 17614 11006 17666
rect 11058 17614 11060 17666
rect 11004 17602 11060 17614
rect 11116 19684 11172 19694
rect 11116 17666 11172 19628
rect 11116 17614 11118 17666
rect 11170 17614 11172 17666
rect 11116 17602 11172 17614
rect 10892 17042 10948 17052
rect 11004 17444 11060 17454
rect 11004 17106 11060 17388
rect 11004 17054 11006 17106
rect 11058 17054 11060 17106
rect 11004 16996 11060 17054
rect 11004 16930 11060 16940
rect 10332 16158 10334 16210
rect 10386 16158 10388 16210
rect 10332 16146 10388 16158
rect 10668 16882 10724 16894
rect 10668 16830 10670 16882
rect 10722 16830 10724 16882
rect 10556 16100 10612 16110
rect 10556 15652 10612 16044
rect 10668 15988 10724 16830
rect 11116 16100 11172 16110
rect 10668 15922 10724 15932
rect 10780 16098 11172 16100
rect 10780 16046 11118 16098
rect 11170 16046 11172 16098
rect 10780 16044 11172 16046
rect 9884 15428 9940 15438
rect 9884 15334 9940 15372
rect 10556 15426 10612 15596
rect 10556 15374 10558 15426
rect 10610 15374 10612 15426
rect 10556 15362 10612 15374
rect 10780 15428 10836 16044
rect 11116 16034 11172 16044
rect 10892 15874 10948 15886
rect 10892 15822 10894 15874
rect 10946 15822 10948 15874
rect 10892 15540 10948 15822
rect 11004 15876 11060 15886
rect 11228 15876 11284 22092
rect 11676 21812 11732 24556
rect 11788 24164 11844 25228
rect 11788 24032 11844 24108
rect 11788 23716 11844 23726
rect 11788 23154 11844 23660
rect 11788 23102 11790 23154
rect 11842 23102 11844 23154
rect 11788 23090 11844 23102
rect 11788 22932 11844 22942
rect 11788 22482 11844 22876
rect 11788 22430 11790 22482
rect 11842 22430 11844 22482
rect 11788 22418 11844 22430
rect 11452 21756 11732 21812
rect 11340 19684 11396 19694
rect 11452 19684 11508 21756
rect 11564 20578 11620 20590
rect 11564 20526 11566 20578
rect 11618 20526 11620 20578
rect 11564 20468 11620 20526
rect 11564 20402 11620 20412
rect 11676 20356 11732 20366
rect 11676 20132 11732 20300
rect 11676 20076 11788 20132
rect 11732 20030 11788 20076
rect 11732 20018 11844 20030
rect 11732 19966 11790 20018
rect 11842 19966 11844 20018
rect 11732 19964 11844 19966
rect 11788 19954 11844 19964
rect 11396 19628 11508 19684
rect 11340 19010 11396 19628
rect 11340 18958 11342 19010
rect 11394 18958 11396 19010
rect 11340 18452 11396 18958
rect 11788 19012 11844 19022
rect 11788 18918 11844 18956
rect 11788 18676 11844 18686
rect 11340 18386 11396 18396
rect 11564 18564 11620 18574
rect 11452 18340 11508 18350
rect 11452 18246 11508 18284
rect 11452 18004 11508 18014
rect 11340 17442 11396 17454
rect 11340 17390 11342 17442
rect 11394 17390 11396 17442
rect 11340 16100 11396 17390
rect 11340 16034 11396 16044
rect 11004 15874 11284 15876
rect 11004 15822 11006 15874
rect 11058 15822 11284 15874
rect 11004 15820 11284 15822
rect 11340 15874 11396 15886
rect 11340 15822 11342 15874
rect 11394 15822 11396 15874
rect 11004 15810 11060 15820
rect 10892 15484 11060 15540
rect 9996 15314 10052 15326
rect 9996 15262 9998 15314
rect 10050 15262 10052 15314
rect 9772 15092 9940 15148
rect 9324 14532 9380 14542
rect 9436 14532 9492 15092
rect 9548 14756 9604 14766
rect 9548 14662 9604 14700
rect 9324 14530 9492 14532
rect 9324 14478 9326 14530
rect 9378 14478 9492 14530
rect 9324 14476 9492 14478
rect 9324 14466 9380 14476
rect 9212 13570 9268 13580
rect 9100 13132 9380 13188
rect 9100 12964 9156 12974
rect 9100 12870 9156 12908
rect 8988 12348 9268 12404
rect 8988 12178 9044 12190
rect 8988 12126 8990 12178
rect 9042 12126 9044 12178
rect 8988 11844 9044 12126
rect 8988 11778 9044 11788
rect 8876 11620 8932 11630
rect 8876 11394 8932 11564
rect 8876 11342 8878 11394
rect 8930 11342 8932 11394
rect 8876 11330 8932 11342
rect 8876 11060 8932 11070
rect 8876 10722 8932 11004
rect 8876 10670 8878 10722
rect 8930 10670 8932 10722
rect 8876 10658 8932 10670
rect 8540 9884 8708 9940
rect 8540 9716 8596 9726
rect 8092 6514 8148 6524
rect 8204 8652 8372 8708
rect 8428 9714 8596 9716
rect 8428 9662 8542 9714
rect 8594 9662 8596 9714
rect 8428 9660 8596 9662
rect 8204 8036 8260 8652
rect 8428 8428 8484 9660
rect 8540 9650 8596 9660
rect 8540 8932 8596 8942
rect 8540 8838 8596 8876
rect 8652 8708 8708 9884
rect 8092 6244 8148 6254
rect 8092 4226 8148 6188
rect 8204 6020 8260 7980
rect 8316 8372 8484 8428
rect 8540 8652 8708 8708
rect 8876 9938 8932 9950
rect 8876 9886 8878 9938
rect 8930 9886 8932 9938
rect 8876 8932 8932 9886
rect 8316 7812 8372 8372
rect 8316 7746 8372 7756
rect 8428 8260 8484 8270
rect 8428 6802 8484 8204
rect 8428 6750 8430 6802
rect 8482 6750 8484 6802
rect 8428 6738 8484 6750
rect 8540 7812 8596 8652
rect 8764 8260 8820 8270
rect 8764 8166 8820 8204
rect 8540 6132 8596 7756
rect 8652 7586 8708 7598
rect 8652 7534 8654 7586
rect 8706 7534 8708 7586
rect 8652 7364 8708 7534
rect 8652 7298 8708 7308
rect 8540 6130 8820 6132
rect 8540 6078 8542 6130
rect 8594 6078 8820 6130
rect 8540 6076 8820 6078
rect 8540 6066 8596 6076
rect 8204 5964 8372 6020
rect 8204 5794 8260 5806
rect 8204 5742 8206 5794
rect 8258 5742 8260 5794
rect 8204 5684 8260 5742
rect 8204 5618 8260 5628
rect 8316 5460 8372 5964
rect 8204 5404 8372 5460
rect 8428 5796 8484 5806
rect 8204 5234 8260 5404
rect 8428 5348 8484 5740
rect 8204 5182 8206 5234
rect 8258 5182 8260 5234
rect 8204 5170 8260 5182
rect 8316 5292 8484 5348
rect 8092 4174 8094 4226
rect 8146 4174 8148 4226
rect 8092 4114 8148 4174
rect 8092 4062 8094 4114
rect 8146 4062 8148 4114
rect 8092 4050 8148 4062
rect 8204 4340 8260 4350
rect 7756 3666 8036 3668
rect 7756 3614 7758 3666
rect 7810 3614 8036 3666
rect 7756 3612 8036 3614
rect 8204 3666 8260 4284
rect 8204 3614 8206 3666
rect 8258 3614 8260 3666
rect 7756 3602 7812 3612
rect 8204 3602 8260 3614
rect 7196 2258 7252 2268
rect 6188 1474 6244 1484
rect 8316 1428 8372 5292
rect 8764 5234 8820 6076
rect 8764 5182 8766 5234
rect 8818 5182 8820 5234
rect 8764 5124 8820 5182
rect 8764 5058 8820 5068
rect 8652 4564 8708 4574
rect 8652 4470 8708 4508
rect 8652 3668 8708 3678
rect 8876 3668 8932 8876
rect 8988 9826 9044 9838
rect 8988 9774 8990 9826
rect 9042 9774 9044 9826
rect 8988 8372 9044 9774
rect 9100 9268 9156 9278
rect 9212 9268 9268 12348
rect 9324 11732 9380 13132
rect 9324 11666 9380 11676
rect 9100 9266 9268 9268
rect 9100 9214 9102 9266
rect 9154 9214 9268 9266
rect 9100 9212 9268 9214
rect 9100 9202 9156 9212
rect 8988 8306 9044 8316
rect 9100 8820 9156 8830
rect 8988 8148 9044 8158
rect 8988 7698 9044 8092
rect 8988 7646 8990 7698
rect 9042 7646 9044 7698
rect 8988 7634 9044 7646
rect 8988 6468 9044 6478
rect 8988 6374 9044 6412
rect 9100 5794 9156 8764
rect 9436 8820 9492 14476
rect 9772 14420 9828 14430
rect 9772 14326 9828 14364
rect 9772 13860 9828 13870
rect 9884 13860 9940 15092
rect 9828 13804 9940 13860
rect 9772 13766 9828 13804
rect 9660 12964 9716 12974
rect 9660 12290 9716 12908
rect 9996 12516 10052 15262
rect 10332 14530 10388 14542
rect 10332 14478 10334 14530
rect 10386 14478 10388 14530
rect 10332 14308 10388 14478
rect 10444 14532 10500 14542
rect 10444 14418 10500 14476
rect 10444 14366 10446 14418
rect 10498 14366 10500 14418
rect 10444 14354 10500 14366
rect 10668 14532 10724 14542
rect 10332 14242 10388 14252
rect 10332 13524 10388 13534
rect 10332 13430 10388 13468
rect 10108 13076 10164 13086
rect 10108 12982 10164 13020
rect 9660 12238 9662 12290
rect 9714 12238 9716 12290
rect 9660 12226 9716 12238
rect 9772 12460 10052 12516
rect 9772 10052 9828 12460
rect 10220 12404 10276 12414
rect 9884 12180 9940 12190
rect 9884 12086 9940 12124
rect 10108 11284 10164 11294
rect 10108 10610 10164 11228
rect 10108 10558 10110 10610
rect 10162 10558 10164 10610
rect 10108 10388 10164 10558
rect 10108 10322 10164 10332
rect 10220 10164 10276 12348
rect 10668 12404 10724 14476
rect 10668 12338 10724 12348
rect 10780 14420 10836 15372
rect 11004 14868 11060 15484
rect 11004 14802 11060 14812
rect 11116 15202 11172 15214
rect 11116 15150 11118 15202
rect 11170 15150 11172 15202
rect 10556 12292 10612 12302
rect 10444 12178 10500 12190
rect 10444 12126 10446 12178
rect 10498 12126 10500 12178
rect 10444 11844 10500 12126
rect 10444 11778 10500 11788
rect 10444 11396 10500 11406
rect 10444 11302 10500 11340
rect 9772 9986 9828 9996
rect 10108 10108 10276 10164
rect 10444 10500 10500 10510
rect 10556 10500 10612 12236
rect 10668 11508 10724 11518
rect 10668 11394 10724 11452
rect 10668 11342 10670 11394
rect 10722 11342 10724 11394
rect 10668 11330 10724 11342
rect 10780 10948 10836 14364
rect 11004 14418 11060 14430
rect 11004 14366 11006 14418
rect 11058 14366 11060 14418
rect 11004 13748 11060 14366
rect 11116 14196 11172 15150
rect 11340 15092 11396 15822
rect 11452 15538 11508 17948
rect 11452 15486 11454 15538
rect 11506 15486 11508 15538
rect 11452 15474 11508 15486
rect 11340 15090 11508 15092
rect 11340 15038 11342 15090
rect 11394 15038 11508 15090
rect 11340 15036 11508 15038
rect 11340 15026 11396 15036
rect 11116 14130 11172 14140
rect 11452 14530 11508 15036
rect 11452 14478 11454 14530
rect 11506 14478 11508 14530
rect 11228 13748 11284 13758
rect 11004 13746 11284 13748
rect 11004 13694 11230 13746
rect 11282 13694 11284 13746
rect 11004 13692 11284 13694
rect 11228 13636 11284 13692
rect 11228 13570 11284 13580
rect 10444 10498 10612 10500
rect 10444 10446 10446 10498
rect 10498 10446 10612 10498
rect 10444 10444 10612 10446
rect 10668 10892 10836 10948
rect 10892 12852 10948 12862
rect 11452 12852 11508 14478
rect 11564 13524 11620 18508
rect 11788 18340 11844 18620
rect 11900 18564 11956 29708
rect 12012 28868 12068 30604
rect 12012 28802 12068 28812
rect 12124 30548 12180 30558
rect 12012 28082 12068 28094
rect 12012 28030 12014 28082
rect 12066 28030 12068 28082
rect 12012 27972 12068 28030
rect 12012 27906 12068 27916
rect 12124 24946 12180 30492
rect 12460 29986 12516 29998
rect 12460 29934 12462 29986
rect 12514 29934 12516 29986
rect 12236 29428 12292 29438
rect 12236 27860 12292 29372
rect 12236 27766 12292 27804
rect 12348 28420 12404 28430
rect 12236 27412 12292 27422
rect 12236 26964 12292 27356
rect 12348 27074 12404 28364
rect 12348 27022 12350 27074
rect 12402 27022 12404 27074
rect 12348 27010 12404 27022
rect 12236 26852 12404 26908
rect 12236 26180 12292 26190
rect 12236 26086 12292 26124
rect 12348 25620 12404 26852
rect 12460 26516 12516 29934
rect 12572 29092 12628 33964
rect 12796 33954 12852 33964
rect 12908 34690 12964 34702
rect 12908 34638 12910 34690
rect 12962 34638 12964 34690
rect 12908 33908 12964 34638
rect 13244 34020 13300 34748
rect 13244 33926 13300 33964
rect 12908 33842 12964 33852
rect 13356 33908 13412 36988
rect 13468 36484 13524 36494
rect 13468 34244 13524 36428
rect 13580 34692 13636 37212
rect 13916 36708 13972 36718
rect 13916 36594 13972 36652
rect 13916 36542 13918 36594
rect 13970 36542 13972 36594
rect 13916 36530 13972 36542
rect 14028 36260 14084 36270
rect 14028 35810 14084 36204
rect 14140 35922 14196 39566
rect 14364 39396 14420 40126
rect 14476 40180 14532 40190
rect 14476 39620 14532 40124
rect 14588 40068 14644 45052
rect 14700 44772 14756 45276
rect 16604 45556 16660 45566
rect 16268 45106 16324 45118
rect 16268 45054 16270 45106
rect 16322 45054 16324 45106
rect 15260 44996 15316 45006
rect 14700 44706 14756 44716
rect 15036 44994 15316 44996
rect 15036 44942 15262 44994
rect 15314 44942 15316 44994
rect 15036 44940 15316 44942
rect 14812 44324 14868 44334
rect 14812 44230 14868 44268
rect 15036 44322 15092 44940
rect 15260 44930 15316 44940
rect 15932 44994 15988 45006
rect 15932 44942 15934 44994
rect 15986 44942 15988 44994
rect 15036 44270 15038 44322
rect 15090 44270 15092 44322
rect 15036 43988 15092 44270
rect 15820 44322 15876 44334
rect 15820 44270 15822 44322
rect 15874 44270 15876 44322
rect 15036 43922 15092 43932
rect 15148 44210 15204 44222
rect 15148 44158 15150 44210
rect 15202 44158 15204 44210
rect 15036 43764 15092 43774
rect 15036 43538 15092 43708
rect 15036 43486 15038 43538
rect 15090 43486 15092 43538
rect 15036 43474 15092 43486
rect 15148 43540 15204 44158
rect 15596 44098 15652 44110
rect 15596 44046 15598 44098
rect 15650 44046 15652 44098
rect 15148 43474 15204 43484
rect 15484 43540 15540 43550
rect 15596 43540 15652 44046
rect 15820 43764 15876 44270
rect 15932 43988 15988 44942
rect 16044 44324 16100 44334
rect 16268 44324 16324 45054
rect 16604 44996 16660 45500
rect 16716 45218 16772 46734
rect 17612 46340 17668 49644
rect 19964 49700 20020 49710
rect 19964 49606 20020 49644
rect 20636 49700 20692 49758
rect 20636 49140 20692 49644
rect 21196 49698 21252 49710
rect 21196 49646 21198 49698
rect 21250 49646 21252 49698
rect 20860 49140 20916 49150
rect 20636 49138 20916 49140
rect 20636 49086 20862 49138
rect 20914 49086 20916 49138
rect 20636 49084 20916 49086
rect 20860 49028 20916 49084
rect 20860 48962 20916 48972
rect 18956 48916 19012 48926
rect 18956 48914 19684 48916
rect 18956 48862 18958 48914
rect 19010 48862 19684 48914
rect 18956 48860 19684 48862
rect 18956 48850 19012 48860
rect 18732 48802 18788 48814
rect 18732 48750 18734 48802
rect 18786 48750 18788 48802
rect 17724 48468 17780 48478
rect 17724 48374 17780 48412
rect 17948 48468 18004 48478
rect 17948 48244 18004 48412
rect 18732 48468 18788 48750
rect 18732 48402 18788 48412
rect 18844 48802 18900 48814
rect 18844 48750 18846 48802
rect 18898 48750 18900 48802
rect 17948 48178 18004 48188
rect 18172 48354 18228 48366
rect 18172 48302 18174 48354
rect 18226 48302 18228 48354
rect 17836 48130 17892 48142
rect 17836 48078 17838 48130
rect 17890 48078 17892 48130
rect 17836 46564 17892 48078
rect 17948 47236 18004 47246
rect 18172 47236 18228 48302
rect 18844 48242 18900 48750
rect 18956 48356 19012 48366
rect 18956 48262 19012 48300
rect 18844 48190 18846 48242
rect 18898 48190 18900 48242
rect 18844 48178 18900 48190
rect 19516 48130 19572 48142
rect 19516 48078 19518 48130
rect 19570 48078 19572 48130
rect 19404 48020 19460 48030
rect 18284 47572 18340 47582
rect 18284 47478 18340 47516
rect 19292 47458 19348 47470
rect 19292 47406 19294 47458
rect 19346 47406 19348 47458
rect 17948 47234 18116 47236
rect 17948 47182 17950 47234
rect 18002 47182 18116 47234
rect 17948 47180 18116 47182
rect 17948 47170 18004 47180
rect 18060 46900 18116 47180
rect 18172 47142 18228 47180
rect 18396 47234 18452 47246
rect 18396 47182 18398 47234
rect 18450 47182 18452 47234
rect 18284 46900 18340 46910
rect 18060 46898 18340 46900
rect 18060 46846 18286 46898
rect 18338 46846 18340 46898
rect 18060 46844 18340 46846
rect 18284 46834 18340 46844
rect 17836 46498 17892 46508
rect 18396 46340 18452 47182
rect 18956 47124 19012 47134
rect 17612 46284 18340 46340
rect 16716 45166 16718 45218
rect 16770 45166 16772 45218
rect 16716 45154 16772 45166
rect 16604 44940 16772 44996
rect 16492 44324 16548 44334
rect 16044 44322 16548 44324
rect 16044 44270 16046 44322
rect 16098 44270 16494 44322
rect 16546 44270 16548 44322
rect 16044 44268 16548 44270
rect 16044 44258 16100 44268
rect 16492 44258 16548 44268
rect 16268 44098 16324 44110
rect 16268 44046 16270 44098
rect 16322 44046 16324 44098
rect 16268 43988 16324 44046
rect 16380 44100 16436 44110
rect 16716 44100 16772 44940
rect 17724 44994 17780 45006
rect 18060 44996 18116 45006
rect 17724 44942 17726 44994
rect 17778 44942 17780 44994
rect 16380 44098 16772 44100
rect 16380 44046 16382 44098
rect 16434 44046 16772 44098
rect 16380 44044 16772 44046
rect 16940 44322 16996 44334
rect 16940 44270 16942 44322
rect 16994 44270 16996 44322
rect 16380 44034 16436 44044
rect 15932 43932 16324 43988
rect 15932 43764 15988 43774
rect 15820 43762 15988 43764
rect 15820 43710 15934 43762
rect 15986 43710 15988 43762
rect 15820 43708 15988 43710
rect 16268 43708 16324 43932
rect 15932 43698 15988 43708
rect 16156 43652 16324 43708
rect 16604 43876 16660 43886
rect 15484 43538 15652 43540
rect 15484 43486 15486 43538
rect 15538 43486 15652 43538
rect 15484 43484 15652 43486
rect 15820 43540 15876 43550
rect 15484 43474 15540 43484
rect 15260 43314 15316 43326
rect 15260 43262 15262 43314
rect 15314 43262 15316 43314
rect 15260 42868 15316 43262
rect 15372 42868 15428 42878
rect 15260 42866 15428 42868
rect 15260 42814 15374 42866
rect 15426 42814 15428 42866
rect 15260 42812 15428 42814
rect 15372 42802 15428 42812
rect 15820 42754 15876 43484
rect 15820 42702 15822 42754
rect 15874 42702 15876 42754
rect 15260 42642 15316 42654
rect 15260 42590 15262 42642
rect 15314 42590 15316 42642
rect 14700 42530 14756 42542
rect 14700 42478 14702 42530
rect 14754 42478 14756 42530
rect 14700 42420 14756 42478
rect 15260 42532 15316 42590
rect 15260 42466 15316 42476
rect 15596 42642 15652 42654
rect 15596 42590 15598 42642
rect 15650 42590 15652 42642
rect 14700 42354 14756 42364
rect 15596 42420 15652 42590
rect 15596 42354 15652 42364
rect 15708 42196 15764 42206
rect 15820 42196 15876 42702
rect 15708 42194 15876 42196
rect 15708 42142 15710 42194
rect 15762 42142 15876 42194
rect 15708 42140 15876 42142
rect 15708 42130 15764 42140
rect 14924 42084 14980 42094
rect 14924 41858 14980 42028
rect 14924 41806 14926 41858
rect 14978 41806 14980 41858
rect 14588 40002 14644 40012
rect 14700 40964 14756 40974
rect 14476 39618 14644 39620
rect 14476 39566 14478 39618
rect 14530 39566 14644 39618
rect 14476 39564 14644 39566
rect 14476 39554 14532 39564
rect 14364 39330 14420 39340
rect 14476 39284 14532 39294
rect 14476 39058 14532 39228
rect 14476 39006 14478 39058
rect 14530 39006 14532 39058
rect 14476 38994 14532 39006
rect 14252 38836 14308 38846
rect 14252 38834 14420 38836
rect 14252 38782 14254 38834
rect 14306 38782 14420 38834
rect 14252 38780 14420 38782
rect 14252 38770 14308 38780
rect 14364 37492 14420 38780
rect 14364 37266 14420 37436
rect 14364 37214 14366 37266
rect 14418 37214 14420 37266
rect 14364 37202 14420 37214
rect 14476 38162 14532 38174
rect 14476 38110 14478 38162
rect 14530 38110 14532 38162
rect 14252 37156 14308 37166
rect 14252 37062 14308 37100
rect 14476 37044 14532 38110
rect 14588 38162 14644 39564
rect 14588 38110 14590 38162
rect 14642 38110 14644 38162
rect 14588 38098 14644 38110
rect 14588 37380 14644 37390
rect 14588 37286 14644 37324
rect 14140 35870 14142 35922
rect 14194 35870 14196 35922
rect 14140 35858 14196 35870
rect 14364 36370 14420 36382
rect 14364 36318 14366 36370
rect 14418 36318 14420 36370
rect 14028 35758 14030 35810
rect 14082 35758 14084 35810
rect 13692 34916 13748 34926
rect 13692 34822 13748 34860
rect 13804 34804 13860 34814
rect 13804 34710 13860 34748
rect 13580 34626 13636 34636
rect 13804 34244 13860 34254
rect 14028 34244 14084 35758
rect 14252 35700 14308 35710
rect 14364 35700 14420 36318
rect 14252 35698 14420 35700
rect 14252 35646 14254 35698
rect 14306 35646 14420 35698
rect 14252 35644 14420 35646
rect 14252 35588 14308 35644
rect 14252 35522 14308 35532
rect 14364 35028 14420 35038
rect 14476 35028 14532 36988
rect 14700 36708 14756 40908
rect 14924 39172 14980 41806
rect 15708 41972 15764 41982
rect 15148 40964 15204 40974
rect 15148 40870 15204 40908
rect 15148 40404 15204 40414
rect 15372 40404 15428 40414
rect 14924 39106 14980 39116
rect 15036 39394 15092 39406
rect 15036 39342 15038 39394
rect 15090 39342 15092 39394
rect 14924 38948 14980 38958
rect 14924 38834 14980 38892
rect 14924 38782 14926 38834
rect 14978 38782 14980 38834
rect 14924 38770 14980 38782
rect 14812 38612 14868 38622
rect 14812 38518 14868 38556
rect 15036 38500 15092 39342
rect 15148 38612 15204 40348
rect 15148 38546 15204 38556
rect 15260 40402 15428 40404
rect 15260 40350 15374 40402
rect 15426 40350 15428 40402
rect 15260 40348 15428 40350
rect 14812 38050 14868 38062
rect 14812 37998 14814 38050
rect 14866 37998 14868 38050
rect 14812 37492 14868 37998
rect 15036 37938 15092 38444
rect 15036 37886 15038 37938
rect 15090 37886 15092 37938
rect 15036 37874 15092 37886
rect 15148 38388 15204 38398
rect 14812 37426 14868 37436
rect 14924 37268 14980 37278
rect 14924 37174 14980 37212
rect 15148 37268 15204 38332
rect 15260 37940 15316 40348
rect 15372 40338 15428 40348
rect 15596 39396 15652 39406
rect 15260 37716 15316 37884
rect 15260 37650 15316 37660
rect 15372 39394 15652 39396
rect 15372 39342 15598 39394
rect 15650 39342 15652 39394
rect 15372 39340 15652 39342
rect 15148 37202 15204 37212
rect 15260 36932 15316 36942
rect 15148 36708 15204 36718
rect 14700 36652 14980 36708
rect 14588 36596 14644 36606
rect 14588 36370 14644 36540
rect 14812 36484 14868 36494
rect 14588 36318 14590 36370
rect 14642 36318 14644 36370
rect 14588 36260 14644 36318
rect 14588 36194 14644 36204
rect 14700 36372 14756 36382
rect 14700 36258 14756 36316
rect 14700 36206 14702 36258
rect 14754 36206 14756 36258
rect 14700 36194 14756 36206
rect 14812 35698 14868 36428
rect 14812 35646 14814 35698
rect 14866 35646 14868 35698
rect 14812 35634 14868 35646
rect 14364 35026 14532 35028
rect 14364 34974 14366 35026
rect 14418 34974 14532 35026
rect 14364 34972 14532 34974
rect 14364 34962 14420 34972
rect 14812 34916 14868 34926
rect 14700 34860 14812 34916
rect 14588 34356 14644 34366
rect 14700 34356 14756 34860
rect 14812 34822 14868 34860
rect 13468 34242 13860 34244
rect 13468 34190 13806 34242
rect 13858 34190 13860 34242
rect 13468 34188 13860 34190
rect 13804 34178 13860 34188
rect 13916 34188 14084 34244
rect 14140 34354 14756 34356
rect 14140 34302 14590 34354
rect 14642 34302 14756 34354
rect 14140 34300 14756 34302
rect 14140 34242 14196 34300
rect 14588 34290 14644 34300
rect 14140 34190 14142 34242
rect 14194 34190 14196 34242
rect 13356 33842 13412 33852
rect 13580 33236 13636 33246
rect 12908 33124 12964 33134
rect 12908 33030 12964 33068
rect 13580 32786 13636 33180
rect 13580 32734 13582 32786
rect 13634 32734 13636 32786
rect 13580 32722 13636 32734
rect 13692 33124 13748 33134
rect 13356 32562 13412 32574
rect 13356 32510 13358 32562
rect 13410 32510 13412 32562
rect 12684 32452 12740 32462
rect 12684 32358 12740 32396
rect 12796 31892 12852 31902
rect 12684 31108 12740 31118
rect 12684 31014 12740 31052
rect 12684 29988 12740 29998
rect 12684 29316 12740 29932
rect 12796 29986 12852 31836
rect 13356 31892 13412 32510
rect 13468 32564 13524 32574
rect 13468 32470 13524 32508
rect 13692 32564 13748 33068
rect 13692 32498 13748 32508
rect 13916 32228 13972 34188
rect 14140 34178 14196 34190
rect 14252 33908 14308 33918
rect 14028 33122 14084 33134
rect 14028 33070 14030 33122
rect 14082 33070 14084 33122
rect 14028 32676 14084 33070
rect 14028 32562 14084 32620
rect 14028 32510 14030 32562
rect 14082 32510 14084 32562
rect 14028 32498 14084 32510
rect 13356 31826 13412 31836
rect 13580 32172 13972 32228
rect 14140 32452 14196 32462
rect 13020 31556 13076 31566
rect 13020 31554 13300 31556
rect 13020 31502 13022 31554
rect 13074 31502 13300 31554
rect 13020 31500 13300 31502
rect 13020 31490 13076 31500
rect 13132 31220 13188 31230
rect 12796 29934 12798 29986
rect 12850 29934 12852 29986
rect 12796 29922 12852 29934
rect 12908 31218 13188 31220
rect 12908 31166 13134 31218
rect 13186 31166 13188 31218
rect 12908 31164 13188 31166
rect 12908 29986 12964 31164
rect 13132 31154 13188 31164
rect 12908 29934 12910 29986
rect 12962 29934 12964 29986
rect 12908 29764 12964 29934
rect 12908 29698 12964 29708
rect 13020 30996 13076 31006
rect 12684 29250 12740 29260
rect 12908 29316 12964 29326
rect 12572 29036 12740 29092
rect 12572 28868 12628 28878
rect 12572 27074 12628 28812
rect 12572 27022 12574 27074
rect 12626 27022 12628 27074
rect 12572 27010 12628 27022
rect 12460 26450 12516 26460
rect 12572 25620 12628 25630
rect 12348 25618 12628 25620
rect 12348 25566 12574 25618
rect 12626 25566 12628 25618
rect 12348 25564 12628 25566
rect 12572 25554 12628 25564
rect 12124 24894 12126 24946
rect 12178 24894 12180 24946
rect 12124 24882 12180 24894
rect 12012 24724 12068 24734
rect 12348 24724 12404 24734
rect 12012 24722 12180 24724
rect 12012 24670 12014 24722
rect 12066 24670 12180 24722
rect 12012 24668 12180 24670
rect 12012 24658 12068 24668
rect 12012 24276 12068 24286
rect 12012 24050 12068 24220
rect 12012 23998 12014 24050
rect 12066 23998 12068 24050
rect 12012 23986 12068 23998
rect 12124 23716 12180 24668
rect 12348 24722 12628 24724
rect 12348 24670 12350 24722
rect 12402 24670 12628 24722
rect 12348 24668 12628 24670
rect 12348 24658 12404 24668
rect 12460 24498 12516 24510
rect 12460 24446 12462 24498
rect 12514 24446 12516 24498
rect 12348 24052 12404 24062
rect 12460 24052 12516 24446
rect 12348 24050 12516 24052
rect 12348 23998 12350 24050
rect 12402 23998 12516 24050
rect 12348 23996 12516 23998
rect 12348 23986 12404 23996
rect 12236 23716 12292 23726
rect 12460 23716 12516 23726
rect 12572 23716 12628 24668
rect 12124 23714 12292 23716
rect 12124 23662 12238 23714
rect 12290 23662 12292 23714
rect 12124 23660 12292 23662
rect 12236 22820 12292 23660
rect 12236 22754 12292 22764
rect 12348 23714 12628 23716
rect 12348 23662 12462 23714
rect 12514 23662 12628 23714
rect 12348 23660 12628 23662
rect 12012 21756 12292 21812
rect 12012 18676 12068 21756
rect 12236 21698 12292 21756
rect 12236 21646 12238 21698
rect 12290 21646 12292 21698
rect 12236 21634 12292 21646
rect 12124 21588 12180 21598
rect 12124 21494 12180 21532
rect 12348 21364 12404 23660
rect 12460 23650 12516 23660
rect 12684 23492 12740 29036
rect 12908 28754 12964 29260
rect 12908 28702 12910 28754
rect 12962 28702 12964 28754
rect 12908 28690 12964 28702
rect 13020 28082 13076 30940
rect 13244 29652 13300 31500
rect 13132 29596 13300 29652
rect 13468 29876 13524 29886
rect 13132 28196 13188 29596
rect 13468 29426 13524 29820
rect 13580 29538 13636 32172
rect 14140 32004 14196 32396
rect 13916 31892 13972 31902
rect 14140 31872 14196 31948
rect 13916 31798 13972 31836
rect 13692 31778 13748 31790
rect 13692 31726 13694 31778
rect 13746 31726 13748 31778
rect 13692 30996 13748 31726
rect 14252 31668 14308 33852
rect 14924 33460 14980 36652
rect 15148 36484 15204 36652
rect 15148 36390 15204 36428
rect 15148 34916 15204 34926
rect 15036 34804 15092 34814
rect 15036 34020 15092 34748
rect 15036 33926 15092 33964
rect 14700 33404 14980 33460
rect 15148 33458 15204 34860
rect 15148 33406 15150 33458
rect 15202 33406 15204 33458
rect 14476 32452 14532 32462
rect 14476 32358 14532 32396
rect 14700 32228 14756 33404
rect 15148 33394 15204 33406
rect 15260 32788 15316 36876
rect 15372 36596 15428 39340
rect 15596 39330 15652 39340
rect 15596 38946 15652 38958
rect 15596 38894 15598 38946
rect 15650 38894 15652 38946
rect 15484 38834 15540 38846
rect 15484 38782 15486 38834
rect 15538 38782 15540 38834
rect 15484 38388 15540 38782
rect 15484 38322 15540 38332
rect 15596 38836 15652 38894
rect 15596 37380 15652 38780
rect 15596 37266 15652 37324
rect 15596 37214 15598 37266
rect 15650 37214 15652 37266
rect 15596 37202 15652 37214
rect 15372 36530 15428 36540
rect 15596 36596 15652 36606
rect 15596 36502 15652 36540
rect 15372 35698 15428 35710
rect 15372 35646 15374 35698
rect 15426 35646 15428 35698
rect 15372 35138 15428 35646
rect 15372 35086 15374 35138
rect 15426 35086 15428 35138
rect 15372 35074 15428 35086
rect 15148 32732 15316 32788
rect 14924 32674 14980 32686
rect 14924 32622 14926 32674
rect 14978 32622 14980 32674
rect 14924 32452 14980 32622
rect 15036 32676 15092 32686
rect 15036 32582 15092 32620
rect 13692 30930 13748 30940
rect 13804 31612 14308 31668
rect 14476 32172 14756 32228
rect 14812 32396 14924 32452
rect 13804 30772 13860 31612
rect 13580 29486 13582 29538
rect 13634 29486 13636 29538
rect 13580 29474 13636 29486
rect 13692 30716 13860 30772
rect 13916 30882 13972 30894
rect 14364 30884 14420 30894
rect 13916 30830 13918 30882
rect 13970 30830 13972 30882
rect 13916 30770 13972 30830
rect 13916 30718 13918 30770
rect 13970 30718 13972 30770
rect 13468 29374 13470 29426
rect 13522 29374 13524 29426
rect 13468 29362 13524 29374
rect 13132 28130 13188 28140
rect 13468 28756 13524 28766
rect 13020 28030 13022 28082
rect 13074 28030 13076 28082
rect 13020 28018 13076 28030
rect 12908 27972 12964 27982
rect 12796 27858 12852 27870
rect 12796 27806 12798 27858
rect 12850 27806 12852 27858
rect 12796 27748 12852 27806
rect 12796 27682 12852 27692
rect 12908 27636 12964 27916
rect 13020 27860 13076 27870
rect 13020 27766 13076 27804
rect 13244 27860 13300 27870
rect 13244 27766 13300 27804
rect 13356 27858 13412 27870
rect 13356 27806 13358 27858
rect 13410 27806 13412 27858
rect 13132 27748 13188 27758
rect 13132 27636 13188 27692
rect 12908 27580 13188 27636
rect 12796 27412 12852 27422
rect 12796 26850 12852 27356
rect 12908 27188 12964 27198
rect 12908 27074 12964 27132
rect 12908 27022 12910 27074
rect 12962 27022 12964 27074
rect 12908 27010 12964 27022
rect 13132 26908 13188 27580
rect 13356 27412 13412 27806
rect 13356 27346 13412 27356
rect 13468 27188 13524 28700
rect 13692 27972 13748 30716
rect 13916 30706 13972 30718
rect 14028 30882 14420 30884
rect 14028 30830 14366 30882
rect 14418 30830 14420 30882
rect 14028 30828 14420 30830
rect 13916 30212 13972 30222
rect 13804 30210 13972 30212
rect 13804 30158 13918 30210
rect 13970 30158 13972 30210
rect 13804 30156 13972 30158
rect 13804 28754 13860 30156
rect 13916 30146 13972 30156
rect 13804 28702 13806 28754
rect 13858 28702 13860 28754
rect 13804 28690 13860 28702
rect 14028 28642 14084 30828
rect 14364 30818 14420 30828
rect 14140 30100 14196 30110
rect 14140 30006 14196 30044
rect 14364 30098 14420 30110
rect 14364 30046 14366 30098
rect 14418 30046 14420 30098
rect 14364 29876 14420 30046
rect 14364 29810 14420 29820
rect 14252 29428 14308 29438
rect 14252 29334 14308 29372
rect 14028 28590 14030 28642
rect 14082 28590 14084 28642
rect 14028 28196 14084 28590
rect 14252 28756 14308 28766
rect 14252 28642 14308 28700
rect 14252 28590 14254 28642
rect 14306 28590 14308 28642
rect 14252 28578 14308 28590
rect 14028 28130 14084 28140
rect 14364 28420 14420 28430
rect 14364 28084 14420 28364
rect 14028 27972 14084 27982
rect 13692 27970 14084 27972
rect 13692 27918 14030 27970
rect 14082 27918 14084 27970
rect 13692 27916 14084 27918
rect 14028 27906 14084 27916
rect 14252 27970 14308 27982
rect 14252 27918 14254 27970
rect 14306 27918 14308 27970
rect 14252 27860 14308 27918
rect 14364 27970 14420 28028
rect 14364 27918 14366 27970
rect 14418 27918 14420 27970
rect 14364 27906 14420 27918
rect 14252 27794 14308 27804
rect 13132 26852 13300 26908
rect 12796 26798 12798 26850
rect 12850 26798 12852 26850
rect 12796 26786 12852 26798
rect 12796 26628 12852 26638
rect 12796 26514 12852 26572
rect 12796 26462 12798 26514
rect 12850 26462 12852 26514
rect 12796 25172 12852 26462
rect 12908 26516 12964 26526
rect 12908 26422 12964 26460
rect 13020 26402 13076 26414
rect 13020 26350 13022 26402
rect 13074 26350 13076 26402
rect 12908 25732 12964 25742
rect 12908 25618 12964 25676
rect 12908 25566 12910 25618
rect 12962 25566 12964 25618
rect 12908 25554 12964 25566
rect 13020 25396 13076 26350
rect 13132 26404 13188 26414
rect 13132 26310 13188 26348
rect 13020 25330 13076 25340
rect 12796 25106 12852 25116
rect 12796 24724 12852 24734
rect 12796 24630 12852 24668
rect 12124 21308 12404 21364
rect 12460 23436 12740 23492
rect 13132 23492 13188 23502
rect 12124 19460 12180 21308
rect 12348 20916 12404 20926
rect 12348 20802 12404 20860
rect 12460 20914 12516 23436
rect 13020 23268 13076 23278
rect 12796 23266 13076 23268
rect 12796 23214 13022 23266
rect 13074 23214 13076 23266
rect 12796 23212 13076 23214
rect 12684 22708 12740 22718
rect 12572 22484 12628 22494
rect 12572 22390 12628 22428
rect 12684 21810 12740 22652
rect 12684 21758 12686 21810
rect 12738 21758 12740 21810
rect 12684 21746 12740 21758
rect 12796 20916 12852 23212
rect 13020 23202 13076 23212
rect 13020 22484 13076 22494
rect 13132 22484 13188 23436
rect 13020 22482 13188 22484
rect 13020 22430 13022 22482
rect 13074 22430 13188 22482
rect 13020 22428 13188 22430
rect 13020 22418 13076 22428
rect 12908 21700 12964 21710
rect 12908 21140 12964 21644
rect 12908 21074 12964 21084
rect 13020 21586 13076 21598
rect 13020 21534 13022 21586
rect 13074 21534 13076 21586
rect 13020 21364 13076 21534
rect 12460 20862 12462 20914
rect 12514 20862 12516 20914
rect 12460 20850 12516 20862
rect 12684 20860 12852 20916
rect 12348 20750 12350 20802
rect 12402 20750 12404 20802
rect 12348 20738 12404 20750
rect 12236 20580 12292 20590
rect 12572 20580 12628 20590
rect 12236 20578 12404 20580
rect 12236 20526 12238 20578
rect 12290 20526 12404 20578
rect 12236 20524 12404 20526
rect 12236 20514 12292 20524
rect 12236 20356 12292 20366
rect 12236 20130 12292 20300
rect 12348 20242 12404 20524
rect 12572 20486 12628 20524
rect 12684 20244 12740 20860
rect 12796 20690 12852 20702
rect 12796 20638 12798 20690
rect 12850 20638 12852 20690
rect 12796 20356 12852 20638
rect 12796 20290 12852 20300
rect 12348 20190 12350 20242
rect 12402 20190 12404 20242
rect 12348 20178 12404 20190
rect 12572 20188 12740 20244
rect 12236 20078 12238 20130
rect 12290 20078 12292 20130
rect 12236 20066 12292 20078
rect 12460 20018 12516 20030
rect 12460 19966 12462 20018
rect 12514 19966 12516 20018
rect 12460 19796 12516 19966
rect 12460 19730 12516 19740
rect 12348 19460 12404 19470
rect 12124 19458 12404 19460
rect 12124 19406 12350 19458
rect 12402 19406 12404 19458
rect 12124 19404 12404 19406
rect 12348 19394 12404 19404
rect 12460 19348 12516 19358
rect 12460 19234 12516 19292
rect 12460 19182 12462 19234
rect 12514 19182 12516 19234
rect 12460 18900 12516 19182
rect 12460 18834 12516 18844
rect 12348 18788 12404 18798
rect 12012 18620 12180 18676
rect 11900 18508 12068 18564
rect 11900 18340 11956 18350
rect 11788 18338 11956 18340
rect 11788 18286 11902 18338
rect 11954 18286 11956 18338
rect 11788 18284 11956 18286
rect 11900 18274 11956 18284
rect 11676 18004 11732 18014
rect 11676 17890 11732 17948
rect 11676 17838 11678 17890
rect 11730 17838 11732 17890
rect 11676 17826 11732 17838
rect 11788 17666 11844 17678
rect 11788 17614 11790 17666
rect 11842 17614 11844 17666
rect 11788 15148 11844 17614
rect 11900 17108 11956 17118
rect 11900 17014 11956 17052
rect 12012 16100 12068 18508
rect 12124 17332 12180 18620
rect 12348 18450 12404 18732
rect 12348 18398 12350 18450
rect 12402 18398 12404 18450
rect 12348 18386 12404 18398
rect 12460 18340 12516 18350
rect 12460 17780 12516 18284
rect 12460 17648 12516 17724
rect 12124 17276 12404 17332
rect 12236 16996 12292 17006
rect 12236 16902 12292 16940
rect 12348 16884 12404 17276
rect 12348 16828 12516 16884
rect 12348 16660 12404 16670
rect 12012 16034 12068 16044
rect 12124 16322 12180 16334
rect 12124 16270 12126 16322
rect 12178 16270 12180 16322
rect 12012 15876 12068 15886
rect 12124 15876 12180 16270
rect 12012 15874 12180 15876
rect 12012 15822 12014 15874
rect 12066 15822 12180 15874
rect 12012 15820 12180 15822
rect 12012 15810 12068 15820
rect 12124 15764 12180 15820
rect 12012 15204 12068 15242
rect 11788 15092 11956 15148
rect 12012 15138 12068 15148
rect 11676 14868 11732 14878
rect 11676 13524 11732 14812
rect 11788 14532 11844 14542
rect 11788 14438 11844 14476
rect 11676 13468 11844 13524
rect 11564 13458 11620 13468
rect 10892 12850 11508 12852
rect 10892 12798 10894 12850
rect 10946 12798 11508 12850
rect 10892 12796 11508 12798
rect 11564 12962 11620 12974
rect 11564 12910 11566 12962
rect 11618 12910 11620 12962
rect 9996 9938 10052 9950
rect 9996 9886 9998 9938
rect 10050 9886 10052 9938
rect 9660 9828 9716 9838
rect 9436 8754 9492 8764
rect 9548 9380 9604 9390
rect 9100 5742 9102 5794
rect 9154 5742 9156 5794
rect 9100 4676 9156 5742
rect 9212 6916 9268 6926
rect 9212 5234 9268 6860
rect 9548 6914 9604 9324
rect 9660 7364 9716 9772
rect 9772 9156 9828 9166
rect 9772 9062 9828 9100
rect 9660 7298 9716 7308
rect 9884 8372 9940 8382
rect 9548 6862 9550 6914
rect 9602 6862 9604 6914
rect 9548 6850 9604 6862
rect 9884 6914 9940 8316
rect 9996 8260 10052 9886
rect 9996 8194 10052 8204
rect 9884 6862 9886 6914
rect 9938 6862 9940 6914
rect 9772 6580 9828 6590
rect 9212 5182 9214 5234
rect 9266 5182 9268 5234
rect 9212 5170 9268 5182
rect 9660 5236 9716 5246
rect 9660 5142 9716 5180
rect 9100 4610 9156 4620
rect 8652 3666 8932 3668
rect 8652 3614 8654 3666
rect 8706 3614 8932 3666
rect 8652 3612 8932 3614
rect 8988 4228 9044 4238
rect 8988 3668 9044 4172
rect 8652 3602 8708 3612
rect 8988 3602 9044 3612
rect 9772 3666 9828 6524
rect 9884 5794 9940 6862
rect 10108 6804 10164 10108
rect 10332 9042 10388 9054
rect 10332 8990 10334 9042
rect 10386 8990 10388 9042
rect 10332 8372 10388 8990
rect 10220 8258 10276 8270
rect 10220 8206 10222 8258
rect 10274 8206 10276 8258
rect 10220 7812 10276 8206
rect 10220 7746 10276 7756
rect 10332 7474 10388 8316
rect 10332 7422 10334 7474
rect 10386 7422 10388 7474
rect 10332 7410 10388 7422
rect 9996 6748 10164 6804
rect 10220 7140 10276 7150
rect 9996 6132 10052 6748
rect 10108 6578 10164 6590
rect 10108 6526 10110 6578
rect 10162 6526 10164 6578
rect 10108 6356 10164 6526
rect 10108 6290 10164 6300
rect 10220 6132 10276 7084
rect 9996 6076 10164 6132
rect 9884 5742 9886 5794
rect 9938 5742 9940 5794
rect 9884 5730 9940 5742
rect 9996 5572 10052 5582
rect 9996 4562 10052 5516
rect 10108 5234 10164 6076
rect 10108 5182 10110 5234
rect 10162 5182 10164 5234
rect 10108 5170 10164 5182
rect 10220 4900 10276 6076
rect 10332 6692 10388 6702
rect 10332 6468 10388 6636
rect 10332 6130 10388 6412
rect 10332 6078 10334 6130
rect 10386 6078 10388 6130
rect 10332 6066 10388 6078
rect 10444 5012 10500 10444
rect 10668 9604 10724 10892
rect 10780 10724 10836 10734
rect 10780 10610 10836 10668
rect 10780 10558 10782 10610
rect 10834 10558 10836 10610
rect 10780 10546 10836 10558
rect 10556 7362 10612 7374
rect 10556 7310 10558 7362
rect 10610 7310 10612 7362
rect 10556 7252 10612 7310
rect 10556 7186 10612 7196
rect 10668 6804 10724 9548
rect 10780 9602 10836 9614
rect 10780 9550 10782 9602
rect 10834 9550 10836 9602
rect 10780 8428 10836 9550
rect 10892 9042 10948 12796
rect 11564 12404 11620 12910
rect 11452 12348 11564 12404
rect 11116 12292 11172 12302
rect 11116 12198 11172 12236
rect 11004 12178 11060 12190
rect 11004 12126 11006 12178
rect 11058 12126 11060 12178
rect 11004 12068 11060 12126
rect 11004 12002 11060 12012
rect 11228 12180 11284 12190
rect 10892 8990 10894 9042
rect 10946 8990 10948 9042
rect 10892 8978 10948 8990
rect 11004 11844 11060 11854
rect 10780 8372 10948 8428
rect 10556 6748 10668 6804
rect 10556 6020 10612 6748
rect 10668 6738 10724 6748
rect 10780 8260 10836 8270
rect 10668 6578 10724 6590
rect 10668 6526 10670 6578
rect 10722 6526 10724 6578
rect 10668 6468 10724 6526
rect 10668 6402 10724 6412
rect 10780 6244 10836 8204
rect 10892 7588 10948 8372
rect 10892 7522 10948 7532
rect 11004 7252 11060 11788
rect 11228 11618 11284 12124
rect 11228 11566 11230 11618
rect 11282 11566 11284 11618
rect 11228 11554 11284 11566
rect 10780 6178 10836 6188
rect 10892 7196 11060 7252
rect 11116 11508 11172 11518
rect 10780 6020 10836 6030
rect 10556 6018 10836 6020
rect 10556 5966 10782 6018
rect 10834 5966 10836 6018
rect 10556 5964 10836 5966
rect 10780 5954 10836 5964
rect 10556 5236 10612 5246
rect 10556 5142 10612 5180
rect 10892 5012 10948 7196
rect 11004 6804 11060 6814
rect 11004 6578 11060 6748
rect 11004 6526 11006 6578
rect 11058 6526 11060 6578
rect 11004 6514 11060 6526
rect 11116 6132 11172 11452
rect 11340 11172 11396 11182
rect 10444 4956 10612 5012
rect 10220 4844 10500 4900
rect 9996 4510 9998 4562
rect 10050 4510 10052 4562
rect 9996 4498 10052 4510
rect 10444 4562 10500 4844
rect 10444 4510 10446 4562
rect 10498 4510 10500 4562
rect 10444 4498 10500 4510
rect 10556 4114 10612 4956
rect 10556 4062 10558 4114
rect 10610 4062 10612 4114
rect 10556 4050 10612 4062
rect 10668 4564 10724 4574
rect 9772 3614 9774 3666
rect 9826 3614 9828 3666
rect 9772 3602 9828 3614
rect 10108 3668 10164 3678
rect 10108 3574 10164 3612
rect 10668 3666 10724 4508
rect 10892 4562 10948 4956
rect 10892 4510 10894 4562
rect 10946 4510 10948 4562
rect 10892 4498 10948 4510
rect 11004 6076 11172 6132
rect 11228 11170 11396 11172
rect 11228 11118 11342 11170
rect 11394 11118 11396 11170
rect 11228 11116 11396 11118
rect 11228 10612 11284 11116
rect 11340 11106 11396 11116
rect 11228 9828 11284 10556
rect 11340 10612 11396 10622
rect 11452 10612 11508 12348
rect 11564 12338 11620 12348
rect 11676 12628 11732 12638
rect 11676 12402 11732 12572
rect 11676 12350 11678 12402
rect 11730 12350 11732 12402
rect 11676 12338 11732 12350
rect 11788 11620 11844 13468
rect 11788 11554 11844 11564
rect 11788 11282 11844 11294
rect 11788 11230 11790 11282
rect 11842 11230 11844 11282
rect 11564 11170 11620 11182
rect 11564 11118 11566 11170
rect 11618 11118 11620 11170
rect 11564 10948 11620 11118
rect 11564 10882 11620 10892
rect 11788 10724 11844 11230
rect 11340 10610 11508 10612
rect 11340 10558 11342 10610
rect 11394 10558 11508 10610
rect 11340 10556 11508 10558
rect 11564 10668 11844 10724
rect 11340 9938 11396 10556
rect 11340 9886 11342 9938
rect 11394 9886 11396 9938
rect 11340 9874 11396 9886
rect 10668 3614 10670 3666
rect 10722 3614 10724 3666
rect 10668 3602 10724 3614
rect 11004 3668 11060 6076
rect 11116 5346 11172 5358
rect 11116 5294 11118 5346
rect 11170 5294 11172 5346
rect 11116 5234 11172 5294
rect 11116 5182 11118 5234
rect 11170 5182 11172 5234
rect 11116 5170 11172 5182
rect 11228 4564 11284 9772
rect 11452 7474 11508 7486
rect 11452 7422 11454 7474
rect 11506 7422 11508 7474
rect 11340 6804 11396 6814
rect 11340 6130 11396 6748
rect 11452 6468 11508 7422
rect 11564 7140 11620 10668
rect 11900 9940 11956 15092
rect 12124 15092 12180 15708
rect 12124 15026 12180 15036
rect 12348 15314 12404 16604
rect 12460 16436 12516 16828
rect 12460 16370 12516 16380
rect 12572 16322 12628 20188
rect 12684 20020 12740 20030
rect 12684 19458 12740 19964
rect 12684 19406 12686 19458
rect 12738 19406 12740 19458
rect 12684 19236 12740 19406
rect 12684 19170 12740 19180
rect 12908 19236 12964 19246
rect 12908 19142 12964 19180
rect 13020 18676 13076 21308
rect 13244 20916 13300 26852
rect 13356 26402 13412 26414
rect 13356 26350 13358 26402
rect 13410 26350 13412 26402
rect 13356 25508 13412 26350
rect 13356 25442 13412 25452
rect 13468 25060 13524 27132
rect 13580 27412 13636 27422
rect 13580 26964 13636 27356
rect 14476 27188 14532 32172
rect 14588 32004 14644 32014
rect 14812 32004 14868 32396
rect 14924 32386 14980 32396
rect 14588 32002 14868 32004
rect 14588 31950 14590 32002
rect 14642 31950 14868 32002
rect 14588 31948 14868 31950
rect 14588 31938 14644 31948
rect 15148 31892 15204 32732
rect 15260 32562 15316 32574
rect 15260 32510 15262 32562
rect 15314 32510 15316 32562
rect 15260 32228 15316 32510
rect 15260 32172 15540 32228
rect 15260 31892 15316 31902
rect 15148 31890 15316 31892
rect 15148 31838 15262 31890
rect 15314 31838 15316 31890
rect 15148 31836 15316 31838
rect 15260 31826 15316 31836
rect 14700 31780 14756 31790
rect 15484 31780 15540 32172
rect 15708 32004 15764 41916
rect 16044 41748 16100 41758
rect 16044 41654 16100 41692
rect 16156 41410 16212 43652
rect 16268 43540 16324 43550
rect 16268 43446 16324 43484
rect 16604 43538 16660 43820
rect 16940 43762 16996 44270
rect 17724 44212 17780 44942
rect 17724 44146 17780 44156
rect 17836 44994 18116 44996
rect 17836 44942 18062 44994
rect 18114 44942 18116 44994
rect 17836 44940 18116 44942
rect 17836 44322 17892 44940
rect 18060 44930 18116 44940
rect 17836 44270 17838 44322
rect 17890 44270 17892 44322
rect 17276 44098 17332 44110
rect 17276 44046 17278 44098
rect 17330 44046 17332 44098
rect 17276 43988 17332 44046
rect 17276 43922 17332 43932
rect 16940 43710 16942 43762
rect 16994 43710 16996 43762
rect 16940 43698 16996 43710
rect 17836 43708 17892 44270
rect 16604 43486 16606 43538
rect 16658 43486 16660 43538
rect 16268 42532 16324 42542
rect 16268 42308 16324 42476
rect 16604 42308 16660 43486
rect 16828 43650 16884 43662
rect 16828 43598 16830 43650
rect 16882 43598 16884 43650
rect 16828 42756 16884 43598
rect 17612 43652 17892 43708
rect 16828 42700 17220 42756
rect 17052 42530 17108 42542
rect 17052 42478 17054 42530
rect 17106 42478 17108 42530
rect 16268 42252 16884 42308
rect 16156 41358 16158 41410
rect 16210 41358 16212 41410
rect 16156 41346 16212 41358
rect 16492 42084 16548 42094
rect 15820 41186 15876 41198
rect 15820 41134 15822 41186
rect 15874 41134 15876 41186
rect 15820 40964 15876 41134
rect 16492 41186 16548 42028
rect 16604 42082 16660 42094
rect 16604 42030 16606 42082
rect 16658 42030 16660 42082
rect 16604 41300 16660 42030
rect 16716 41972 16772 41982
rect 16716 41878 16772 41916
rect 16828 41860 16884 42252
rect 17052 42084 17108 42478
rect 17052 42018 17108 42028
rect 17164 42532 17220 42700
rect 16828 41804 17108 41860
rect 16604 41234 16660 41244
rect 16492 41134 16494 41186
rect 16546 41134 16548 41186
rect 16492 41122 16548 41134
rect 15820 40898 15876 40908
rect 16380 40514 16436 40526
rect 16380 40462 16382 40514
rect 16434 40462 16436 40514
rect 16044 40404 16100 40442
rect 16044 40338 16100 40348
rect 16380 40404 16436 40462
rect 16044 40180 16100 40190
rect 16044 39394 16100 40124
rect 16044 39342 16046 39394
rect 16098 39342 16100 39394
rect 16044 39284 16100 39342
rect 15820 38834 15876 38846
rect 15820 38782 15822 38834
rect 15874 38782 15876 38834
rect 15820 38276 15876 38782
rect 16044 38836 16100 39228
rect 16044 38770 16100 38780
rect 16156 38722 16212 38734
rect 16156 38670 16158 38722
rect 16210 38670 16212 38722
rect 16156 38500 16212 38670
rect 16156 38434 16212 38444
rect 15820 38220 16324 38276
rect 16044 37940 16100 37950
rect 16044 37846 16100 37884
rect 16156 37938 16212 37950
rect 16156 37886 16158 37938
rect 16210 37886 16212 37938
rect 15820 37826 15876 37838
rect 15820 37774 15822 37826
rect 15874 37774 15876 37826
rect 15820 36596 15876 37774
rect 15932 37828 15988 37838
rect 15932 37734 15988 37772
rect 16156 37828 16212 37886
rect 16268 37938 16324 38220
rect 16268 37886 16270 37938
rect 16322 37886 16324 37938
rect 16268 37874 16324 37886
rect 16156 37762 16212 37772
rect 16380 37492 16436 40348
rect 16940 40402 16996 40414
rect 16940 40350 16942 40402
rect 16994 40350 16996 40402
rect 16940 40180 16996 40350
rect 16940 40114 16996 40124
rect 16828 39394 16884 39406
rect 16828 39342 16830 39394
rect 16882 39342 16884 39394
rect 16828 38946 16884 39342
rect 16828 38894 16830 38946
rect 16882 38894 16884 38946
rect 16604 38836 16660 38846
rect 16604 38742 16660 38780
rect 16828 38668 16884 38894
rect 16940 39396 16996 39406
rect 16940 38946 16996 39340
rect 16940 38894 16942 38946
rect 16994 38894 16996 38946
rect 16940 38882 16996 38894
rect 16716 38612 16996 38668
rect 16044 37268 16100 37278
rect 16044 37044 16100 37212
rect 16044 36988 16212 37044
rect 15820 36530 15876 36540
rect 16044 36484 16100 36494
rect 16044 35586 16100 36428
rect 16044 35534 16046 35586
rect 16098 35534 16100 35586
rect 15820 34802 15876 34814
rect 15820 34750 15822 34802
rect 15874 34750 15876 34802
rect 15820 34244 15876 34750
rect 15932 34804 15988 34814
rect 15932 34710 15988 34748
rect 16044 34802 16100 35534
rect 16044 34750 16046 34802
rect 16098 34750 16100 34802
rect 15820 34188 15988 34244
rect 15820 34020 15876 34030
rect 15820 33926 15876 33964
rect 15932 33908 15988 34188
rect 15932 33842 15988 33852
rect 15932 33684 15988 33694
rect 15820 33572 15876 33582
rect 15820 32450 15876 33516
rect 15820 32398 15822 32450
rect 15874 32398 15876 32450
rect 15820 32386 15876 32398
rect 15708 31948 15876 32004
rect 15708 31780 15764 31790
rect 15484 31778 15764 31780
rect 15484 31726 15710 31778
rect 15762 31726 15764 31778
rect 15484 31724 15764 31726
rect 14700 31218 14756 31724
rect 15708 31714 15764 31724
rect 14700 31166 14702 31218
rect 14754 31166 14756 31218
rect 14700 31154 14756 31166
rect 15260 30882 15316 30894
rect 15260 30830 15262 30882
rect 15314 30830 15316 30882
rect 14700 30770 14756 30782
rect 14700 30718 14702 30770
rect 14754 30718 14756 30770
rect 14588 30098 14644 30110
rect 14588 30046 14590 30098
rect 14642 30046 14644 30098
rect 14588 29428 14644 30046
rect 14588 29362 14644 29372
rect 14700 28532 14756 30718
rect 15148 30100 15204 30110
rect 15148 30006 15204 30044
rect 15260 29876 15316 30830
rect 15372 30548 15428 30558
rect 15372 30434 15428 30492
rect 15372 30382 15374 30434
rect 15426 30382 15428 30434
rect 15372 30370 15428 30382
rect 15708 30436 15764 30446
rect 15820 30436 15876 31948
rect 15708 30434 15876 30436
rect 15708 30382 15710 30434
rect 15762 30382 15876 30434
rect 15708 30380 15876 30382
rect 15708 30370 15764 30380
rect 15260 29810 15316 29820
rect 15820 29540 15876 29550
rect 15708 29426 15764 29438
rect 15708 29374 15710 29426
rect 15762 29374 15764 29426
rect 15596 29316 15652 29326
rect 14588 28476 14756 28532
rect 15484 28644 15540 28654
rect 14588 27860 14644 28476
rect 14588 27794 14644 27804
rect 14700 28308 14756 28318
rect 14588 27188 14644 27198
rect 14476 27186 14644 27188
rect 14476 27134 14590 27186
rect 14642 27134 14644 27186
rect 14476 27132 14644 27134
rect 14588 27122 14644 27132
rect 14700 27074 14756 28252
rect 15484 28308 15540 28588
rect 15596 28530 15652 29260
rect 15708 29204 15764 29374
rect 15708 29138 15764 29148
rect 15596 28478 15598 28530
rect 15650 28478 15652 28530
rect 15596 28466 15652 28478
rect 15820 28530 15876 29484
rect 15820 28478 15822 28530
rect 15874 28478 15876 28530
rect 15820 28466 15876 28478
rect 15260 27860 15316 27870
rect 15260 27766 15316 27804
rect 15484 27748 15540 28252
rect 15708 28418 15764 28430
rect 15708 28366 15710 28418
rect 15762 28366 15764 28418
rect 15708 27972 15764 28366
rect 15708 27906 15764 27916
rect 15820 28196 15876 28206
rect 15708 27748 15764 27758
rect 15484 27746 15764 27748
rect 15484 27694 15710 27746
rect 15762 27694 15764 27746
rect 15484 27692 15764 27694
rect 15708 27682 15764 27692
rect 15148 27634 15204 27646
rect 15148 27582 15150 27634
rect 15202 27582 15204 27634
rect 14924 27412 14980 27422
rect 14924 27186 14980 27356
rect 15148 27298 15204 27582
rect 15148 27246 15150 27298
rect 15202 27246 15204 27298
rect 15148 27234 15204 27246
rect 14924 27134 14926 27186
rect 14978 27134 14980 27186
rect 14924 27122 14980 27134
rect 14700 27022 14702 27074
rect 14754 27022 14756 27074
rect 14700 27010 14756 27022
rect 15372 27076 15428 27086
rect 13580 26898 13636 26908
rect 13804 26964 13860 27002
rect 15372 26982 15428 27020
rect 14476 26962 14532 26974
rect 14476 26910 14478 26962
rect 14530 26910 14532 26962
rect 14476 26908 14532 26910
rect 13804 26898 13860 26908
rect 14364 26852 14532 26908
rect 14588 26964 14644 26974
rect 14588 26852 14756 26908
rect 14364 26292 14420 26852
rect 14700 26514 14756 26852
rect 15596 26852 15652 26862
rect 14700 26462 14702 26514
rect 14754 26462 14756 26514
rect 14700 26450 14756 26462
rect 14924 26740 14980 26750
rect 14588 26404 14644 26414
rect 14588 26310 14644 26348
rect 14364 26226 14420 26236
rect 14476 26180 14532 26190
rect 14476 26086 14532 26124
rect 14364 25956 14420 25966
rect 14364 25508 14420 25900
rect 14476 25620 14532 25630
rect 14476 25526 14532 25564
rect 14140 25506 14420 25508
rect 14140 25454 14366 25506
rect 14418 25454 14420 25506
rect 14140 25452 14420 25454
rect 14028 25396 14084 25406
rect 14028 25302 14084 25340
rect 13692 25284 13748 25294
rect 13692 25282 13860 25284
rect 13692 25230 13694 25282
rect 13746 25230 13860 25282
rect 13692 25228 13860 25230
rect 13692 25218 13748 25228
rect 13356 25004 13524 25060
rect 13356 24052 13412 25004
rect 13468 24722 13524 24734
rect 13468 24670 13470 24722
rect 13522 24670 13524 24722
rect 13468 24612 13524 24670
rect 13468 24276 13524 24556
rect 13468 24210 13524 24220
rect 13804 24164 13860 25228
rect 13916 25282 13972 25294
rect 13916 25230 13918 25282
rect 13970 25230 13972 25282
rect 13916 25172 13972 25230
rect 13916 25106 13972 25116
rect 14028 24724 14084 24734
rect 14140 24724 14196 25452
rect 14364 25442 14420 25452
rect 14476 25396 14532 25406
rect 14476 25284 14532 25340
rect 14028 24722 14196 24724
rect 14028 24670 14030 24722
rect 14082 24670 14196 24722
rect 14028 24668 14196 24670
rect 14364 25228 14532 25284
rect 14028 24658 14084 24668
rect 13356 23996 13524 24052
rect 13468 23380 13524 23996
rect 13804 24050 13860 24108
rect 13804 23998 13806 24050
rect 13858 23998 13860 24050
rect 13804 23986 13860 23998
rect 13916 23940 13972 23950
rect 13804 23828 13860 23838
rect 13804 23734 13860 23772
rect 13468 23314 13524 23324
rect 13580 23156 13636 23166
rect 13356 23154 13636 23156
rect 13356 23102 13582 23154
rect 13634 23102 13636 23154
rect 13356 23100 13636 23102
rect 13356 21924 13412 23100
rect 13580 23090 13636 23100
rect 13356 21858 13412 21868
rect 13468 22596 13524 22606
rect 13468 21252 13524 22540
rect 13804 22484 13860 22494
rect 13916 22484 13972 23884
rect 13804 22482 13972 22484
rect 13804 22430 13806 22482
rect 13858 22430 13972 22482
rect 13804 22428 13972 22430
rect 14028 23826 14084 23838
rect 14028 23774 14030 23826
rect 14082 23774 14084 23826
rect 13804 22418 13860 22428
rect 13916 22148 13972 22158
rect 13244 20850 13300 20860
rect 13356 21196 13524 21252
rect 13580 21476 13636 21486
rect 13580 21252 13636 21420
rect 13020 18610 13076 18620
rect 13132 19348 13188 19358
rect 12684 18452 12740 18462
rect 12684 17108 12740 18396
rect 12796 18338 12852 18350
rect 12796 18286 12798 18338
rect 12850 18286 12852 18338
rect 12796 17220 12852 18286
rect 12908 18226 12964 18238
rect 12908 18174 12910 18226
rect 12962 18174 12964 18226
rect 12908 17778 12964 18174
rect 12908 17726 12910 17778
rect 12962 17726 12964 17778
rect 12908 17668 12964 17726
rect 12908 17602 12964 17612
rect 12796 17164 12964 17220
rect 12684 17042 12740 17052
rect 12796 16884 12852 16894
rect 12572 16270 12574 16322
rect 12626 16270 12628 16322
rect 12572 16258 12628 16270
rect 12684 16882 12852 16884
rect 12684 16830 12798 16882
rect 12850 16830 12852 16882
rect 12684 16828 12852 16830
rect 12572 15874 12628 15886
rect 12572 15822 12574 15874
rect 12626 15822 12628 15874
rect 12572 15652 12628 15822
rect 12572 15586 12628 15596
rect 12348 15262 12350 15314
rect 12402 15262 12404 15314
rect 12124 14756 12180 14766
rect 12124 14662 12180 14700
rect 12012 14420 12068 14430
rect 12012 14326 12068 14364
rect 12124 13746 12180 13758
rect 12124 13694 12126 13746
rect 12178 13694 12180 13746
rect 12012 13636 12068 13646
rect 12012 12180 12068 13580
rect 12124 13412 12180 13694
rect 12124 13346 12180 13356
rect 12348 13300 12404 15262
rect 12684 14756 12740 16828
rect 12796 16818 12852 16828
rect 12908 16660 12964 17164
rect 13132 17108 13188 19292
rect 13356 18564 13412 21196
rect 13580 20914 13636 21196
rect 13580 20862 13582 20914
rect 13634 20862 13636 20914
rect 13580 20850 13636 20862
rect 13692 21028 13748 21038
rect 13692 19906 13748 20972
rect 13692 19854 13694 19906
rect 13746 19854 13748 19906
rect 13244 18508 13412 18564
rect 13468 19572 13524 19582
rect 13244 18226 13300 18508
rect 13356 18340 13412 18350
rect 13356 18246 13412 18284
rect 13244 18174 13246 18226
rect 13298 18174 13300 18226
rect 13244 17556 13300 18174
rect 13468 17780 13524 19516
rect 13692 19012 13748 19854
rect 13804 19908 13860 19918
rect 13804 19814 13860 19852
rect 13916 19572 13972 22092
rect 14028 21812 14084 23774
rect 14252 22708 14308 22718
rect 14252 22370 14308 22652
rect 14252 22318 14254 22370
rect 14306 22318 14308 22370
rect 14252 22260 14308 22318
rect 14252 22194 14308 22204
rect 14140 21812 14196 21822
rect 14028 21756 14140 21812
rect 14140 21474 14196 21756
rect 14140 21422 14142 21474
rect 14194 21422 14196 21474
rect 14028 20020 14084 20030
rect 14028 19926 14084 19964
rect 14140 19796 14196 21422
rect 14252 21362 14308 21374
rect 14252 21310 14254 21362
rect 14306 21310 14308 21362
rect 14252 20914 14308 21310
rect 14252 20862 14254 20914
rect 14306 20862 14308 20914
rect 14252 20850 14308 20862
rect 14364 20804 14420 25228
rect 14812 24612 14868 24622
rect 14924 24612 14980 26684
rect 15484 26404 15540 26414
rect 15260 26402 15540 26404
rect 15260 26350 15486 26402
rect 15538 26350 15540 26402
rect 15260 26348 15540 26350
rect 15260 25508 15316 26348
rect 15484 26338 15540 26348
rect 15596 26404 15652 26796
rect 15596 26272 15652 26348
rect 15484 26068 15540 26078
rect 15484 25974 15540 26012
rect 15260 25506 15428 25508
rect 15260 25454 15262 25506
rect 15314 25454 15428 25506
rect 15260 25452 15428 25454
rect 15260 25442 15316 25452
rect 15036 25394 15092 25406
rect 15036 25342 15038 25394
rect 15090 25342 15092 25394
rect 15036 25284 15092 25342
rect 15036 25228 15204 25284
rect 15148 25060 15204 25228
rect 15148 24994 15204 25004
rect 15260 25172 15316 25182
rect 14812 24610 14980 24612
rect 14812 24558 14814 24610
rect 14866 24558 14980 24610
rect 14812 24556 14980 24558
rect 15036 24836 15092 24846
rect 14812 24546 14868 24556
rect 14476 24276 14532 24286
rect 14476 21362 14532 24220
rect 14700 23938 14756 23950
rect 14700 23886 14702 23938
rect 14754 23886 14756 23938
rect 14700 23828 14756 23886
rect 14588 23268 14644 23278
rect 14588 23174 14644 23212
rect 14588 22260 14644 22270
rect 14700 22260 14756 23772
rect 14924 23828 14980 23838
rect 14924 23714 14980 23772
rect 14924 23662 14926 23714
rect 14978 23662 14980 23714
rect 14812 23156 14868 23166
rect 14812 23062 14868 23100
rect 14588 22258 14756 22260
rect 14588 22206 14590 22258
rect 14642 22206 14756 22258
rect 14588 22204 14756 22206
rect 14588 22148 14644 22204
rect 14588 22082 14644 22092
rect 14700 21588 14756 21598
rect 14700 21494 14756 21532
rect 14924 21588 14980 23662
rect 15036 22260 15092 24780
rect 15148 24610 15204 24622
rect 15148 24558 15150 24610
rect 15202 24558 15204 24610
rect 15148 24276 15204 24558
rect 15260 24388 15316 25116
rect 15260 24322 15316 24332
rect 15148 23716 15204 24220
rect 15372 23938 15428 25452
rect 15484 25282 15540 25294
rect 15484 25230 15486 25282
rect 15538 25230 15540 25282
rect 15484 25172 15540 25230
rect 15484 25106 15540 25116
rect 15596 25282 15652 25294
rect 15596 25230 15598 25282
rect 15650 25230 15652 25282
rect 15596 24836 15652 25230
rect 15372 23886 15374 23938
rect 15426 23886 15428 23938
rect 15372 23874 15428 23886
rect 15484 24780 15652 24836
rect 15708 25060 15764 25070
rect 15708 24836 15764 25004
rect 15148 23650 15204 23660
rect 15036 22194 15092 22204
rect 15148 23380 15204 23390
rect 15148 23156 15204 23324
rect 15260 23268 15316 23278
rect 15260 23174 15316 23212
rect 15148 22146 15204 23100
rect 15148 22094 15150 22146
rect 15202 22094 15204 22146
rect 14924 21586 15092 21588
rect 14924 21534 14926 21586
rect 14978 21534 15092 21586
rect 14924 21532 15092 21534
rect 14924 21522 14980 21532
rect 14476 21310 14478 21362
rect 14530 21310 14532 21362
rect 14476 21298 14532 21310
rect 14812 21474 14868 21486
rect 14812 21422 14814 21474
rect 14866 21422 14868 21474
rect 14812 20916 14868 21422
rect 14700 20860 14868 20916
rect 14588 20804 14644 20814
rect 14364 20748 14532 20804
rect 14252 20692 14308 20702
rect 14252 20598 14308 20636
rect 14364 20578 14420 20590
rect 14364 20526 14366 20578
rect 14418 20526 14420 20578
rect 13916 19506 13972 19516
rect 14028 19740 14196 19796
rect 14252 19796 14308 19806
rect 13916 19348 13972 19358
rect 13804 19236 13860 19274
rect 13916 19254 13972 19292
rect 13804 19170 13860 19180
rect 13692 18956 13860 19012
rect 13804 18562 13860 18956
rect 13916 18788 13972 18798
rect 13916 18674 13972 18732
rect 13916 18622 13918 18674
rect 13970 18622 13972 18674
rect 13916 18610 13972 18622
rect 13804 18510 13806 18562
rect 13858 18510 13860 18562
rect 13804 18498 13860 18510
rect 13468 17714 13524 17724
rect 13580 18228 13636 18238
rect 14028 18228 14084 19740
rect 14252 19458 14308 19740
rect 14252 19406 14254 19458
rect 14306 19406 14308 19458
rect 14140 19234 14196 19246
rect 14140 19182 14142 19234
rect 14194 19182 14196 19234
rect 14140 19124 14196 19182
rect 14140 19058 14196 19068
rect 14252 19012 14308 19406
rect 14252 18946 14308 18956
rect 14140 18452 14196 18462
rect 14364 18452 14420 20526
rect 14140 18450 14420 18452
rect 14140 18398 14142 18450
rect 14194 18398 14420 18450
rect 14140 18396 14420 18398
rect 14140 18386 14196 18396
rect 14476 18340 14532 20748
rect 14588 20710 14644 20748
rect 14700 20244 14756 20860
rect 14812 20690 14868 20702
rect 14812 20638 14814 20690
rect 14866 20638 14868 20690
rect 14812 20580 14868 20638
rect 14812 20514 14868 20524
rect 14700 20178 14756 20188
rect 15036 20130 15092 21532
rect 15036 20078 15038 20130
rect 15090 20078 15092 20130
rect 15036 20066 15092 20078
rect 14700 19908 14756 19918
rect 14700 19460 14756 19852
rect 14700 18674 14756 19404
rect 14700 18622 14702 18674
rect 14754 18622 14756 18674
rect 14924 19236 14980 19246
rect 14700 18610 14756 18622
rect 14812 18618 14868 18630
rect 14812 18566 14814 18618
rect 14866 18566 14868 18618
rect 14476 18284 14644 18340
rect 14028 18172 14532 18228
rect 13244 17500 13524 17556
rect 13132 17052 13412 17108
rect 13244 16884 13300 16894
rect 13244 16790 13300 16828
rect 12908 16594 12964 16604
rect 12908 16212 12964 16222
rect 12908 16118 12964 16156
rect 13356 16212 13412 17052
rect 13356 16146 13412 16156
rect 13020 16100 13076 16110
rect 13020 15538 13076 16044
rect 13020 15486 13022 15538
rect 13074 15486 13076 15538
rect 13020 15474 13076 15486
rect 13132 15876 13188 15886
rect 12908 15428 12964 15438
rect 12908 15314 12964 15372
rect 12908 15262 12910 15314
rect 12962 15262 12964 15314
rect 12908 15250 12964 15262
rect 13020 15204 13076 15214
rect 12684 14690 12740 14700
rect 12908 14756 12964 14766
rect 13020 14756 13076 15148
rect 12908 14754 13076 14756
rect 12908 14702 12910 14754
rect 12962 14702 13076 14754
rect 12908 14700 13076 14702
rect 12908 14690 12964 14700
rect 12908 14532 12964 14542
rect 13132 14532 13188 15820
rect 12908 14530 13188 14532
rect 12908 14478 12910 14530
rect 12962 14478 13188 14530
rect 12908 14476 13188 14478
rect 13356 15652 13412 15662
rect 12908 14466 12964 14476
rect 12572 14418 12628 14430
rect 12572 14366 12574 14418
rect 12626 14366 12628 14418
rect 12572 14084 12628 14366
rect 12348 13234 12404 13244
rect 12460 14028 12572 14084
rect 12236 12404 12292 12414
rect 12236 12310 12292 12348
rect 12012 12124 12180 12180
rect 12012 11620 12068 11630
rect 12012 10834 12068 11564
rect 12012 10782 12014 10834
rect 12066 10782 12068 10834
rect 12012 10770 12068 10782
rect 11900 9874 11956 9884
rect 12012 9604 12068 9614
rect 12124 9604 12180 12124
rect 12460 11508 12516 14028
rect 12572 14018 12628 14028
rect 12796 14308 12852 14318
rect 12684 12852 12740 12862
rect 12796 12852 12852 14252
rect 13244 14084 13300 14094
rect 12740 12850 12852 12852
rect 12740 12798 12798 12850
rect 12850 12798 12852 12850
rect 12740 12796 12852 12798
rect 12684 12786 12740 12796
rect 12796 12786 12852 12796
rect 12908 12962 12964 12974
rect 12908 12910 12910 12962
rect 12962 12910 12964 12962
rect 12908 12852 12964 12910
rect 12908 12786 12964 12796
rect 12572 12628 12628 12638
rect 12572 12402 12628 12572
rect 13020 12628 13076 12638
rect 12572 12350 12574 12402
rect 12626 12350 12628 12402
rect 12572 12338 12628 12350
rect 12796 12516 12852 12526
rect 11900 9602 12180 9604
rect 11900 9550 12014 9602
rect 12066 9550 12180 9602
rect 11900 9548 12180 9550
rect 12236 11452 12516 11508
rect 12796 12292 12852 12460
rect 11676 9268 11732 9278
rect 11676 9174 11732 9212
rect 11676 8372 11732 8382
rect 11676 7924 11732 8316
rect 11788 8148 11844 8158
rect 11788 8054 11844 8092
rect 11676 7858 11732 7868
rect 11564 7074 11620 7084
rect 11788 7700 11844 7710
rect 11564 6804 11620 6814
rect 11788 6804 11844 7644
rect 11564 6802 11844 6804
rect 11564 6750 11566 6802
rect 11618 6750 11844 6802
rect 11564 6748 11844 6750
rect 11564 6738 11620 6748
rect 11452 6402 11508 6412
rect 11340 6078 11342 6130
rect 11394 6078 11396 6130
rect 11340 5346 11396 6078
rect 11340 5294 11342 5346
rect 11394 5294 11396 5346
rect 11340 5282 11396 5294
rect 11564 5236 11620 5246
rect 11228 4498 11284 4508
rect 11340 5124 11396 5134
rect 11228 4340 11284 4350
rect 11340 4340 11396 5068
rect 11228 4338 11396 4340
rect 11228 4286 11230 4338
rect 11282 4286 11396 4338
rect 11228 4284 11396 4286
rect 11228 4274 11284 4284
rect 11340 4228 11396 4284
rect 11340 4162 11396 4172
rect 11116 3668 11172 3678
rect 11004 3666 11172 3668
rect 11004 3614 11118 3666
rect 11170 3614 11172 3666
rect 11004 3612 11172 3614
rect 11116 3602 11172 3612
rect 11564 3556 11620 5180
rect 11788 5012 11844 6748
rect 11900 5236 11956 9548
rect 12012 9538 12068 9548
rect 12236 9268 12292 11452
rect 12348 11284 12404 11294
rect 12404 11228 12516 11284
rect 12348 11190 12404 11228
rect 12012 9212 12292 9268
rect 12348 10610 12404 10622
rect 12348 10558 12350 10610
rect 12402 10558 12404 10610
rect 12012 7700 12068 9212
rect 12012 7634 12068 7644
rect 12236 9044 12292 9054
rect 12124 7588 12180 7598
rect 12124 7494 12180 7532
rect 12236 7028 12292 8988
rect 12348 8260 12404 10558
rect 12348 7252 12404 8204
rect 12348 7186 12404 7196
rect 12460 7700 12516 11228
rect 12684 11170 12740 11182
rect 12684 11118 12686 11170
rect 12738 11118 12740 11170
rect 12684 10052 12740 11118
rect 12796 10834 12852 12236
rect 12796 10782 12798 10834
rect 12850 10782 12852 10834
rect 12796 10770 12852 10782
rect 12908 11844 12964 11854
rect 12684 9986 12740 9996
rect 12796 9940 12852 9950
rect 12572 9602 12628 9614
rect 12572 9550 12574 9602
rect 12626 9550 12628 9602
rect 12572 9154 12628 9550
rect 12572 9102 12574 9154
rect 12626 9102 12628 9154
rect 12572 9044 12628 9102
rect 12572 8978 12628 8988
rect 12796 8370 12852 9884
rect 12908 9714 12964 11788
rect 12908 9662 12910 9714
rect 12962 9662 12964 9714
rect 12908 9650 12964 9662
rect 13020 9492 13076 12572
rect 13132 12404 13188 12414
rect 13132 12310 13188 12348
rect 12796 8318 12798 8370
rect 12850 8318 12852 8370
rect 12796 8306 12852 8318
rect 12908 9436 13076 9492
rect 12236 6972 12404 7028
rect 12236 6804 12292 6814
rect 12236 6710 12292 6748
rect 12124 6692 12180 6702
rect 12012 6636 12124 6692
rect 12012 5906 12068 6636
rect 12124 6598 12180 6636
rect 12236 6132 12292 6142
rect 12348 6132 12404 6972
rect 12236 6130 12404 6132
rect 12236 6078 12238 6130
rect 12290 6078 12404 6130
rect 12236 6076 12404 6078
rect 12236 6066 12292 6076
rect 12012 5854 12014 5906
rect 12066 5854 12068 5906
rect 12012 5842 12068 5854
rect 12460 5572 12516 7644
rect 12460 5506 12516 5516
rect 12684 7588 12740 7598
rect 12684 7362 12740 7532
rect 12684 7310 12686 7362
rect 12738 7310 12740 7362
rect 11900 5170 11956 5180
rect 12348 5348 12404 5358
rect 12236 5124 12292 5134
rect 12012 5122 12292 5124
rect 12012 5070 12238 5122
rect 12290 5070 12292 5122
rect 12012 5068 12292 5070
rect 12012 5012 12068 5068
rect 12236 5058 12292 5068
rect 11788 4956 12068 5012
rect 12348 4562 12404 5292
rect 12348 4510 12350 4562
rect 12402 4510 12404 4562
rect 12348 4498 12404 4510
rect 12684 4340 12740 7310
rect 12908 6690 12964 9436
rect 13244 9266 13300 14028
rect 13356 13188 13412 15596
rect 13468 14532 13524 17500
rect 13580 16994 13636 18172
rect 13916 17780 13972 17790
rect 13804 17668 13860 17678
rect 13804 17444 13860 17612
rect 13804 17378 13860 17388
rect 13580 16942 13582 16994
rect 13634 16942 13636 16994
rect 13580 16930 13636 16942
rect 13916 16884 13972 17724
rect 14028 17668 14084 17678
rect 14364 17668 14420 17678
rect 14028 17666 14308 17668
rect 14028 17614 14030 17666
rect 14082 17614 14308 17666
rect 14028 17612 14308 17614
rect 14028 17602 14084 17612
rect 13916 16882 14196 16884
rect 13916 16830 13918 16882
rect 13970 16830 14196 16882
rect 13916 16828 14196 16830
rect 13916 16818 13972 16828
rect 13916 15986 13972 15998
rect 13916 15934 13918 15986
rect 13970 15934 13972 15986
rect 13580 15874 13636 15886
rect 13580 15822 13582 15874
rect 13634 15822 13636 15874
rect 13580 15428 13636 15822
rect 13804 15876 13860 15914
rect 13804 15810 13860 15820
rect 13580 15362 13636 15372
rect 13804 15652 13860 15662
rect 13692 15314 13748 15326
rect 13692 15262 13694 15314
rect 13746 15262 13748 15314
rect 13692 14868 13748 15262
rect 13692 14802 13748 14812
rect 13804 15092 13860 15596
rect 13692 14532 13748 14542
rect 13468 14530 13748 14532
rect 13468 14478 13694 14530
rect 13746 14478 13748 14530
rect 13468 14476 13748 14478
rect 13692 14466 13748 14476
rect 13804 14308 13860 15036
rect 13692 14306 13860 14308
rect 13692 14254 13806 14306
rect 13858 14254 13860 14306
rect 13692 14252 13860 14254
rect 13692 14084 13748 14252
rect 13804 14242 13860 14252
rect 13916 14418 13972 15934
rect 14028 15314 14084 15326
rect 14028 15262 14030 15314
rect 14082 15262 14084 15314
rect 14028 14756 14084 15262
rect 14028 14690 14084 14700
rect 13916 14366 13918 14418
rect 13970 14366 13972 14418
rect 13692 14018 13748 14028
rect 13916 14084 13972 14366
rect 13468 13972 13524 13982
rect 13468 13748 13524 13916
rect 13468 13746 13748 13748
rect 13468 13694 13470 13746
rect 13522 13694 13748 13746
rect 13468 13692 13748 13694
rect 13468 13682 13524 13692
rect 13356 13122 13412 13132
rect 13580 13412 13636 13422
rect 13468 12292 13524 12302
rect 13468 12198 13524 12236
rect 13580 11396 13636 13356
rect 13468 11394 13636 11396
rect 13468 11342 13582 11394
rect 13634 11342 13636 11394
rect 13468 11340 13636 11342
rect 13356 10612 13412 10622
rect 13356 10518 13412 10556
rect 13244 9214 13246 9266
rect 13298 9214 13300 9266
rect 13244 9202 13300 9214
rect 12908 6638 12910 6690
rect 12962 6638 12964 6690
rect 12908 6356 12964 6638
rect 12908 6290 12964 6300
rect 13020 7362 13076 7374
rect 13020 7310 13022 7362
rect 13074 7310 13076 7362
rect 13020 6692 13076 7310
rect 12796 6132 12852 6142
rect 13020 6132 13076 6636
rect 12796 6130 13076 6132
rect 12796 6078 12798 6130
rect 12850 6078 13076 6130
rect 12796 6076 13076 6078
rect 13244 6356 13300 6366
rect 12796 6066 12852 6076
rect 13132 6020 13188 6030
rect 13132 5926 13188 5964
rect 13244 5908 13300 6300
rect 13244 5842 13300 5852
rect 13468 5682 13524 11340
rect 13580 11330 13636 11340
rect 13692 9492 13748 13692
rect 13804 12740 13860 12750
rect 13804 12646 13860 12684
rect 13916 12628 13972 14028
rect 14140 13972 14196 16828
rect 14252 15764 14308 17612
rect 14364 17574 14420 17612
rect 14476 17444 14532 18172
rect 14364 17388 14532 17444
rect 14364 16212 14420 17388
rect 14476 17108 14532 17118
rect 14476 16994 14532 17052
rect 14476 16942 14478 16994
rect 14530 16942 14532 16994
rect 14476 16930 14532 16942
rect 14476 16212 14532 16222
rect 14364 16210 14532 16212
rect 14364 16158 14478 16210
rect 14530 16158 14532 16210
rect 14364 16156 14532 16158
rect 14476 16146 14532 16156
rect 14252 14980 14308 15708
rect 14588 15204 14644 18284
rect 14700 18228 14756 18238
rect 14700 15540 14756 18172
rect 14812 17108 14868 18566
rect 14924 17892 14980 19180
rect 15148 18452 15204 22094
rect 15372 22370 15428 22382
rect 15372 22318 15374 22370
rect 15426 22318 15428 22370
rect 15372 21924 15428 22318
rect 15372 21858 15428 21868
rect 15372 21588 15428 21598
rect 15372 21494 15428 21532
rect 15484 21476 15540 24780
rect 15596 24612 15652 24622
rect 15708 24612 15764 24780
rect 15596 24610 15764 24612
rect 15596 24558 15598 24610
rect 15650 24558 15764 24610
rect 15596 24556 15764 24558
rect 15596 24546 15652 24556
rect 15708 23826 15764 23838
rect 15708 23774 15710 23826
rect 15762 23774 15764 23826
rect 15596 23716 15652 23726
rect 15596 23622 15652 23660
rect 15708 23492 15764 23774
rect 15596 23436 15764 23492
rect 15596 23044 15652 23436
rect 15708 23266 15764 23278
rect 15708 23214 15710 23266
rect 15762 23214 15764 23266
rect 15708 23156 15764 23214
rect 15708 23090 15764 23100
rect 15596 22708 15652 22988
rect 15596 22642 15652 22652
rect 15820 22708 15876 28140
rect 15932 27634 15988 33628
rect 16044 33460 16100 34750
rect 16156 34356 16212 36988
rect 16268 36596 16324 36606
rect 16380 36596 16436 37436
rect 16492 38500 16548 38510
rect 16492 36932 16548 38444
rect 16604 37828 16660 37838
rect 16604 37154 16660 37772
rect 16604 37102 16606 37154
rect 16658 37102 16660 37154
rect 16604 37090 16660 37102
rect 16716 37378 16772 38612
rect 16940 38546 16996 38556
rect 16716 37326 16718 37378
rect 16770 37326 16772 37378
rect 16716 37156 16772 37326
rect 16716 37100 16884 37156
rect 16492 36876 16660 36932
rect 16268 36594 16436 36596
rect 16268 36542 16270 36594
rect 16322 36542 16436 36594
rect 16268 36540 16436 36542
rect 16268 36530 16324 36540
rect 16492 36260 16548 36270
rect 16492 34916 16548 36204
rect 16604 35922 16660 36876
rect 16828 36596 16884 37100
rect 16940 37042 16996 37054
rect 16940 36990 16942 37042
rect 16994 36990 16996 37042
rect 16940 36820 16996 36990
rect 16940 36754 16996 36764
rect 16716 36540 16884 36596
rect 16716 36482 16772 36540
rect 16716 36430 16718 36482
rect 16770 36430 16772 36482
rect 16716 36418 16772 36430
rect 17052 36484 17108 41804
rect 17164 39508 17220 42476
rect 17612 42530 17668 43652
rect 17836 43586 17892 43596
rect 17948 44772 18004 44782
rect 17612 42478 17614 42530
rect 17666 42478 17668 42530
rect 17612 42308 17668 42478
rect 17612 42242 17668 42252
rect 17724 41858 17780 41870
rect 17724 41806 17726 41858
rect 17778 41806 17780 41858
rect 17724 41746 17780 41806
rect 17724 41694 17726 41746
rect 17778 41694 17780 41746
rect 17612 41188 17668 41198
rect 17724 41188 17780 41694
rect 17612 41186 17780 41188
rect 17612 41134 17614 41186
rect 17666 41134 17780 41186
rect 17612 41132 17780 41134
rect 17836 41300 17892 41310
rect 17612 40516 17668 41132
rect 17612 40450 17668 40460
rect 17724 40404 17780 40414
rect 17724 40310 17780 40348
rect 17164 39442 17220 39452
rect 17612 40178 17668 40190
rect 17612 40126 17614 40178
rect 17666 40126 17668 40178
rect 17276 39396 17332 39406
rect 17612 39396 17668 40126
rect 17276 39394 17668 39396
rect 17276 39342 17278 39394
rect 17330 39342 17668 39394
rect 17276 39340 17668 39342
rect 17276 39330 17332 39340
rect 17164 38724 17220 38734
rect 17164 36820 17220 38668
rect 17388 38500 17444 38510
rect 17388 38162 17444 38444
rect 17388 38110 17390 38162
rect 17442 38110 17444 38162
rect 17388 38098 17444 38110
rect 17612 38052 17668 39340
rect 17836 39618 17892 41244
rect 17836 39566 17838 39618
rect 17890 39566 17892 39618
rect 17724 38836 17780 38846
rect 17724 38742 17780 38780
rect 17612 37958 17668 37996
rect 17724 38388 17780 38398
rect 17724 37156 17780 38332
rect 17724 37062 17780 37100
rect 17164 36754 17220 36764
rect 17052 36418 17108 36428
rect 17276 36370 17332 36382
rect 17276 36318 17278 36370
rect 17330 36318 17332 36370
rect 17164 36260 17220 36270
rect 16604 35870 16606 35922
rect 16658 35870 16660 35922
rect 16604 35858 16660 35870
rect 16940 36258 17220 36260
rect 16940 36206 17166 36258
rect 17218 36206 17220 36258
rect 16940 36204 17220 36206
rect 16940 35922 16996 36204
rect 17164 36036 17220 36204
rect 17276 36260 17332 36318
rect 17276 36194 17332 36204
rect 17724 36260 17780 36270
rect 17724 36166 17780 36204
rect 17164 35980 17780 36036
rect 16940 35870 16942 35922
rect 16994 35870 16996 35922
rect 16492 34850 16548 34860
rect 16940 34914 16996 35870
rect 17724 35922 17780 35980
rect 17724 35870 17726 35922
rect 17778 35870 17780 35922
rect 17724 35858 17780 35870
rect 17836 35700 17892 39566
rect 17948 39172 18004 44716
rect 18172 44324 18228 44334
rect 18060 44098 18116 44110
rect 18060 44046 18062 44098
rect 18114 44046 18116 44098
rect 18060 43762 18116 44046
rect 18060 43710 18062 43762
rect 18114 43710 18116 43762
rect 18060 43698 18116 43710
rect 18172 43540 18228 44268
rect 18284 43708 18340 46284
rect 18396 46274 18452 46284
rect 18508 46786 18564 46798
rect 18508 46734 18510 46786
rect 18562 46734 18564 46786
rect 18508 45556 18564 46734
rect 18620 46676 18676 46686
rect 18620 46582 18676 46620
rect 18508 45490 18564 45500
rect 18508 45108 18564 45118
rect 18508 45014 18564 45052
rect 18732 45108 18788 45118
rect 18396 44212 18452 44222
rect 18396 44118 18452 44156
rect 18620 43876 18676 43886
rect 18284 43652 18452 43708
rect 18396 43650 18452 43652
rect 18396 43598 18398 43650
rect 18450 43598 18452 43650
rect 18396 43586 18452 43598
rect 18508 43652 18564 43662
rect 18508 43558 18564 43596
rect 18284 43540 18340 43550
rect 18172 43538 18340 43540
rect 18172 43486 18286 43538
rect 18338 43486 18340 43538
rect 18172 43484 18340 43486
rect 18060 42532 18116 42542
rect 18060 42438 18116 42476
rect 18060 41972 18116 41982
rect 18060 41878 18116 41916
rect 18284 41748 18340 43484
rect 18620 42084 18676 43820
rect 18732 42644 18788 45052
rect 18844 44212 18900 44222
rect 18844 43540 18900 44156
rect 18956 43876 19012 47068
rect 19068 46452 19124 46462
rect 19068 45780 19124 46396
rect 19180 46340 19236 46350
rect 19180 46114 19236 46284
rect 19180 46062 19182 46114
rect 19234 46062 19236 46114
rect 19180 46050 19236 46062
rect 19068 45332 19124 45724
rect 19292 45666 19348 47406
rect 19292 45614 19294 45666
rect 19346 45614 19348 45666
rect 19292 45556 19348 45614
rect 19292 45490 19348 45500
rect 19180 45332 19236 45342
rect 19068 45330 19236 45332
rect 19068 45278 19182 45330
rect 19234 45278 19236 45330
rect 19068 45276 19236 45278
rect 19068 45106 19124 45118
rect 19068 45054 19070 45106
rect 19122 45054 19124 45106
rect 19068 44324 19124 45054
rect 19068 44258 19124 44268
rect 18956 43810 19012 43820
rect 19068 43540 19124 43550
rect 18844 43538 19124 43540
rect 18844 43486 19070 43538
rect 19122 43486 19124 43538
rect 18844 43484 19124 43486
rect 18844 42866 18900 43484
rect 19068 43474 19124 43484
rect 18844 42814 18846 42866
rect 18898 42814 18900 42866
rect 18844 42802 18900 42814
rect 18732 42588 19012 42644
rect 18284 41298 18340 41692
rect 18284 41246 18286 41298
rect 18338 41246 18340 41298
rect 18284 41234 18340 41246
rect 18508 42028 18676 42084
rect 18844 42420 18900 42430
rect 18172 40292 18228 40302
rect 18060 39396 18116 39406
rect 18060 39302 18116 39340
rect 17948 39116 18116 39172
rect 17948 38948 18004 38958
rect 17948 38834 18004 38892
rect 18060 38946 18116 39116
rect 18060 38894 18062 38946
rect 18114 38894 18116 38946
rect 18060 38882 18116 38894
rect 17948 38782 17950 38834
rect 18002 38782 18004 38834
rect 17948 38724 18004 38782
rect 18172 38724 18228 40236
rect 18284 40290 18340 40302
rect 18284 40238 18286 40290
rect 18338 40238 18340 40290
rect 18284 40178 18340 40238
rect 18284 40126 18286 40178
rect 18338 40126 18340 40178
rect 18284 40114 18340 40126
rect 18508 39172 18564 42028
rect 18620 41858 18676 41870
rect 18620 41806 18622 41858
rect 18674 41806 18676 41858
rect 18620 41746 18676 41806
rect 18620 41694 18622 41746
rect 18674 41694 18676 41746
rect 18620 41682 18676 41694
rect 18844 41188 18900 42364
rect 18956 41972 19012 42588
rect 19180 42532 19236 45276
rect 19404 45330 19460 47964
rect 19516 47796 19572 48078
rect 19516 47730 19572 47740
rect 19628 47682 19684 48860
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 21196 48468 21252 49646
rect 21196 48374 21252 48412
rect 19628 47630 19630 47682
rect 19682 47630 19684 47682
rect 19404 45278 19406 45330
rect 19458 45278 19460 45330
rect 19404 45266 19460 45278
rect 19516 47570 19572 47582
rect 19516 47518 19518 47570
rect 19570 47518 19572 47570
rect 19516 46676 19572 47518
rect 19516 45778 19572 46620
rect 19628 46674 19684 47630
rect 19740 48242 19796 48254
rect 19740 48190 19742 48242
rect 19794 48190 19796 48242
rect 19740 47572 19796 48190
rect 19740 47506 19796 47516
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 19628 46622 19630 46674
rect 19682 46622 19684 46674
rect 19628 46610 19684 46622
rect 19740 46564 19796 46574
rect 19740 46470 19796 46508
rect 20188 46452 20244 46462
rect 20188 46358 20244 46396
rect 19516 45726 19518 45778
rect 19570 45726 19572 45778
rect 19516 44324 19572 45726
rect 19964 45780 20020 45790
rect 19964 45686 20020 45724
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20300 45332 20356 45342
rect 21420 45332 21476 56028
rect 27020 56082 27076 56094
rect 27020 56030 27022 56082
rect 27074 56030 27076 56082
rect 27020 55972 27076 56030
rect 27020 55906 27076 55916
rect 27580 55972 27636 55982
rect 27580 55878 27636 55916
rect 23660 55860 23716 55870
rect 23324 55186 23380 55198
rect 23324 55134 23326 55186
rect 23378 55134 23380 55186
rect 22876 55076 22932 55086
rect 22876 54982 22932 55020
rect 23324 55076 23380 55134
rect 23660 55186 23716 55804
rect 27132 55300 27188 55310
rect 26796 55188 26852 55198
rect 23660 55134 23662 55186
rect 23714 55134 23716 55186
rect 23660 55122 23716 55134
rect 26572 55186 26852 55188
rect 26572 55134 26798 55186
rect 26850 55134 26852 55186
rect 26572 55132 26852 55134
rect 23324 55010 23380 55020
rect 23548 51604 23604 51614
rect 24668 51604 24724 51614
rect 23548 51602 24724 51604
rect 23548 51550 23550 51602
rect 23602 51550 24670 51602
rect 24722 51550 24724 51602
rect 23548 51548 24724 51550
rect 23548 51538 23604 51548
rect 24668 51538 24724 51548
rect 26236 51490 26292 51502
rect 26236 51438 26238 51490
rect 26290 51438 26292 51490
rect 23436 51378 23492 51390
rect 23436 51326 23438 51378
rect 23490 51326 23492 51378
rect 21868 51266 21924 51278
rect 21868 51214 21870 51266
rect 21922 51214 21924 51266
rect 21532 49812 21588 49822
rect 21532 49718 21588 49756
rect 21756 49140 21812 49150
rect 21756 49046 21812 49084
rect 21644 49028 21700 49038
rect 21644 48934 21700 48972
rect 21868 48916 21924 51214
rect 22204 50594 22260 50606
rect 22204 50542 22206 50594
rect 22258 50542 22260 50594
rect 22204 49812 22260 50542
rect 22540 50594 22596 50606
rect 22540 50542 22542 50594
rect 22594 50542 22596 50594
rect 22540 50372 22596 50542
rect 22764 50596 22820 50606
rect 22764 50502 22820 50540
rect 23212 50372 23268 50382
rect 22540 50370 23268 50372
rect 22540 50318 23214 50370
rect 23266 50318 23268 50370
rect 22540 50316 23268 50318
rect 22204 49746 22260 49756
rect 22428 49812 22484 49822
rect 22428 49718 22484 49756
rect 22540 49586 22596 50316
rect 23212 50306 23268 50316
rect 23436 49812 23492 51326
rect 23660 51378 23716 51390
rect 23660 51326 23662 51378
rect 23714 51326 23716 51378
rect 23660 50372 23716 51326
rect 24108 51380 24164 51390
rect 24108 51286 24164 51324
rect 24556 51378 24612 51390
rect 24556 51326 24558 51378
rect 24610 51326 24612 51378
rect 24220 51156 24276 51166
rect 24108 50596 24164 50606
rect 23660 50306 23716 50316
rect 23772 50594 24164 50596
rect 23772 50542 24110 50594
rect 24162 50542 24164 50594
rect 23772 50540 24164 50542
rect 23660 49812 23716 49822
rect 23492 49810 23716 49812
rect 23492 49758 23662 49810
rect 23714 49758 23716 49810
rect 23492 49756 23716 49758
rect 23436 49746 23492 49756
rect 23436 49588 23492 49598
rect 22540 49534 22542 49586
rect 22594 49534 22596 49586
rect 21980 48916 22036 48926
rect 21868 48914 22036 48916
rect 21868 48862 21982 48914
rect 22034 48862 22036 48914
rect 21868 48860 22036 48862
rect 21868 48468 21924 48860
rect 21980 48850 22036 48860
rect 21868 48374 21924 48412
rect 22428 48802 22484 48814
rect 22428 48750 22430 48802
rect 22482 48750 22484 48802
rect 22428 48468 22484 48750
rect 22540 48804 22596 49534
rect 23324 49532 23436 49588
rect 23324 49028 23380 49532
rect 23436 49456 23492 49532
rect 23436 49252 23492 49262
rect 23548 49252 23604 49756
rect 23660 49746 23716 49756
rect 23436 49250 23604 49252
rect 23436 49198 23438 49250
rect 23490 49198 23604 49250
rect 23436 49196 23604 49198
rect 23772 49250 23828 50540
rect 24108 50530 24164 50540
rect 23772 49198 23774 49250
rect 23826 49198 23828 49250
rect 23436 49186 23492 49196
rect 23772 49186 23828 49198
rect 23996 50372 24052 50382
rect 23996 49810 24052 50316
rect 24220 49922 24276 51100
rect 24220 49870 24222 49922
rect 24274 49870 24276 49922
rect 24220 49858 24276 49870
rect 23996 49758 23998 49810
rect 24050 49758 24052 49810
rect 23660 49140 23716 49150
rect 23324 48972 23604 49028
rect 22876 48804 22932 48814
rect 22540 48802 22932 48804
rect 22540 48750 22878 48802
rect 22930 48750 22932 48802
rect 22540 48748 22932 48750
rect 21980 48356 22036 48366
rect 21980 48262 22036 48300
rect 22316 48356 22372 48366
rect 21868 48018 21924 48030
rect 21868 47966 21870 48018
rect 21922 47966 21924 48018
rect 21868 47460 21924 47966
rect 22316 47682 22372 48300
rect 22428 48132 22484 48412
rect 22428 48066 22484 48076
rect 22316 47630 22318 47682
rect 22370 47630 22372 47682
rect 22316 47618 22372 47630
rect 22876 47572 22932 48748
rect 23212 48242 23268 48254
rect 23212 48190 23214 48242
rect 23266 48190 23268 48242
rect 23212 48132 23268 48190
rect 23436 48244 23492 48254
rect 23436 48150 23492 48188
rect 23212 48066 23268 48076
rect 23548 48130 23604 48972
rect 23660 48914 23716 49084
rect 23996 49140 24052 49758
rect 24108 49588 24164 49598
rect 24556 49588 24612 51326
rect 24108 49586 24612 49588
rect 24108 49534 24110 49586
rect 24162 49534 24612 49586
rect 24108 49532 24612 49534
rect 24668 51380 24724 51390
rect 24668 50706 24724 51324
rect 24668 50654 24670 50706
rect 24722 50654 24724 50706
rect 24668 49588 24724 50654
rect 24108 49522 24164 49532
rect 24668 49522 24724 49532
rect 24892 51378 24948 51390
rect 24892 51326 24894 51378
rect 24946 51326 24948 51378
rect 23996 49074 24052 49084
rect 23660 48862 23662 48914
rect 23714 48862 23716 48914
rect 23660 48850 23716 48862
rect 24892 48804 24948 51326
rect 26124 51156 26180 51166
rect 26124 51062 26180 51100
rect 26124 50932 26180 50942
rect 26124 50594 26180 50876
rect 26124 50542 26126 50594
rect 26178 50542 26180 50594
rect 25004 50482 25060 50494
rect 25004 50430 25006 50482
rect 25058 50430 25060 50482
rect 25004 49924 25060 50430
rect 25004 49858 25060 49868
rect 25228 50484 25284 50494
rect 24892 48738 24948 48748
rect 24332 48356 24388 48366
rect 24332 48262 24388 48300
rect 24108 48244 24164 48254
rect 24108 48150 24164 48188
rect 24444 48242 24500 48254
rect 24444 48190 24446 48242
rect 24498 48190 24500 48242
rect 23548 48078 23550 48130
rect 23602 48078 23604 48130
rect 23548 48066 23604 48078
rect 22876 47570 23268 47572
rect 22876 47518 22878 47570
rect 22930 47518 23268 47570
rect 22876 47516 23268 47518
rect 22876 47506 22932 47516
rect 22652 47460 22708 47470
rect 21868 47394 21924 47404
rect 22540 47458 22708 47460
rect 22540 47406 22654 47458
rect 22706 47406 22708 47458
rect 22540 47404 22708 47406
rect 22540 46674 22596 47404
rect 22652 47394 22708 47404
rect 22988 47348 23044 47358
rect 22652 46900 22708 46910
rect 22652 46806 22708 46844
rect 22876 46900 22932 46910
rect 22988 46900 23044 47292
rect 22876 46898 23044 46900
rect 22876 46846 22878 46898
rect 22930 46846 23044 46898
rect 22876 46844 23044 46846
rect 23212 46900 23268 47516
rect 23436 47460 23492 47470
rect 23436 47366 23492 47404
rect 23772 47460 23828 47470
rect 23772 47366 23828 47404
rect 23548 47348 23604 47358
rect 23548 47254 23604 47292
rect 24444 47348 24500 48190
rect 24892 48132 24948 48142
rect 24892 48038 24948 48076
rect 24444 47282 24500 47292
rect 24892 47796 24948 47806
rect 22876 46834 22932 46844
rect 23212 46806 23268 46844
rect 24108 47234 24164 47246
rect 24108 47182 24110 47234
rect 24162 47182 24164 47234
rect 24108 46900 24164 47182
rect 22540 46622 22542 46674
rect 22594 46622 22596 46674
rect 22540 46116 22596 46622
rect 23324 46676 23380 46686
rect 22540 46060 22708 46116
rect 20300 45330 20468 45332
rect 20300 45278 20302 45330
rect 20354 45278 20468 45330
rect 20300 45276 20468 45278
rect 20300 45266 20356 45276
rect 19964 45108 20020 45118
rect 19964 45014 20020 45052
rect 20300 44996 20356 45006
rect 20300 44902 20356 44940
rect 20188 44882 20244 44894
rect 20188 44830 20190 44882
rect 20242 44830 20244 44882
rect 20188 44660 20244 44830
rect 20188 44604 20356 44660
rect 19740 44324 19796 44334
rect 19516 44322 19796 44324
rect 19516 44270 19742 44322
rect 19794 44270 19796 44322
rect 19516 44268 19796 44270
rect 19740 44258 19796 44268
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19180 42466 19236 42476
rect 19404 43762 19460 43774
rect 19404 43710 19406 43762
rect 19458 43710 19460 43762
rect 19404 43540 19460 43710
rect 20300 43708 20356 44604
rect 20412 44322 20468 45276
rect 21420 45266 21476 45276
rect 20972 45220 21028 45230
rect 20412 44270 20414 44322
rect 20466 44270 20468 44322
rect 20412 44258 20468 44270
rect 20524 44996 20580 45006
rect 20524 43708 20580 44940
rect 20860 44996 20916 45006
rect 20860 44902 20916 44940
rect 20636 44436 20692 44446
rect 20636 44434 20916 44436
rect 20636 44382 20638 44434
rect 20690 44382 20916 44434
rect 20636 44380 20916 44382
rect 20636 44370 20692 44380
rect 20300 43652 20468 43708
rect 20524 43652 20804 43708
rect 20300 43540 20356 43550
rect 19404 43484 20300 43540
rect 18956 41970 19348 41972
rect 18956 41918 18958 41970
rect 19010 41918 19348 41970
rect 18956 41916 19348 41918
rect 18956 41906 19012 41916
rect 18844 41132 19012 41188
rect 18844 40962 18900 40974
rect 18844 40910 18846 40962
rect 18898 40910 18900 40962
rect 18732 40402 18788 40414
rect 18732 40350 18734 40402
rect 18786 40350 18788 40402
rect 18732 40292 18788 40350
rect 18844 40404 18900 40910
rect 18844 40338 18900 40348
rect 18732 40226 18788 40236
rect 18956 39956 19012 41132
rect 19292 41186 19348 41916
rect 19404 41860 19460 43484
rect 20300 43446 20356 43484
rect 20076 43314 20132 43326
rect 20076 43262 20078 43314
rect 20130 43262 20132 43314
rect 20076 42980 20132 43262
rect 20412 43316 20468 43652
rect 20636 43316 20692 43326
rect 20412 43314 20692 43316
rect 20412 43262 20638 43314
rect 20690 43262 20692 43314
rect 20412 43260 20692 43262
rect 20300 42980 20356 42990
rect 20076 42978 20356 42980
rect 20076 42926 20302 42978
rect 20354 42926 20356 42978
rect 20076 42924 20356 42926
rect 20300 42914 20356 42924
rect 19516 42754 19572 42766
rect 20524 42756 20580 42766
rect 19516 42702 19518 42754
rect 19570 42702 19572 42754
rect 19516 42644 19572 42702
rect 19516 42196 19572 42588
rect 20412 42754 20580 42756
rect 20412 42702 20526 42754
rect 20578 42702 20580 42754
rect 20412 42700 20580 42702
rect 20412 42642 20468 42700
rect 20524 42690 20580 42700
rect 20412 42590 20414 42642
rect 20466 42590 20468 42642
rect 20412 42578 20468 42590
rect 19740 42532 19796 42570
rect 19740 42466 19796 42476
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19964 42196 20020 42206
rect 19516 42194 20020 42196
rect 19516 42142 19966 42194
rect 20018 42142 20020 42194
rect 19516 42140 20020 42142
rect 19964 42130 20020 42140
rect 20188 42196 20244 42206
rect 20636 42196 20692 43260
rect 20748 42756 20804 43652
rect 20860 43316 20916 44380
rect 20972 43762 21028 45164
rect 20972 43710 20974 43762
rect 21026 43710 21028 43762
rect 20972 43698 21028 43710
rect 22428 43764 22484 43774
rect 21420 43540 21476 43550
rect 21420 43446 21476 43484
rect 22316 43428 22372 43438
rect 22428 43428 22484 43708
rect 22652 43708 22708 46060
rect 23324 46114 23380 46620
rect 23324 46062 23326 46114
rect 23378 46062 23380 46114
rect 23324 46050 23380 46062
rect 22876 46002 22932 46014
rect 22876 45950 22878 46002
rect 22930 45950 22932 46002
rect 22876 45218 22932 45950
rect 22876 45166 22878 45218
rect 22930 45166 22932 45218
rect 22876 44660 22932 45166
rect 22988 45890 23044 45902
rect 22988 45838 22990 45890
rect 23042 45838 23044 45890
rect 22988 45220 23044 45838
rect 23212 45892 23268 45902
rect 23212 45330 23268 45836
rect 23212 45278 23214 45330
rect 23266 45278 23268 45330
rect 23212 45266 23268 45278
rect 22988 45126 23044 45164
rect 22876 44604 23268 44660
rect 23212 44434 23268 44604
rect 23212 44382 23214 44434
rect 23266 44382 23268 44434
rect 23212 44370 23268 44382
rect 22764 44324 22820 44334
rect 23100 44324 23156 44334
rect 22764 44322 22932 44324
rect 22764 44270 22766 44322
rect 22818 44270 22932 44322
rect 22764 44268 22932 44270
rect 22764 44258 22820 44268
rect 22876 43708 22932 44268
rect 23100 43764 23156 44268
rect 23660 44324 23716 44334
rect 23660 44230 23716 44268
rect 24108 43708 24164 46844
rect 24892 46898 24948 47740
rect 24892 46846 24894 46898
rect 24946 46846 24948 46898
rect 24892 46834 24948 46846
rect 24220 46674 24276 46686
rect 24220 46622 24222 46674
rect 24274 46622 24276 46674
rect 24220 45892 24276 46622
rect 24668 46676 24724 46686
rect 24668 46582 24724 46620
rect 24780 46562 24836 46574
rect 24780 46510 24782 46562
rect 24834 46510 24836 46562
rect 24780 46004 24836 46510
rect 24780 45938 24836 45948
rect 25004 46228 25060 46238
rect 24220 45826 24276 45836
rect 24892 45892 24948 45902
rect 24892 45798 24948 45836
rect 24220 45444 24276 45454
rect 24220 44546 24276 45388
rect 24220 44494 24222 44546
rect 24274 44494 24276 44546
rect 24220 44482 24276 44494
rect 24668 44436 24724 44446
rect 24332 44324 24388 44334
rect 22652 43652 22820 43708
rect 22876 43652 23044 43708
rect 23100 43652 23268 43708
rect 24108 43652 24276 43708
rect 22316 43426 22484 43428
rect 22316 43374 22318 43426
rect 22370 43374 22484 43426
rect 22316 43372 22484 43374
rect 22316 43362 22372 43372
rect 20860 43222 20916 43260
rect 21196 43204 21252 43214
rect 20748 42754 20916 42756
rect 20748 42702 20750 42754
rect 20802 42702 20916 42754
rect 20748 42700 20916 42702
rect 20748 42690 20804 42700
rect 20860 42642 20916 42700
rect 20860 42590 20862 42642
rect 20914 42590 20916 42642
rect 20188 42102 20244 42140
rect 20412 42140 20692 42196
rect 20748 42532 20804 42542
rect 20748 42194 20804 42476
rect 20748 42142 20750 42194
rect 20802 42142 20804 42194
rect 19852 41972 19908 41982
rect 19404 41794 19460 41804
rect 19516 41970 19908 41972
rect 19516 41918 19854 41970
rect 19906 41918 19908 41970
rect 19516 41916 19908 41918
rect 19292 41134 19294 41186
rect 19346 41134 19348 41186
rect 19292 41122 19348 41134
rect 19516 40626 19572 41916
rect 19852 41906 19908 41916
rect 19628 40964 19684 40974
rect 19628 40870 19684 40908
rect 20188 40962 20244 40974
rect 20188 40910 20190 40962
rect 20242 40910 20244 40962
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19516 40574 19518 40626
rect 19570 40574 19572 40626
rect 19516 40562 19572 40574
rect 19404 40516 19460 40526
rect 19404 40422 19460 40460
rect 19292 40404 19348 40414
rect 19292 40310 19348 40348
rect 19740 40402 19796 40414
rect 19740 40350 19742 40402
rect 19794 40350 19796 40402
rect 18844 39900 19012 39956
rect 18620 39396 18676 39406
rect 18620 39394 18788 39396
rect 18620 39342 18622 39394
rect 18674 39342 18788 39394
rect 18620 39340 18788 39342
rect 18620 39330 18676 39340
rect 18508 39116 18676 39172
rect 17948 38668 18228 38724
rect 18284 38610 18340 38622
rect 18284 38558 18286 38610
rect 18338 38558 18340 38610
rect 17948 37826 18004 37838
rect 17948 37774 17950 37826
rect 18002 37774 18004 37826
rect 17948 37716 18004 37774
rect 18284 37716 18340 38558
rect 18508 38610 18564 38622
rect 18508 38558 18510 38610
rect 18562 38558 18564 38610
rect 18508 38274 18564 38558
rect 18508 38222 18510 38274
rect 18562 38222 18564 38274
rect 18508 38210 18564 38222
rect 18620 38052 18676 39116
rect 18732 38388 18788 39340
rect 18732 38322 18788 38332
rect 18844 38164 18900 39900
rect 19628 39844 19684 39854
rect 19740 39844 19796 40350
rect 20188 40068 20244 40910
rect 20300 40404 20356 40414
rect 20300 40310 20356 40348
rect 20412 40292 20468 42140
rect 20748 42130 20804 42142
rect 20636 41970 20692 41982
rect 20636 41918 20638 41970
rect 20690 41918 20692 41970
rect 20636 40626 20692 41918
rect 20748 41748 20804 41758
rect 20748 41654 20804 41692
rect 20860 41524 20916 42590
rect 20636 40574 20638 40626
rect 20690 40574 20692 40626
rect 20636 40562 20692 40574
rect 20748 41468 20916 41524
rect 20524 40516 20580 40526
rect 20524 40422 20580 40460
rect 20412 40236 20692 40292
rect 20188 40012 20580 40068
rect 19628 39842 19796 39844
rect 19628 39790 19630 39842
rect 19682 39790 19796 39842
rect 19628 39788 19796 39790
rect 19628 39778 19684 39788
rect 18956 39732 19012 39742
rect 18956 38836 19012 39676
rect 20524 39732 20580 40012
rect 19964 39620 20020 39630
rect 19404 39508 19460 39518
rect 19068 39394 19124 39406
rect 19068 39342 19070 39394
rect 19122 39342 19124 39394
rect 19068 39060 19124 39342
rect 19404 39060 19460 39452
rect 19964 39396 20020 39564
rect 20188 39508 20244 39518
rect 20188 39414 20244 39452
rect 20524 39506 20580 39676
rect 20524 39454 20526 39506
rect 20578 39454 20580 39506
rect 20524 39442 20580 39454
rect 19964 39330 20020 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19068 39004 19460 39060
rect 19180 38836 19236 38846
rect 18956 38834 19236 38836
rect 18956 38782 19182 38834
rect 19234 38782 19236 38834
rect 18956 38780 19236 38782
rect 19180 38500 19236 38780
rect 19180 38434 19236 38444
rect 18508 37996 18676 38052
rect 18732 38108 18900 38164
rect 17948 37660 18452 37716
rect 18172 37492 18228 37502
rect 18060 37380 18116 37390
rect 17388 35644 17892 35700
rect 17948 36484 18004 36494
rect 17388 35026 17444 35644
rect 17388 34974 17390 35026
rect 17442 34974 17444 35026
rect 17388 34962 17444 34974
rect 16940 34862 16942 34914
rect 16994 34862 16996 34914
rect 16940 34850 16996 34862
rect 16268 34356 16324 34366
rect 16156 34354 16324 34356
rect 16156 34302 16270 34354
rect 16322 34302 16324 34354
rect 16156 34300 16324 34302
rect 16268 34290 16324 34300
rect 16604 34356 16660 34366
rect 16604 34020 16660 34300
rect 17948 34242 18004 36428
rect 18060 35812 18116 37324
rect 18172 37154 18228 37436
rect 18396 37266 18452 37660
rect 18396 37214 18398 37266
rect 18450 37214 18452 37266
rect 18396 37202 18452 37214
rect 18172 37102 18174 37154
rect 18226 37102 18228 37154
rect 18172 37044 18228 37102
rect 18172 36978 18228 36988
rect 18172 36820 18228 36830
rect 18172 36260 18228 36764
rect 18172 36258 18452 36260
rect 18172 36206 18174 36258
rect 18226 36206 18452 36258
rect 18172 36204 18452 36206
rect 18172 36194 18228 36204
rect 18060 35810 18228 35812
rect 18060 35758 18062 35810
rect 18114 35758 18228 35810
rect 18060 35756 18228 35758
rect 18060 35746 18116 35756
rect 17948 34190 17950 34242
rect 18002 34190 18004 34242
rect 17948 34178 18004 34190
rect 18172 34244 18228 35756
rect 18172 34178 18228 34188
rect 18284 35588 18340 35598
rect 18284 35138 18340 35532
rect 18284 35086 18286 35138
rect 18338 35086 18340 35138
rect 16604 33954 16660 33964
rect 18060 34130 18116 34142
rect 18060 34078 18062 34130
rect 18114 34078 18116 34130
rect 16044 33394 16100 33404
rect 17612 33796 17668 33806
rect 17612 33458 17668 33740
rect 18060 33796 18116 34078
rect 18060 33730 18116 33740
rect 17612 33406 17614 33458
rect 17666 33406 17668 33458
rect 17612 33394 17668 33406
rect 16156 33124 16212 33134
rect 16044 33122 16212 33124
rect 16044 33070 16158 33122
rect 16210 33070 16212 33122
rect 16044 33068 16212 33070
rect 16044 31892 16100 33068
rect 16156 33058 16212 33068
rect 16268 33122 16324 33134
rect 16268 33070 16270 33122
rect 16322 33070 16324 33122
rect 16156 32564 16212 32574
rect 16156 32228 16212 32508
rect 16268 32450 16324 33070
rect 16380 33122 16436 33134
rect 16604 33124 16660 33134
rect 16380 33070 16382 33122
rect 16434 33070 16436 33122
rect 16380 32564 16436 33070
rect 16492 33068 16604 33124
rect 16492 32676 16548 33068
rect 16604 33030 16660 33068
rect 17276 33122 17332 33134
rect 17276 33070 17278 33122
rect 17330 33070 17332 33122
rect 16492 32610 16548 32620
rect 16380 32498 16436 32508
rect 16604 32562 16660 32574
rect 16604 32510 16606 32562
rect 16658 32510 16660 32562
rect 16268 32398 16270 32450
rect 16322 32398 16324 32450
rect 16268 32386 16324 32398
rect 16156 32162 16212 32172
rect 16044 31798 16100 31836
rect 16156 32004 16212 32014
rect 16044 30884 16100 30894
rect 16044 30790 16100 30828
rect 15932 27582 15934 27634
rect 15986 27582 15988 27634
rect 15932 27570 15988 27582
rect 16044 28644 16100 28654
rect 16044 28082 16100 28588
rect 16044 28030 16046 28082
rect 16098 28030 16100 28082
rect 16044 27636 16100 28030
rect 16044 27570 16100 27580
rect 15932 27298 15988 27310
rect 15932 27246 15934 27298
rect 15986 27246 15988 27298
rect 15932 26850 15988 27246
rect 15932 26798 15934 26850
rect 15986 26798 15988 26850
rect 15932 25172 15988 26798
rect 16044 25284 16100 25294
rect 16044 25190 16100 25228
rect 15932 25106 15988 25116
rect 16044 24610 16100 24622
rect 16044 24558 16046 24610
rect 16098 24558 16100 24610
rect 16044 24388 16100 24558
rect 16044 23492 16100 24332
rect 16044 23426 16100 23436
rect 15820 22642 15876 22652
rect 16044 23268 16100 23278
rect 16044 22594 16100 23212
rect 16044 22542 16046 22594
rect 16098 22542 16100 22594
rect 16044 22530 16100 22542
rect 15932 22258 15988 22270
rect 15932 22206 15934 22258
rect 15986 22206 15988 22258
rect 15708 22148 15764 22158
rect 15708 21700 15764 22092
rect 15708 21634 15764 21644
rect 15820 21924 15876 21934
rect 15820 21698 15876 21868
rect 15820 21646 15822 21698
rect 15874 21646 15876 21698
rect 15820 21634 15876 21646
rect 15484 21420 15652 21476
rect 15372 21028 15428 21038
rect 15372 20914 15428 20972
rect 15372 20862 15374 20914
rect 15426 20862 15428 20914
rect 15372 20850 15428 20862
rect 15372 19572 15428 19582
rect 15372 19346 15428 19516
rect 15484 19460 15540 19470
rect 15484 19366 15540 19404
rect 15372 19294 15374 19346
rect 15426 19294 15428 19346
rect 15372 19282 15428 19294
rect 15260 19124 15316 19134
rect 15260 19030 15316 19068
rect 15596 18788 15652 21420
rect 15820 21140 15876 21150
rect 15820 20914 15876 21084
rect 15820 20862 15822 20914
rect 15874 20862 15876 20914
rect 15820 20850 15876 20862
rect 15484 18732 15652 18788
rect 15708 20132 15764 20142
rect 15372 18564 15428 18574
rect 15372 18470 15428 18508
rect 15148 18396 15316 18452
rect 14924 17826 14980 17836
rect 15148 17668 15204 17678
rect 15148 17574 15204 17612
rect 15036 17108 15092 17118
rect 14868 17106 15092 17108
rect 14868 17054 15038 17106
rect 15090 17054 15092 17106
rect 14868 17052 15092 17054
rect 14812 16976 14868 17052
rect 15036 17042 15092 17052
rect 14700 15474 14756 15484
rect 14924 16772 14980 16782
rect 14924 15316 14980 16716
rect 15260 16212 15316 18396
rect 15372 18004 15428 18014
rect 15372 17106 15428 17948
rect 15484 17778 15540 18732
rect 15708 18676 15764 20076
rect 15932 19908 15988 22206
rect 16044 22146 16100 22158
rect 16044 22094 16046 22146
rect 16098 22094 16100 22146
rect 16044 22036 16100 22094
rect 16044 21364 16100 21980
rect 16156 21924 16212 31948
rect 16492 32004 16548 32014
rect 16492 31218 16548 31948
rect 16604 31556 16660 32510
rect 17276 32004 17332 33070
rect 17724 33124 17780 33134
rect 17724 32786 17780 33068
rect 17724 32734 17726 32786
rect 17778 32734 17780 32786
rect 17724 32722 17780 32734
rect 17276 31938 17332 31948
rect 17724 32564 17780 32574
rect 17724 31890 17780 32508
rect 18060 32564 18116 32574
rect 18060 32470 18116 32508
rect 17724 31838 17726 31890
rect 17778 31838 17780 31890
rect 17724 31826 17780 31838
rect 18060 32004 18116 32014
rect 18060 31778 18116 31948
rect 18060 31726 18062 31778
rect 18114 31726 18116 31778
rect 18060 31714 18116 31726
rect 16604 31490 16660 31500
rect 17948 31556 18004 31566
rect 16492 31166 16494 31218
rect 16546 31166 16548 31218
rect 16492 31154 16548 31166
rect 16940 30882 16996 30894
rect 17724 30884 17780 30894
rect 16940 30830 16942 30882
rect 16994 30830 16996 30882
rect 16268 29988 16324 29998
rect 16268 29986 16436 29988
rect 16268 29934 16270 29986
rect 16322 29934 16436 29986
rect 16268 29932 16436 29934
rect 16268 29922 16324 29932
rect 16268 29428 16324 29438
rect 16268 29334 16324 29372
rect 16380 29204 16436 29932
rect 16828 29986 16884 29998
rect 16828 29934 16830 29986
rect 16882 29934 16884 29986
rect 16380 29138 16436 29148
rect 16492 29540 16548 29550
rect 16268 28642 16324 28654
rect 16268 28590 16270 28642
rect 16322 28590 16324 28642
rect 16268 28084 16324 28590
rect 16268 28018 16324 28028
rect 16492 27524 16548 29484
rect 16828 29540 16884 29934
rect 16828 29446 16884 29484
rect 16940 28868 16996 30830
rect 17388 30882 17780 30884
rect 17388 30830 17726 30882
rect 17778 30830 17780 30882
rect 17388 30828 17780 30830
rect 17276 29988 17332 29998
rect 17276 29894 17332 29932
rect 16940 28802 16996 28812
rect 17276 29428 17332 29438
rect 16828 28642 16884 28654
rect 16828 28590 16830 28642
rect 16882 28590 16884 28642
rect 16716 27970 16772 27982
rect 16716 27918 16718 27970
rect 16770 27918 16772 27970
rect 16268 27468 16548 27524
rect 16604 27858 16660 27870
rect 16604 27806 16606 27858
rect 16658 27806 16660 27858
rect 16268 27298 16324 27468
rect 16268 27246 16270 27298
rect 16322 27246 16324 27298
rect 16268 27234 16324 27246
rect 16492 27300 16548 27310
rect 16492 26404 16548 27244
rect 16604 27188 16660 27806
rect 16716 27860 16772 27918
rect 16716 27794 16772 27804
rect 16604 27122 16660 27132
rect 16716 27300 16772 27310
rect 16716 27074 16772 27244
rect 16828 27186 16884 28590
rect 17276 28642 17332 29372
rect 17276 28590 17278 28642
rect 17330 28590 17332 28642
rect 17276 28578 17332 28590
rect 16940 28084 16996 28094
rect 16940 27990 16996 28028
rect 16828 27134 16830 27186
rect 16882 27134 16884 27186
rect 16828 27122 16884 27134
rect 17052 27860 17108 27870
rect 16716 27022 16718 27074
rect 16770 27022 16772 27074
rect 16716 27010 16772 27022
rect 16940 26962 16996 26974
rect 16940 26910 16942 26962
rect 16994 26910 16996 26962
rect 16940 26908 16996 26910
rect 16604 26852 16660 26862
rect 16604 26758 16660 26796
rect 16716 26852 16996 26908
rect 16716 26516 16772 26852
rect 16268 26290 16324 26302
rect 16268 26238 16270 26290
rect 16322 26238 16324 26290
rect 16268 25620 16324 26238
rect 16268 25554 16324 25564
rect 16380 25284 16436 25294
rect 16492 25284 16548 26348
rect 16380 25282 16548 25284
rect 16380 25230 16382 25282
rect 16434 25230 16548 25282
rect 16380 25228 16548 25230
rect 16380 25218 16436 25228
rect 16380 24948 16436 24958
rect 16380 24162 16436 24892
rect 16380 24110 16382 24162
rect 16434 24110 16436 24162
rect 16380 24098 16436 24110
rect 16492 24610 16548 25228
rect 16492 24558 16494 24610
rect 16546 24558 16548 24610
rect 16492 23940 16548 24558
rect 16604 26460 16772 26516
rect 16828 26516 16884 26526
rect 17052 26516 17108 27804
rect 17164 27748 17220 27758
rect 17164 27074 17220 27692
rect 17164 27022 17166 27074
rect 17218 27022 17220 27074
rect 17164 26740 17220 27022
rect 17388 26908 17444 30828
rect 17724 30818 17780 30828
rect 17724 30324 17780 30334
rect 17724 28308 17780 30268
rect 17724 28242 17780 28252
rect 17836 29428 17892 29438
rect 17724 27746 17780 27758
rect 17724 27694 17726 27746
rect 17778 27694 17780 27746
rect 17724 27636 17780 27694
rect 17724 27570 17780 27580
rect 17836 27188 17892 29372
rect 17948 28866 18004 31500
rect 18060 29988 18116 29998
rect 18060 29650 18116 29932
rect 18060 29598 18062 29650
rect 18114 29598 18116 29650
rect 18060 29586 18116 29598
rect 17948 28814 17950 28866
rect 18002 28814 18004 28866
rect 17948 28802 18004 28814
rect 18172 28756 18228 28766
rect 18172 28642 18228 28700
rect 18172 28590 18174 28642
rect 18226 28590 18228 28642
rect 18172 28578 18228 28590
rect 18060 28420 18116 28430
rect 18060 27524 18116 28364
rect 18172 27972 18228 27982
rect 18172 27878 18228 27916
rect 18060 27468 18228 27524
rect 17948 27188 18004 27198
rect 18172 27188 18228 27468
rect 17836 27186 18116 27188
rect 17836 27134 17950 27186
rect 18002 27134 18116 27186
rect 17836 27132 18116 27134
rect 17948 27122 18004 27132
rect 17164 26674 17220 26684
rect 17276 26852 17444 26908
rect 17724 27076 17780 27086
rect 16828 26514 17108 26516
rect 16828 26462 16830 26514
rect 16882 26462 17108 26514
rect 16828 26460 17108 26462
rect 16604 24050 16660 26460
rect 16828 26450 16884 26460
rect 16716 26290 16772 26302
rect 16940 26292 16996 26302
rect 16716 26238 16718 26290
rect 16770 26238 16772 26290
rect 16716 26068 16772 26238
rect 16716 26002 16772 26012
rect 16828 26290 16996 26292
rect 16828 26238 16942 26290
rect 16994 26238 16996 26290
rect 16828 26236 16996 26238
rect 16604 23998 16606 24050
rect 16658 23998 16660 24050
rect 16604 23986 16660 23998
rect 16716 25732 16772 25742
rect 16380 23938 16548 23940
rect 16380 23886 16494 23938
rect 16546 23886 16548 23938
rect 16380 23884 16548 23886
rect 16156 21868 16324 21924
rect 16156 21698 16212 21710
rect 16156 21646 16158 21698
rect 16210 21646 16212 21698
rect 16156 21588 16212 21646
rect 16156 21522 16212 21532
rect 16044 21298 16100 21308
rect 15596 18564 15652 18574
rect 15596 18470 15652 18508
rect 15708 18562 15764 18620
rect 15708 18510 15710 18562
rect 15762 18510 15764 18562
rect 15708 18498 15764 18510
rect 15820 19796 15876 19806
rect 15820 18340 15876 19740
rect 15932 19460 15988 19852
rect 15932 19394 15988 19404
rect 16044 20132 16212 20188
rect 16044 19124 16100 20132
rect 16156 20130 16212 20132
rect 16156 20078 16158 20130
rect 16210 20078 16212 20130
rect 16156 20066 16212 20078
rect 16156 19908 16212 19918
rect 16156 19346 16212 19852
rect 16156 19294 16158 19346
rect 16210 19294 16212 19346
rect 16156 19282 16212 19294
rect 16044 19058 16100 19068
rect 16044 18900 16100 18910
rect 15932 18676 15988 18686
rect 15932 18562 15988 18620
rect 15932 18510 15934 18562
rect 15986 18510 15988 18562
rect 15932 18498 15988 18510
rect 15484 17726 15486 17778
rect 15538 17726 15540 17778
rect 15484 17714 15540 17726
rect 15596 18284 15876 18340
rect 15372 17054 15374 17106
rect 15426 17054 15428 17106
rect 15372 17042 15428 17054
rect 15484 16996 15540 17006
rect 15372 16212 15428 16222
rect 15260 16210 15428 16212
rect 15260 16158 15374 16210
rect 15426 16158 15428 16210
rect 15260 16156 15428 16158
rect 15372 16146 15428 16156
rect 15148 15540 15204 15550
rect 15036 15316 15092 15326
rect 14924 15314 15092 15316
rect 14924 15262 15038 15314
rect 15090 15262 15092 15314
rect 14924 15260 15092 15262
rect 14252 14914 14308 14924
rect 14364 15148 14644 15204
rect 15036 15204 15092 15260
rect 13916 12562 13972 12572
rect 14028 13916 14196 13972
rect 14028 12402 14084 13916
rect 14028 12350 14030 12402
rect 14082 12350 14084 12402
rect 14028 12338 14084 12350
rect 14140 13746 14196 13758
rect 14140 13694 14142 13746
rect 14194 13694 14196 13746
rect 13804 11506 13860 11518
rect 13804 11454 13806 11506
rect 13858 11454 13860 11506
rect 13804 11396 13860 11454
rect 13804 11330 13860 11340
rect 14140 11284 14196 13694
rect 14252 13748 14308 13758
rect 14252 12850 14308 13692
rect 14252 12798 14254 12850
rect 14306 12798 14308 12850
rect 14252 12628 14308 12798
rect 14252 12562 14308 12572
rect 14364 12404 14420 15148
rect 15036 15138 15092 15148
rect 14476 14418 14532 14430
rect 14476 14366 14478 14418
rect 14530 14366 14532 14418
rect 14476 14196 14532 14366
rect 14476 13748 14532 14140
rect 14924 14420 14980 14430
rect 14700 13972 14756 13982
rect 14700 13878 14756 13916
rect 14476 13682 14532 13692
rect 14588 13636 14644 13646
rect 14588 12850 14644 13580
rect 14588 12798 14590 12850
rect 14642 12798 14644 12850
rect 14588 12786 14644 12798
rect 14140 11218 14196 11228
rect 14252 12348 14420 12404
rect 14924 12628 14980 14364
rect 15148 13972 15204 15484
rect 15148 13906 15204 13916
rect 15260 14868 15316 14878
rect 15148 13748 15204 13758
rect 14252 11506 14308 12348
rect 14252 11454 14254 11506
rect 14306 11454 14308 11506
rect 13916 10498 13972 10510
rect 13916 10446 13918 10498
rect 13970 10446 13972 10498
rect 13916 10276 13972 10446
rect 13916 10210 13972 10220
rect 14252 10052 14308 11454
rect 14364 12178 14420 12190
rect 14364 12126 14366 12178
rect 14418 12126 14420 12178
rect 14364 11172 14420 12126
rect 14700 11394 14756 11406
rect 14700 11342 14702 11394
rect 14754 11342 14756 11394
rect 14364 11106 14420 11116
rect 14476 11284 14532 11294
rect 14252 9986 14308 9996
rect 14140 9940 14196 9950
rect 14140 9846 14196 9884
rect 13580 9436 13748 9492
rect 13804 9826 13860 9838
rect 13804 9774 13806 9826
rect 13858 9774 13860 9826
rect 13580 8372 13636 9436
rect 13692 9268 13748 9278
rect 13692 9174 13748 9212
rect 13580 8306 13636 8316
rect 13580 8148 13636 8158
rect 13804 8148 13860 9774
rect 14028 9828 14084 9838
rect 13916 9714 13972 9726
rect 13916 9662 13918 9714
rect 13970 9662 13972 9714
rect 13916 9044 13972 9662
rect 14028 9154 14084 9772
rect 14364 9828 14420 9838
rect 14364 9734 14420 9772
rect 14476 9268 14532 11228
rect 14700 10836 14756 11342
rect 14588 10722 14644 10734
rect 14588 10670 14590 10722
rect 14642 10670 14644 10722
rect 14700 10704 14756 10780
rect 14812 11172 14868 11182
rect 14812 10722 14868 11116
rect 14588 10612 14644 10670
rect 14588 10546 14644 10556
rect 14812 10670 14814 10722
rect 14866 10670 14868 10722
rect 14812 10612 14868 10670
rect 14812 10546 14868 10556
rect 14924 10388 14980 12572
rect 15036 13188 15092 13198
rect 15036 13074 15092 13132
rect 15036 13022 15038 13074
rect 15090 13022 15092 13074
rect 15036 12180 15092 13022
rect 15148 12852 15204 13692
rect 15260 13746 15316 14812
rect 15260 13694 15262 13746
rect 15314 13694 15316 13746
rect 15260 13636 15316 13694
rect 15484 13748 15540 16940
rect 15596 14642 15652 18284
rect 15596 14590 15598 14642
rect 15650 14590 15652 14642
rect 15596 14578 15652 14590
rect 15708 17892 15764 17902
rect 15708 13972 15764 17836
rect 16044 17332 16100 18844
rect 16156 18338 16212 18350
rect 16156 18286 16158 18338
rect 16210 18286 16212 18338
rect 16156 17666 16212 18286
rect 16268 17778 16324 21868
rect 16380 21476 16436 23884
rect 16492 23874 16548 23884
rect 16716 23380 16772 25676
rect 16828 23716 16884 26236
rect 16940 26226 16996 26236
rect 16940 25620 16996 25630
rect 16940 25526 16996 25564
rect 17052 25284 17108 25294
rect 16940 24948 16996 24958
rect 17052 24948 17108 25228
rect 16940 24946 17108 24948
rect 16940 24894 16942 24946
rect 16994 24894 17108 24946
rect 16940 24892 17108 24894
rect 16940 24882 16996 24892
rect 16940 24164 16996 24174
rect 16940 24070 16996 24108
rect 17276 24164 17332 26852
rect 17612 26292 17668 26302
rect 17500 26236 17612 26292
rect 17500 25394 17556 26236
rect 17612 26198 17668 26236
rect 17612 25620 17668 25630
rect 17724 25620 17780 27020
rect 17836 26740 17892 26750
rect 17836 26514 17892 26684
rect 17836 26462 17838 26514
rect 17890 26462 17892 26514
rect 17836 26450 17892 26462
rect 17948 26290 18004 26302
rect 17948 26238 17950 26290
rect 18002 26238 18004 26290
rect 17948 25844 18004 26238
rect 17948 25778 18004 25788
rect 17612 25618 17780 25620
rect 17612 25566 17614 25618
rect 17666 25566 17780 25618
rect 17612 25564 17780 25566
rect 17612 25554 17668 25564
rect 17500 25342 17502 25394
rect 17554 25342 17556 25394
rect 17500 25330 17556 25342
rect 17724 25396 17780 25406
rect 17724 25302 17780 25340
rect 18060 25284 18116 27132
rect 18060 25218 18116 25228
rect 18172 25060 18228 27132
rect 17948 25004 18228 25060
rect 17836 24724 17892 24734
rect 17276 24098 17332 24108
rect 17724 24722 17892 24724
rect 17724 24670 17838 24722
rect 17890 24670 17892 24722
rect 17724 24668 17892 24670
rect 17052 24052 17108 24062
rect 17108 23996 17220 24052
rect 17052 23986 17108 23996
rect 17164 23938 17220 23996
rect 17164 23886 17166 23938
rect 17218 23886 17220 23938
rect 17164 23874 17220 23886
rect 17724 23828 17780 24668
rect 17836 24658 17892 24668
rect 17724 23762 17780 23772
rect 17836 23826 17892 23838
rect 17836 23774 17838 23826
rect 17890 23774 17892 23826
rect 17836 23716 17892 23774
rect 16828 23660 17668 23716
rect 17612 23380 17668 23660
rect 17836 23650 17892 23660
rect 17836 23380 17892 23390
rect 17612 23378 17892 23380
rect 17612 23326 17838 23378
rect 17890 23326 17892 23378
rect 17612 23324 17892 23326
rect 16716 23314 16772 23324
rect 17836 23314 17892 23324
rect 16716 23156 16772 23166
rect 16492 23044 16548 23082
rect 16492 22978 16548 22988
rect 16492 22820 16548 22830
rect 16492 21588 16548 22764
rect 16604 22708 16660 22718
rect 16604 22370 16660 22652
rect 16604 22318 16606 22370
rect 16658 22318 16660 22370
rect 16604 22306 16660 22318
rect 16716 21812 16772 23100
rect 17724 23154 17780 23166
rect 17724 23102 17726 23154
rect 17778 23102 17780 23154
rect 16940 23042 16996 23054
rect 16940 22990 16942 23042
rect 16994 22990 16996 23042
rect 16940 22932 16996 22990
rect 17724 23044 17780 23102
rect 17724 22978 17780 22988
rect 16940 22866 16996 22876
rect 17612 22932 17668 22942
rect 17276 22708 17332 22718
rect 16940 22596 16996 22606
rect 16940 22370 16996 22540
rect 16940 22318 16942 22370
rect 16994 22318 16996 22370
rect 16940 22306 16996 22318
rect 16828 22146 16884 22158
rect 16828 22094 16830 22146
rect 16882 22094 16884 22146
rect 16828 22036 16884 22094
rect 16828 21970 16884 21980
rect 16828 21812 16884 21822
rect 16716 21810 16884 21812
rect 16716 21758 16830 21810
rect 16882 21758 16884 21810
rect 16716 21756 16884 21758
rect 16716 21588 16772 21598
rect 16492 21586 16772 21588
rect 16492 21534 16718 21586
rect 16770 21534 16772 21586
rect 16492 21532 16772 21534
rect 16380 21420 16660 21476
rect 16492 20916 16548 20926
rect 16492 20822 16548 20860
rect 16380 20578 16436 20590
rect 16380 20526 16382 20578
rect 16434 20526 16436 20578
rect 16380 17892 16436 20526
rect 16604 20578 16660 21420
rect 16604 20526 16606 20578
rect 16658 20526 16660 20578
rect 16604 19906 16660 20526
rect 16604 19854 16606 19906
rect 16658 19854 16660 19906
rect 16604 19796 16660 19854
rect 16716 19908 16772 21532
rect 16716 19842 16772 19852
rect 16604 19730 16660 19740
rect 16828 19572 16884 21756
rect 17052 21700 17108 21710
rect 17052 21606 17108 21644
rect 16940 21588 16996 21598
rect 16940 20802 16996 21532
rect 16940 20750 16942 20802
rect 16994 20750 16996 20802
rect 16940 20738 16996 20750
rect 16604 19516 16884 19572
rect 17164 19796 17220 19806
rect 16604 19346 16660 19516
rect 16604 19294 16606 19346
rect 16658 19294 16660 19346
rect 16604 19282 16660 19294
rect 16380 17826 16436 17836
rect 16604 19012 16660 19022
rect 16604 18564 16660 18956
rect 16268 17726 16270 17778
rect 16322 17726 16324 17778
rect 16268 17714 16324 17726
rect 16156 17614 16158 17666
rect 16210 17614 16212 17666
rect 16156 17602 16212 17614
rect 16492 17554 16548 17566
rect 16492 17502 16494 17554
rect 16546 17502 16548 17554
rect 16044 17276 16436 17332
rect 16156 16884 16212 16894
rect 16044 16772 16100 16782
rect 16044 16678 16100 16716
rect 16156 16436 16212 16828
rect 16044 16380 16212 16436
rect 16268 16436 16324 16446
rect 16380 16436 16436 17276
rect 16492 16660 16548 17502
rect 16604 17106 16660 18508
rect 16716 18452 16772 19516
rect 17164 19346 17220 19740
rect 17164 19294 17166 19346
rect 17218 19294 17220 19346
rect 17164 19282 17220 19294
rect 16716 18386 16772 18396
rect 17164 18452 17220 18462
rect 17052 18338 17108 18350
rect 17052 18286 17054 18338
rect 17106 18286 17108 18338
rect 17052 18228 17108 18286
rect 17052 18162 17108 18172
rect 17052 17892 17108 17902
rect 16604 17054 16606 17106
rect 16658 17054 16660 17106
rect 16604 17042 16660 17054
rect 16940 17108 16996 17118
rect 16492 16594 16548 16604
rect 16380 16380 16548 16436
rect 15820 16324 15876 16334
rect 15820 16098 15876 16268
rect 15820 16046 15822 16098
rect 15874 16046 15876 16098
rect 15820 16034 15876 16046
rect 16044 16098 16100 16380
rect 16044 16046 16046 16098
rect 16098 16046 16100 16098
rect 16044 15652 16100 16046
rect 16044 15586 16100 15596
rect 16156 16212 16212 16222
rect 16156 15538 16212 16156
rect 16268 15986 16324 16380
rect 16268 15934 16270 15986
rect 16322 15934 16324 15986
rect 16268 15922 16324 15934
rect 16380 15988 16436 15998
rect 16380 15894 16436 15932
rect 16492 15876 16548 16380
rect 16492 15820 16772 15876
rect 16156 15486 16158 15538
rect 16210 15486 16212 15538
rect 16156 15474 16212 15486
rect 16380 15764 16436 15774
rect 16044 15428 16100 15438
rect 16044 15334 16100 15372
rect 16380 15426 16436 15708
rect 16380 15374 16382 15426
rect 16434 15374 16436 15426
rect 16380 15362 16436 15374
rect 16492 15540 16548 15550
rect 15932 15314 15988 15326
rect 15932 15262 15934 15314
rect 15986 15262 15988 15314
rect 15932 15092 15988 15262
rect 15932 14308 15988 15036
rect 16268 15316 16324 15326
rect 16044 14420 16100 14430
rect 16044 14326 16100 14364
rect 16268 14308 16324 15260
rect 16380 14308 16436 14318
rect 16268 14306 16436 14308
rect 16268 14254 16382 14306
rect 16434 14254 16436 14306
rect 16268 14252 16436 14254
rect 15932 14242 15988 14252
rect 15708 13906 15764 13916
rect 16380 13972 16436 14252
rect 16380 13906 16436 13916
rect 16492 13970 16548 15484
rect 16492 13918 16494 13970
rect 16546 13918 16548 13970
rect 16492 13906 16548 13918
rect 15484 13682 15540 13692
rect 15708 13748 15764 13758
rect 15260 13188 15316 13580
rect 15596 13636 15652 13646
rect 15260 13122 15316 13132
rect 15484 13524 15540 13534
rect 15596 13524 15652 13580
rect 15484 13522 15652 13524
rect 15484 13470 15486 13522
rect 15538 13470 15652 13522
rect 15484 13468 15652 13470
rect 15484 12964 15540 13468
rect 15708 13188 15764 13692
rect 15820 13748 15876 13758
rect 16380 13748 16436 13758
rect 16604 13748 16660 13758
rect 15820 13746 16436 13748
rect 15820 13694 15822 13746
rect 15874 13694 16382 13746
rect 16434 13694 16436 13746
rect 15820 13692 16436 13694
rect 15820 13682 15876 13692
rect 16380 13682 16436 13692
rect 16492 13746 16660 13748
rect 16492 13694 16606 13746
rect 16658 13694 16660 13746
rect 16492 13692 16660 13694
rect 15708 13132 15988 13188
rect 15484 12908 15876 12964
rect 15148 12796 15540 12852
rect 15148 12404 15204 12414
rect 15148 12310 15204 12348
rect 15036 12114 15092 12124
rect 15260 11732 15316 11742
rect 15260 10834 15316 11676
rect 15260 10782 15262 10834
rect 15314 10782 15316 10834
rect 15260 10770 15316 10782
rect 15484 11172 15540 12796
rect 15596 12738 15652 12750
rect 15596 12686 15598 12738
rect 15650 12686 15652 12738
rect 15596 11956 15652 12686
rect 15708 12404 15764 12414
rect 15708 12310 15764 12348
rect 15596 11890 15652 11900
rect 15820 11284 15876 12908
rect 15932 11506 15988 13132
rect 16492 13186 16548 13692
rect 16604 13682 16660 13692
rect 16492 13134 16494 13186
rect 16546 13134 16548 13186
rect 16492 13122 16548 13134
rect 16044 12964 16100 12974
rect 16044 12870 16100 12908
rect 16604 12962 16660 12974
rect 16604 12910 16606 12962
rect 16658 12910 16660 12962
rect 16604 12852 16660 12910
rect 16380 12796 16660 12852
rect 16156 12740 16212 12750
rect 16044 12516 16100 12526
rect 16044 12402 16100 12460
rect 16044 12350 16046 12402
rect 16098 12350 16100 12402
rect 16044 12180 16100 12350
rect 16044 12114 16100 12124
rect 15932 11454 15934 11506
rect 15986 11454 15988 11506
rect 15932 11442 15988 11454
rect 15820 11228 15988 11284
rect 14812 10332 14980 10388
rect 14028 9102 14030 9154
rect 14082 9102 14084 9154
rect 14028 9090 14084 9102
rect 14140 9212 14532 9268
rect 14700 9828 14756 9838
rect 14700 9266 14756 9772
rect 14812 9604 14868 10332
rect 14924 10052 14980 10062
rect 14980 9996 15428 10052
rect 14924 9986 14980 9996
rect 14924 9828 14980 9838
rect 14924 9734 14980 9772
rect 15260 9828 15316 9838
rect 15260 9734 15316 9772
rect 15372 9714 15428 9996
rect 15372 9662 15374 9714
rect 15426 9662 15428 9714
rect 14812 9548 15092 9604
rect 14700 9214 14702 9266
rect 14754 9214 14756 9266
rect 13916 8978 13972 8988
rect 14028 8148 14084 8158
rect 13804 8146 14084 8148
rect 13804 8094 14030 8146
rect 14082 8094 14084 8146
rect 13804 8092 14084 8094
rect 13580 8036 13636 8092
rect 13692 8036 13748 8046
rect 13580 8034 13748 8036
rect 13580 7982 13694 8034
rect 13746 7982 13748 8034
rect 13580 7980 13748 7982
rect 13580 7698 13636 7980
rect 13692 7970 13748 7980
rect 14028 8036 14084 8092
rect 14028 7970 14084 7980
rect 13580 7646 13582 7698
rect 13634 7646 13636 7698
rect 13580 7634 13636 7646
rect 13804 7924 13860 7934
rect 13692 7474 13748 7486
rect 13692 7422 13694 7474
rect 13746 7422 13748 7474
rect 13692 7364 13748 7422
rect 13580 6692 13636 6702
rect 13580 6598 13636 6636
rect 13692 6580 13748 7308
rect 13692 6514 13748 6524
rect 13692 6132 13748 6142
rect 13804 6132 13860 7868
rect 14028 6580 14084 6590
rect 14028 6486 14084 6524
rect 13692 6130 13860 6132
rect 13692 6078 13694 6130
rect 13746 6078 13860 6130
rect 13692 6076 13860 6078
rect 13916 6466 13972 6478
rect 13916 6414 13918 6466
rect 13970 6414 13972 6466
rect 13692 6066 13748 6076
rect 13468 5630 13470 5682
rect 13522 5630 13524 5682
rect 13468 5618 13524 5630
rect 12908 5572 12964 5582
rect 12908 5234 12964 5516
rect 12908 5182 12910 5234
rect 12962 5182 12964 5234
rect 12908 5170 12964 5182
rect 13020 4564 13076 4574
rect 13020 4470 13076 4508
rect 13804 4452 13860 4462
rect 13804 4358 13860 4396
rect 12684 4274 12740 4284
rect 11676 4226 11732 4238
rect 11676 4174 11678 4226
rect 11730 4174 11732 4226
rect 11676 4114 11732 4174
rect 11676 4062 11678 4114
rect 11730 4062 11732 4114
rect 11676 4050 11732 4062
rect 13580 3668 13636 3678
rect 13580 3574 13636 3612
rect 11340 3500 11620 3556
rect 12796 3556 12852 3566
rect 11340 3332 11396 3500
rect 12796 3462 12852 3500
rect 11676 3442 11732 3454
rect 11676 3390 11678 3442
rect 11730 3390 11732 3442
rect 11676 3388 11732 3390
rect 11340 3266 11396 3276
rect 11452 3332 11732 3388
rect 8316 1362 8372 1372
rect 11452 800 11508 3332
rect 13916 3220 13972 6414
rect 14028 6244 14084 6254
rect 14028 5234 14084 6188
rect 14140 6130 14196 9212
rect 14700 8146 14756 9214
rect 14812 9380 14868 9390
rect 14812 9266 14868 9324
rect 14812 9214 14814 9266
rect 14866 9214 14868 9266
rect 14812 9202 14868 9214
rect 14924 9156 14980 9166
rect 14924 9062 14980 9100
rect 14700 8094 14702 8146
rect 14754 8094 14756 8146
rect 14700 8082 14756 8094
rect 14812 8932 14868 8942
rect 15036 8932 15092 9548
rect 14252 7700 14308 7710
rect 14252 7606 14308 7644
rect 14588 7476 14644 7486
rect 14588 7382 14644 7420
rect 14140 6078 14142 6130
rect 14194 6078 14196 6130
rect 14140 5460 14196 6078
rect 14140 5394 14196 5404
rect 14252 6580 14308 6590
rect 14252 5572 14308 6524
rect 14812 6020 14868 8876
rect 14924 8876 15092 8932
rect 15260 9044 15316 9054
rect 14924 6244 14980 8876
rect 15036 8034 15092 8046
rect 15036 7982 15038 8034
rect 15090 7982 15092 8034
rect 15036 7700 15092 7982
rect 15148 7700 15204 7710
rect 15036 7698 15204 7700
rect 15036 7646 15150 7698
rect 15202 7646 15204 7698
rect 15036 7644 15204 7646
rect 15036 7476 15092 7644
rect 15148 7634 15204 7644
rect 15036 6914 15092 7420
rect 15036 6862 15038 6914
rect 15090 6862 15092 6914
rect 15036 6850 15092 6862
rect 15148 6580 15204 6590
rect 15148 6486 15204 6524
rect 14924 6178 14980 6188
rect 15148 6132 15204 6142
rect 15148 6038 15204 6076
rect 14812 5964 14980 6020
rect 14028 5182 14030 5234
rect 14082 5182 14084 5234
rect 14028 5170 14084 5182
rect 14140 4564 14196 4574
rect 14140 4470 14196 4508
rect 14252 3666 14308 5516
rect 14588 5794 14644 5806
rect 14588 5742 14590 5794
rect 14642 5742 14644 5794
rect 14588 5682 14644 5742
rect 14588 5630 14590 5682
rect 14642 5630 14644 5682
rect 14588 4788 14644 5630
rect 14812 5236 14868 5246
rect 14812 5142 14868 5180
rect 14588 4722 14644 4732
rect 14588 4564 14644 4574
rect 14588 4470 14644 4508
rect 14252 3614 14254 3666
rect 14306 3614 14308 3666
rect 14252 3602 14308 3614
rect 14700 3668 14756 3678
rect 14924 3668 14980 5964
rect 14700 3666 14980 3668
rect 14700 3614 14702 3666
rect 14754 3614 14980 3666
rect 14700 3612 14980 3614
rect 15148 4564 15204 4574
rect 15148 4116 15204 4508
rect 15148 3666 15204 4060
rect 15148 3614 15150 3666
rect 15202 3614 15204 3666
rect 14700 3602 14756 3612
rect 15148 3602 15204 3614
rect 15260 3668 15316 8988
rect 15372 5234 15428 9662
rect 15484 6132 15540 11116
rect 15820 10724 15876 10734
rect 15708 10722 15876 10724
rect 15708 10670 15822 10722
rect 15874 10670 15876 10722
rect 15708 10668 15876 10670
rect 15484 6066 15540 6076
rect 15596 10612 15652 10622
rect 15372 5182 15374 5234
rect 15426 5182 15428 5234
rect 15372 5170 15428 5182
rect 15372 4788 15428 4798
rect 15372 4226 15428 4732
rect 15372 4174 15374 4226
rect 15426 4174 15428 4226
rect 15372 4004 15428 4174
rect 15596 4788 15652 10556
rect 15708 8148 15764 10668
rect 15820 10658 15876 10668
rect 15932 10500 15988 11228
rect 15820 10444 15988 10500
rect 16044 10612 16100 10622
rect 15820 9492 15876 10444
rect 16044 10276 16100 10556
rect 16044 10210 16100 10220
rect 16156 10052 16212 12684
rect 16268 12628 16324 12638
rect 16268 10498 16324 12572
rect 16268 10446 16270 10498
rect 16322 10446 16324 10498
rect 16268 10434 16324 10446
rect 16380 11844 16436 12796
rect 16604 12404 16660 12414
rect 16716 12404 16772 15820
rect 16940 15764 16996 17052
rect 17052 17106 17108 17836
rect 17052 17054 17054 17106
rect 17106 17054 17108 17106
rect 17052 17042 17108 17054
rect 17052 16212 17108 16222
rect 17052 16098 17108 16156
rect 17052 16046 17054 16098
rect 17106 16046 17108 16098
rect 17052 16034 17108 16046
rect 16828 15708 16996 15764
rect 16828 13972 16884 15708
rect 17052 15652 17108 15662
rect 16940 15540 16996 15550
rect 17052 15540 17108 15596
rect 16940 15538 17108 15540
rect 16940 15486 16942 15538
rect 16994 15486 17108 15538
rect 16940 15484 17108 15486
rect 16940 15474 16996 15484
rect 17052 14754 17108 14766
rect 17052 14702 17054 14754
rect 17106 14702 17108 14754
rect 17052 14642 17108 14702
rect 17052 14590 17054 14642
rect 17106 14590 17108 14642
rect 17052 14578 17108 14590
rect 17164 14532 17220 18396
rect 17276 17778 17332 22652
rect 17500 21812 17556 21822
rect 17500 21364 17556 21756
rect 17500 21298 17556 21308
rect 17612 20692 17668 22876
rect 17836 22148 17892 22158
rect 17836 22054 17892 22092
rect 17948 21924 18004 25004
rect 18172 24834 18228 24846
rect 18172 24782 18174 24834
rect 18226 24782 18228 24834
rect 18172 24724 18228 24782
rect 18172 24388 18228 24668
rect 18172 24322 18228 24332
rect 18284 24164 18340 35086
rect 18396 35476 18452 36204
rect 18396 35026 18452 35420
rect 18396 34974 18398 35026
rect 18450 34974 18452 35026
rect 18396 34962 18452 34974
rect 18508 32676 18564 37996
rect 18620 37826 18676 37838
rect 18620 37774 18622 37826
rect 18674 37774 18676 37826
rect 18620 37492 18676 37774
rect 18620 37426 18676 37436
rect 18732 37380 18788 38108
rect 18956 38052 19012 38062
rect 18844 37940 18900 37950
rect 18956 37940 19012 37996
rect 18844 37938 19012 37940
rect 18844 37886 18846 37938
rect 18898 37886 19012 37938
rect 18844 37884 19012 37886
rect 18844 37874 18900 37884
rect 18620 37156 18676 37166
rect 18620 37042 18676 37100
rect 18620 36990 18622 37042
rect 18674 36990 18676 37042
rect 18620 34580 18676 36990
rect 18732 36594 18788 37324
rect 18732 36542 18734 36594
rect 18786 36542 18788 36594
rect 18732 36530 18788 36542
rect 18844 35586 18900 35598
rect 18844 35534 18846 35586
rect 18898 35534 18900 35586
rect 18844 35476 18900 35534
rect 18956 35588 19012 37884
rect 19068 37268 19124 37278
rect 19068 37174 19124 37212
rect 18956 35522 19012 35532
rect 19180 36258 19236 36270
rect 19180 36206 19182 36258
rect 19234 36206 19236 36258
rect 18844 35364 18900 35420
rect 18844 35308 19012 35364
rect 18844 34802 18900 34814
rect 18844 34750 18846 34802
rect 18898 34750 18900 34802
rect 18620 34524 18788 34580
rect 18620 34130 18676 34142
rect 18620 34078 18622 34130
rect 18674 34078 18676 34130
rect 18620 33124 18676 34078
rect 18620 33058 18676 33068
rect 18620 32676 18676 32686
rect 18508 32674 18676 32676
rect 18508 32622 18622 32674
rect 18674 32622 18676 32674
rect 18508 32620 18676 32622
rect 18620 32610 18676 32620
rect 18732 32452 18788 34524
rect 18844 34356 18900 34750
rect 18844 34290 18900 34300
rect 18620 32396 18788 32452
rect 18508 31666 18564 31678
rect 18508 31614 18510 31666
rect 18562 31614 18564 31666
rect 18508 31556 18564 31614
rect 18508 31490 18564 31500
rect 18396 30882 18452 30894
rect 18396 30830 18398 30882
rect 18450 30830 18452 30882
rect 18396 30324 18452 30830
rect 18396 30258 18452 30268
rect 18508 30770 18564 30782
rect 18508 30718 18510 30770
rect 18562 30718 18564 30770
rect 18396 29988 18452 29998
rect 18396 29894 18452 29932
rect 18508 28868 18564 30718
rect 18620 29876 18676 32396
rect 18844 30882 18900 30894
rect 18844 30830 18846 30882
rect 18898 30830 18900 30882
rect 18844 30770 18900 30830
rect 18844 30718 18846 30770
rect 18898 30718 18900 30770
rect 18844 30706 18900 30718
rect 18956 30324 19012 35308
rect 19180 34356 19236 36206
rect 19292 35588 19348 35598
rect 19292 35494 19348 35532
rect 19180 34290 19236 34300
rect 19292 34692 19348 34702
rect 19292 33796 19348 34636
rect 19292 33730 19348 33740
rect 19180 33124 19236 33134
rect 19180 33030 19236 33068
rect 19404 32676 19460 39004
rect 20412 38948 20468 38958
rect 20412 38854 20468 38892
rect 19852 38722 19908 38734
rect 19852 38670 19854 38722
rect 19906 38670 19908 38722
rect 19852 38668 19908 38670
rect 19852 38612 20132 38668
rect 19852 38546 19908 38556
rect 19740 38500 19796 38510
rect 19516 38388 19572 38398
rect 19516 38050 19572 38332
rect 19516 37998 19518 38050
rect 19570 37998 19572 38050
rect 19516 37986 19572 37998
rect 19740 38050 19796 38444
rect 19740 37998 19742 38050
rect 19794 37998 19796 38050
rect 19740 37986 19796 37998
rect 20076 37938 20132 38612
rect 20076 37886 20078 37938
rect 20130 37886 20132 37938
rect 19628 37826 19684 37838
rect 19628 37774 19630 37826
rect 19682 37774 19684 37826
rect 19628 37492 19684 37774
rect 20076 37828 20132 37886
rect 20076 37762 20132 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19628 37436 19908 37492
rect 19852 37378 19908 37436
rect 20636 37490 20692 40236
rect 20636 37438 20638 37490
rect 20690 37438 20692 37490
rect 20636 37426 20692 37438
rect 19852 37326 19854 37378
rect 19906 37326 19908 37378
rect 19852 36482 19908 37326
rect 19964 37268 20020 37278
rect 20020 37212 20244 37268
rect 19964 37174 20020 37212
rect 19852 36430 19854 36482
rect 19906 36430 19908 36482
rect 19852 36418 19908 36430
rect 20188 36482 20244 37212
rect 20636 37266 20692 37278
rect 20636 37214 20638 37266
rect 20690 37214 20692 37266
rect 20188 36430 20190 36482
rect 20242 36430 20244 36482
rect 20188 36418 20244 36430
rect 20524 36596 20580 36606
rect 20412 36372 20468 36382
rect 20412 36278 20468 36316
rect 20076 36260 20132 36270
rect 20076 36258 20244 36260
rect 20076 36206 20078 36258
rect 20130 36206 20244 36258
rect 20076 36204 20244 36206
rect 20076 36194 20132 36204
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20188 35924 20244 36204
rect 20076 35868 20244 35924
rect 19852 35698 19908 35710
rect 19852 35646 19854 35698
rect 19906 35646 19908 35698
rect 19852 35026 19908 35646
rect 20076 35698 20132 35868
rect 20412 35812 20468 35822
rect 20524 35812 20580 36540
rect 20412 35810 20580 35812
rect 20412 35758 20414 35810
rect 20466 35758 20580 35810
rect 20412 35756 20580 35758
rect 20412 35746 20468 35756
rect 20076 35646 20078 35698
rect 20130 35646 20132 35698
rect 20076 35634 20132 35646
rect 20300 35474 20356 35486
rect 20300 35422 20302 35474
rect 20354 35422 20356 35474
rect 20300 35364 20356 35422
rect 20300 35298 20356 35308
rect 20412 35140 20468 35150
rect 19852 34974 19854 35026
rect 19906 34974 19908 35026
rect 19852 34962 19908 34974
rect 20300 35028 20356 35038
rect 20412 35028 20468 35084
rect 20300 35026 20468 35028
rect 20300 34974 20302 35026
rect 20354 34974 20468 35026
rect 20300 34972 20468 34974
rect 20300 34962 20356 34972
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19740 34130 19796 34142
rect 19740 34078 19742 34130
rect 19794 34078 19796 34130
rect 19740 33796 19796 34078
rect 19740 33730 19796 33740
rect 20412 34018 20468 34972
rect 20524 34914 20580 34926
rect 20524 34862 20526 34914
rect 20578 34862 20580 34914
rect 20524 34804 20580 34862
rect 20524 34738 20580 34748
rect 20636 34242 20692 37214
rect 20748 36708 20804 41468
rect 20860 40964 20916 40974
rect 20860 40870 20916 40908
rect 20860 40404 20916 40414
rect 20860 39284 20916 40348
rect 20972 40402 21028 40414
rect 20972 40350 20974 40402
rect 21026 40350 21028 40402
rect 20972 39732 21028 40350
rect 20972 39666 21028 39676
rect 21084 39620 21140 39630
rect 20860 39228 21028 39284
rect 20860 38948 20916 38958
rect 20860 38854 20916 38892
rect 20860 38388 20916 38398
rect 20860 38162 20916 38332
rect 20860 38110 20862 38162
rect 20914 38110 20916 38162
rect 20860 37940 20916 38110
rect 20860 37874 20916 37884
rect 20860 37380 20916 37390
rect 20972 37380 21028 39228
rect 21084 39172 21140 39564
rect 21084 39058 21140 39116
rect 21084 39006 21086 39058
rect 21138 39006 21140 39058
rect 21084 38994 21140 39006
rect 21196 38836 21252 43148
rect 21308 42532 21364 42542
rect 21308 42194 21364 42476
rect 21308 42142 21310 42194
rect 21362 42142 21364 42194
rect 21308 42130 21364 42142
rect 21868 41186 21924 41198
rect 21868 41134 21870 41186
rect 21922 41134 21924 41186
rect 21644 41074 21700 41086
rect 21644 41022 21646 41074
rect 21698 41022 21700 41074
rect 21644 40964 21700 41022
rect 21644 40898 21700 40908
rect 21644 40516 21700 40526
rect 21644 40514 21812 40516
rect 21644 40462 21646 40514
rect 21698 40462 21812 40514
rect 21644 40460 21812 40462
rect 21644 40450 21700 40460
rect 21532 40402 21588 40414
rect 21532 40350 21534 40402
rect 21586 40350 21588 40402
rect 20860 37378 21028 37380
rect 20860 37326 20862 37378
rect 20914 37326 21028 37378
rect 20860 37324 21028 37326
rect 21084 38780 21252 38836
rect 21308 39396 21364 39406
rect 20860 37044 20916 37324
rect 20860 36978 20916 36988
rect 20748 36642 20804 36652
rect 20860 35586 20916 35598
rect 20860 35534 20862 35586
rect 20914 35534 20916 35586
rect 20860 35364 20916 35534
rect 20860 35298 20916 35308
rect 20636 34190 20638 34242
rect 20690 34190 20692 34242
rect 20636 34178 20692 34190
rect 21084 34916 21140 38780
rect 21308 38668 21364 39340
rect 21532 39396 21588 40350
rect 21644 40178 21700 40190
rect 21644 40126 21646 40178
rect 21698 40126 21700 40178
rect 21644 39618 21700 40126
rect 21644 39566 21646 39618
rect 21698 39566 21700 39618
rect 21644 39554 21700 39566
rect 21532 39330 21588 39340
rect 21756 39172 21812 40460
rect 21868 40404 21924 41134
rect 22204 40964 22260 40974
rect 22204 40870 22260 40908
rect 21868 40338 21924 40348
rect 22204 40292 22260 40302
rect 21980 40290 22260 40292
rect 21980 40238 22206 40290
rect 22258 40238 22260 40290
rect 21980 40236 22260 40238
rect 21756 39106 21812 39116
rect 21868 40068 21924 40078
rect 21756 38948 21812 38958
rect 21756 38854 21812 38892
rect 21196 38612 21252 38622
rect 21308 38612 21476 38668
rect 21196 38518 21252 38556
rect 21420 36820 21476 38612
rect 21532 37828 21588 37838
rect 21532 37734 21588 37772
rect 21532 37380 21588 37390
rect 21532 37266 21588 37324
rect 21532 37214 21534 37266
rect 21586 37214 21588 37266
rect 21532 37202 21588 37214
rect 21868 37156 21924 40012
rect 21980 39394 22036 40236
rect 22204 40226 22260 40236
rect 22092 39732 22148 39742
rect 22092 39638 22148 39676
rect 21980 39342 21982 39394
rect 22034 39342 22036 39394
rect 21980 38834 22036 39342
rect 22204 39396 22260 39406
rect 22204 39302 22260 39340
rect 21980 38782 21982 38834
rect 22034 38782 22036 38834
rect 21980 38388 22036 38782
rect 22204 38724 22260 38734
rect 22428 38668 22484 43372
rect 22764 41412 22820 43652
rect 22988 43650 23044 43652
rect 22988 43598 22990 43650
rect 23042 43598 23044 43650
rect 22988 42978 23044 43598
rect 23212 43650 23268 43652
rect 23212 43598 23214 43650
rect 23266 43598 23268 43650
rect 23212 43586 23268 43598
rect 23100 43540 23156 43550
rect 23100 43446 23156 43484
rect 22988 42926 22990 42978
rect 23042 42926 23044 42978
rect 22988 42914 23044 42926
rect 23884 43316 23940 43326
rect 23324 42868 23380 42878
rect 23324 42774 23380 42812
rect 22876 42754 22932 42766
rect 22876 42702 22878 42754
rect 22930 42702 22932 42754
rect 22876 42196 22932 42702
rect 22876 42130 22932 42140
rect 23324 42084 23380 42094
rect 23100 41412 23156 41422
rect 22764 41410 23156 41412
rect 22764 41358 23102 41410
rect 23154 41358 23156 41410
rect 22764 41356 23156 41358
rect 23100 41346 23156 41356
rect 22764 41076 22820 41086
rect 22540 41074 22820 41076
rect 22540 41022 22766 41074
rect 22818 41022 22820 41074
rect 22540 41020 22820 41022
rect 22540 39058 22596 41020
rect 22764 41010 22820 41020
rect 22988 40964 23044 40974
rect 22988 40870 23044 40908
rect 23324 40404 23380 42028
rect 23884 40514 23940 43260
rect 23884 40462 23886 40514
rect 23938 40462 23940 40514
rect 23884 40450 23940 40462
rect 24108 42868 24164 42878
rect 24108 42642 24164 42812
rect 24108 42590 24110 42642
rect 24162 42590 24164 42642
rect 23548 40404 23604 40414
rect 23324 40402 23548 40404
rect 23324 40350 23326 40402
rect 23378 40350 23548 40402
rect 23324 40348 23548 40350
rect 23324 40338 23380 40348
rect 22652 40290 22708 40302
rect 22652 40238 22654 40290
rect 22706 40238 22708 40290
rect 22652 39396 22708 40238
rect 22652 39330 22708 39340
rect 22764 40292 22820 40302
rect 22764 39730 22820 40236
rect 22764 39678 22766 39730
rect 22818 39678 22820 39730
rect 22540 39006 22542 39058
rect 22594 39006 22596 39058
rect 22540 38994 22596 39006
rect 22204 38630 22260 38668
rect 21980 38322 22036 38332
rect 22316 38612 22484 38668
rect 22540 38836 22596 38846
rect 22764 38836 22820 39678
rect 23212 39396 23268 39406
rect 23212 39302 23268 39340
rect 22988 38948 23044 38958
rect 22988 38854 23044 38892
rect 22540 38834 22820 38836
rect 22540 38782 22542 38834
rect 22594 38782 22820 38834
rect 22540 38780 22820 38782
rect 22204 38050 22260 38062
rect 22204 37998 22206 38050
rect 22258 37998 22260 38050
rect 22204 37828 22260 37998
rect 21868 37100 22148 37156
rect 21756 37044 21812 37054
rect 21812 36988 22036 37044
rect 21756 36978 21812 36988
rect 21084 34132 21140 34860
rect 21308 36764 21476 36820
rect 21196 34132 21252 34142
rect 21084 34130 21252 34132
rect 21084 34078 21198 34130
rect 21250 34078 21252 34130
rect 21084 34076 21252 34078
rect 21196 34066 21252 34076
rect 20412 33966 20414 34018
rect 20466 33966 20468 34018
rect 19852 33124 19908 33134
rect 19292 32620 19460 32676
rect 19628 33122 19908 33124
rect 19628 33070 19854 33122
rect 19906 33070 19908 33122
rect 19628 33068 19908 33070
rect 20412 33124 20468 33966
rect 21308 33908 21364 36764
rect 21644 36372 21700 36382
rect 21644 36278 21700 36316
rect 21980 36370 22036 36988
rect 21980 36318 21982 36370
rect 22034 36318 22036 36370
rect 21980 36306 22036 36318
rect 21420 35586 21476 35598
rect 21420 35534 21422 35586
rect 21474 35534 21476 35586
rect 21420 34692 21476 35534
rect 21868 35586 21924 35598
rect 21868 35534 21870 35586
rect 21922 35534 21924 35586
rect 21868 35140 21924 35534
rect 21868 35074 21924 35084
rect 21980 34804 22036 34814
rect 21980 34710 22036 34748
rect 21420 34626 21476 34636
rect 21644 34692 21700 34702
rect 21644 34598 21700 34636
rect 21196 33852 21364 33908
rect 21420 34356 21476 34366
rect 20860 33124 20916 33134
rect 20412 33122 21028 33124
rect 20412 33070 20862 33122
rect 20914 33070 21028 33122
rect 20412 33068 21028 33070
rect 19292 30436 19348 32620
rect 19516 32562 19572 32574
rect 19516 32510 19518 32562
rect 19570 32510 19572 32562
rect 19404 32450 19460 32462
rect 19404 32398 19406 32450
rect 19458 32398 19460 32450
rect 19404 31892 19460 32398
rect 19404 31826 19460 31836
rect 19404 31668 19460 31678
rect 19404 31554 19460 31612
rect 19404 31502 19406 31554
rect 19458 31502 19460 31554
rect 19404 31108 19460 31502
rect 19404 30976 19460 31052
rect 19516 30996 19572 32510
rect 19516 30930 19572 30940
rect 19628 32004 19684 33068
rect 19852 33058 19908 33068
rect 20860 33058 20916 33068
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 20636 32676 20692 32686
rect 20636 32582 20692 32620
rect 20860 32676 20916 32686
rect 20524 32564 20580 32574
rect 20524 32470 20580 32508
rect 19628 30772 19684 31948
rect 20188 31892 20244 31902
rect 20860 31892 20916 32620
rect 20972 32340 21028 33068
rect 20972 32284 21140 32340
rect 20188 31798 20244 31836
rect 20636 31890 20916 31892
rect 20636 31838 20862 31890
rect 20914 31838 20916 31890
rect 20636 31836 20916 31838
rect 20076 31668 20132 31678
rect 20076 31574 20132 31612
rect 20300 31554 20356 31566
rect 20300 31502 20302 31554
rect 20354 31502 20356 31554
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19964 31108 20020 31118
rect 19628 30706 19684 30716
rect 19852 30996 19908 31006
rect 19292 30380 19572 30436
rect 18956 30258 19012 30268
rect 18732 30100 18788 30110
rect 19292 30100 19348 30110
rect 18788 30098 19348 30100
rect 18788 30046 19294 30098
rect 19346 30046 19348 30098
rect 18788 30044 19348 30046
rect 18732 30006 18788 30044
rect 19292 30034 19348 30044
rect 18620 29820 18788 29876
rect 18620 29428 18676 29438
rect 18620 29334 18676 29372
rect 18508 28812 18676 28868
rect 18508 28644 18564 28654
rect 18508 28550 18564 28588
rect 18396 28084 18452 28094
rect 18620 28084 18676 28812
rect 18396 25618 18452 28028
rect 18508 28028 18676 28084
rect 18732 28082 18788 29820
rect 19180 29314 19236 29326
rect 19180 29262 19182 29314
rect 19234 29262 19236 29314
rect 18732 28030 18734 28082
rect 18786 28030 18788 28082
rect 18508 27300 18564 28028
rect 18732 28018 18788 28030
rect 18844 28308 18900 28318
rect 18844 28082 18900 28252
rect 18844 28030 18846 28082
rect 18898 28030 18900 28082
rect 18844 28018 18900 28030
rect 19180 28084 19236 29262
rect 19404 28754 19460 28766
rect 19404 28702 19406 28754
rect 19458 28702 19460 28754
rect 19292 28642 19348 28654
rect 19292 28590 19294 28642
rect 19346 28590 19348 28642
rect 19292 28308 19348 28590
rect 19292 28242 19348 28252
rect 19180 28028 19348 28084
rect 18620 27860 18676 27870
rect 18620 27766 18676 27804
rect 19180 27858 19236 27870
rect 19180 27806 19182 27858
rect 19234 27806 19236 27858
rect 19180 27636 19236 27806
rect 19292 27860 19348 28028
rect 19292 27794 19348 27804
rect 19180 27570 19236 27580
rect 18508 27234 18564 27244
rect 18844 27412 18900 27422
rect 18844 27186 18900 27356
rect 18844 27134 18846 27186
rect 18898 27134 18900 27186
rect 18844 27122 18900 27134
rect 18508 27076 18564 27086
rect 18508 26982 18564 27020
rect 19292 26964 19348 27002
rect 19292 26898 19348 26908
rect 18620 26852 18676 26862
rect 18508 26068 18564 26078
rect 18508 25974 18564 26012
rect 18396 25566 18398 25618
rect 18450 25566 18452 25618
rect 18396 25554 18452 25566
rect 18396 24724 18452 24734
rect 18396 24498 18452 24668
rect 18396 24446 18398 24498
rect 18450 24446 18452 24498
rect 18396 24434 18452 24446
rect 18172 24108 18340 24164
rect 18396 24162 18452 24174
rect 18396 24110 18398 24162
rect 18450 24110 18452 24162
rect 18060 23828 18116 23838
rect 18060 23734 18116 23772
rect 18060 23268 18116 23278
rect 18060 22372 18116 23212
rect 18172 23044 18228 24108
rect 18396 24052 18452 24110
rect 18396 23986 18452 23996
rect 18508 24164 18564 24174
rect 18508 23938 18564 24108
rect 18508 23886 18510 23938
rect 18562 23886 18564 23938
rect 18284 23714 18340 23726
rect 18284 23662 18286 23714
rect 18338 23662 18340 23714
rect 18284 23266 18340 23662
rect 18284 23214 18286 23266
rect 18338 23214 18340 23266
rect 18284 23202 18340 23214
rect 18508 23044 18564 23886
rect 18172 22988 18340 23044
rect 18172 22372 18228 22382
rect 18060 22370 18228 22372
rect 18060 22318 18174 22370
rect 18226 22318 18228 22370
rect 18060 22316 18228 22318
rect 18172 22306 18228 22316
rect 17836 21868 18004 21924
rect 17836 21810 17892 21868
rect 17836 21758 17838 21810
rect 17890 21758 17892 21810
rect 17836 21746 17892 21758
rect 18172 21812 18228 21822
rect 17948 21698 18004 21710
rect 17948 21646 17950 21698
rect 18002 21646 18004 21698
rect 17724 21586 17780 21598
rect 17724 21534 17726 21586
rect 17778 21534 17780 21586
rect 17724 20916 17780 21534
rect 17724 20850 17780 20860
rect 17724 20692 17780 20702
rect 17612 20690 17780 20692
rect 17612 20638 17726 20690
rect 17778 20638 17780 20690
rect 17612 20636 17780 20638
rect 17724 20626 17780 20636
rect 17948 20132 18004 21646
rect 18060 21700 18116 21738
rect 18060 21634 18116 21644
rect 18172 21698 18228 21756
rect 18172 21646 18174 21698
rect 18226 21646 18228 21698
rect 18060 21364 18116 21374
rect 18060 20804 18116 21308
rect 18172 21028 18228 21646
rect 18284 21364 18340 22988
rect 18508 22978 18564 22988
rect 18620 22596 18676 26796
rect 19292 26516 19348 26526
rect 19404 26516 19460 28702
rect 19516 28084 19572 30380
rect 19740 30324 19796 30334
rect 19740 30210 19796 30268
rect 19740 30158 19742 30210
rect 19794 30158 19796 30210
rect 19740 30146 19796 30158
rect 19852 29988 19908 30940
rect 19964 30324 20020 31052
rect 19964 30258 20020 30268
rect 20076 30996 20132 31006
rect 20076 30210 20132 30940
rect 20300 30324 20356 31502
rect 20300 30258 20356 30268
rect 20076 30158 20078 30210
rect 20130 30158 20132 30210
rect 20076 30146 20132 30158
rect 20636 30212 20692 31836
rect 20860 31826 20916 31836
rect 20860 30324 20916 30334
rect 20636 30210 20804 30212
rect 20636 30158 20638 30210
rect 20690 30158 20804 30210
rect 20636 30156 20804 30158
rect 20636 30146 20692 30156
rect 19628 29986 19908 29988
rect 19628 29934 19854 29986
rect 19906 29934 19908 29986
rect 19628 29932 19908 29934
rect 19628 29652 19684 29932
rect 19852 29922 19908 29932
rect 20748 29876 20804 30156
rect 20860 30098 20916 30268
rect 20860 30046 20862 30098
rect 20914 30046 20916 30098
rect 20860 30034 20916 30046
rect 19836 29820 20100 29830
rect 20748 29820 21028 29876
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 20972 29652 21028 29820
rect 19628 29596 19796 29652
rect 19628 29428 19684 29438
rect 19628 29334 19684 29372
rect 19740 28530 19796 29596
rect 19740 28478 19742 28530
rect 19794 28478 19796 28530
rect 19740 28466 19796 28478
rect 20188 29538 20244 29550
rect 20188 29486 20190 29538
rect 20242 29486 20244 29538
rect 20972 29520 21028 29596
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19516 28028 20132 28084
rect 19740 27860 19796 27870
rect 19740 27766 19796 27804
rect 20076 27186 20132 28028
rect 20188 27412 20244 29486
rect 20412 29428 20468 29438
rect 20412 29334 20468 29372
rect 20748 29428 20804 29438
rect 20524 28420 20580 28430
rect 20188 27346 20244 27356
rect 20300 28418 20580 28420
rect 20300 28366 20526 28418
rect 20578 28366 20580 28418
rect 20300 28364 20580 28366
rect 20300 27858 20356 28364
rect 20524 28354 20580 28364
rect 20300 27806 20302 27858
rect 20354 27806 20356 27858
rect 20076 27134 20078 27186
rect 20130 27134 20132 27186
rect 20076 27122 20132 27134
rect 20188 27188 20244 27198
rect 20188 27074 20244 27132
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 20188 27010 20244 27022
rect 20300 27076 20356 27806
rect 20636 28084 20692 28094
rect 20636 27748 20692 28028
rect 20748 28082 20804 29372
rect 20972 28644 21028 28654
rect 20972 28550 21028 28588
rect 20748 28030 20750 28082
rect 20802 28030 20804 28082
rect 20748 28018 20804 28030
rect 21084 27972 21140 32284
rect 21196 29428 21252 33852
rect 21308 32450 21364 32462
rect 21308 32398 21310 32450
rect 21362 32398 21364 32450
rect 21308 32340 21364 32398
rect 21308 32274 21364 32284
rect 21196 29362 21252 29372
rect 21420 28420 21476 34300
rect 21756 34132 21812 34142
rect 21532 32676 21588 32686
rect 21532 30994 21588 32620
rect 21756 32676 21812 34076
rect 22092 33458 22148 37100
rect 22092 33406 22094 33458
rect 22146 33406 22148 33458
rect 22092 33236 22148 33406
rect 22092 33170 22148 33180
rect 21868 32788 21924 32798
rect 21868 32786 22148 32788
rect 21868 32734 21870 32786
rect 21922 32734 22148 32786
rect 21868 32732 22148 32734
rect 21868 32722 21924 32732
rect 21756 32610 21812 32620
rect 21644 32562 21700 32574
rect 21644 32510 21646 32562
rect 21698 32510 21700 32562
rect 21644 31890 21700 32510
rect 21980 32562 22036 32574
rect 21980 32510 21982 32562
rect 22034 32510 22036 32562
rect 21980 32004 22036 32510
rect 21644 31838 21646 31890
rect 21698 31838 21700 31890
rect 21644 31826 21700 31838
rect 21756 31948 22036 32004
rect 21756 31892 21812 31948
rect 21644 31332 21700 31342
rect 21644 31218 21700 31276
rect 21644 31166 21646 31218
rect 21698 31166 21700 31218
rect 21644 31154 21700 31166
rect 21532 30942 21534 30994
rect 21586 30942 21588 30994
rect 21532 30930 21588 30942
rect 21756 30434 21812 31836
rect 21868 31780 21924 31790
rect 21868 31686 21924 31724
rect 22092 31220 22148 32732
rect 22204 32228 22260 37772
rect 22204 32162 22260 32172
rect 22204 32004 22260 32014
rect 22316 32004 22372 38612
rect 22428 37940 22484 37950
rect 22540 37940 22596 38780
rect 23212 38164 23268 38174
rect 23212 38070 23268 38108
rect 22428 37938 22596 37940
rect 22428 37886 22430 37938
rect 22482 37886 22596 37938
rect 22428 37884 22596 37886
rect 22428 37874 22484 37884
rect 22652 37380 22708 37390
rect 22652 37286 22708 37324
rect 23436 37380 23492 37390
rect 23436 37266 23492 37324
rect 23436 37214 23438 37266
rect 23490 37214 23492 37266
rect 23436 37202 23492 37214
rect 23212 34916 23268 34926
rect 23212 34822 23268 34860
rect 22428 34804 22484 34814
rect 22428 34710 22484 34748
rect 23548 33572 23604 40348
rect 23660 38724 23716 38734
rect 23660 38722 23828 38724
rect 23660 38670 23662 38722
rect 23714 38670 23828 38722
rect 23660 38668 23828 38670
rect 23660 38658 23716 38668
rect 23772 38612 23828 38668
rect 23772 36260 23828 38556
rect 23996 38164 24052 38174
rect 23996 38050 24052 38108
rect 23996 37998 23998 38050
rect 24050 37998 24052 38050
rect 23996 37986 24052 37998
rect 24108 37378 24164 42590
rect 24108 37326 24110 37378
rect 24162 37326 24164 37378
rect 24108 37314 24164 37326
rect 23884 37266 23940 37278
rect 23884 37214 23886 37266
rect 23938 37214 23940 37266
rect 23884 36708 23940 37214
rect 24220 36820 24276 43652
rect 24332 42866 24388 44268
rect 24556 44322 24612 44334
rect 24556 44270 24558 44322
rect 24610 44270 24612 44322
rect 24556 43540 24612 44270
rect 24556 43474 24612 43484
rect 24668 44322 24724 44380
rect 24668 44270 24670 44322
rect 24722 44270 24724 44322
rect 24332 42814 24334 42866
rect 24386 42814 24388 42866
rect 24332 42802 24388 42814
rect 24332 42530 24388 42542
rect 24332 42478 24334 42530
rect 24386 42478 24388 42530
rect 24332 42196 24388 42478
rect 24332 42130 24388 42140
rect 24668 40962 24724 44270
rect 25004 42868 25060 46172
rect 25116 45890 25172 45902
rect 25116 45838 25118 45890
rect 25170 45838 25172 45890
rect 25116 44100 25172 45838
rect 25116 44034 25172 44044
rect 25004 42802 25060 42812
rect 25228 42196 25284 50428
rect 26124 50484 26180 50542
rect 26236 50596 26292 51438
rect 26460 51154 26516 51166
rect 26460 51102 26462 51154
rect 26514 51102 26516 51154
rect 26460 50932 26516 51102
rect 26460 50866 26516 50876
rect 26348 50596 26404 50606
rect 26236 50540 26348 50596
rect 26348 50502 26404 50540
rect 26124 50418 26180 50428
rect 26572 50372 26628 55132
rect 26796 55122 26852 55132
rect 27132 55186 27188 55244
rect 27132 55134 27134 55186
rect 27186 55134 27188 55186
rect 27132 55122 27188 55134
rect 29596 55186 29652 55198
rect 29596 55134 29598 55186
rect 29650 55134 29652 55186
rect 28028 53284 28084 53294
rect 26796 51938 26852 51950
rect 26796 51886 26798 51938
rect 26850 51886 26852 51938
rect 26796 50932 26852 51886
rect 28028 51490 28084 53228
rect 29596 53284 29652 55134
rect 29932 55186 29988 56140
rect 29932 55134 29934 55186
rect 29986 55134 29988 55186
rect 29932 55122 29988 55134
rect 31052 55524 31108 55534
rect 31612 55468 31668 59200
rect 36988 56642 37044 59200
rect 43036 57092 43092 59200
rect 43036 57026 43092 57036
rect 43596 57092 43652 57102
rect 36988 56590 36990 56642
rect 37042 56590 37044 56642
rect 36988 56578 37044 56590
rect 37884 56642 37940 56654
rect 37884 56590 37886 56642
rect 37938 56590 37940 56642
rect 29596 53218 29652 53228
rect 28028 51438 28030 51490
rect 28082 51438 28084 51490
rect 28028 51426 28084 51438
rect 26796 50866 26852 50876
rect 27356 51378 27412 51390
rect 27356 51326 27358 51378
rect 27410 51326 27412 51378
rect 26460 50316 26628 50372
rect 27020 50484 27076 50494
rect 27356 50484 27412 51326
rect 27692 51266 27748 51278
rect 27692 51214 27694 51266
rect 27746 51214 27748 51266
rect 27468 50932 27524 50942
rect 27468 50706 27524 50876
rect 27468 50654 27470 50706
rect 27522 50654 27524 50706
rect 27468 50642 27524 50654
rect 27020 50482 27412 50484
rect 27020 50430 27022 50482
rect 27074 50430 27412 50482
rect 27020 50428 27412 50430
rect 26124 49812 26180 49822
rect 26124 49250 26180 49756
rect 26124 49198 26126 49250
rect 26178 49198 26180 49250
rect 26124 49186 26180 49198
rect 25228 42130 25284 42140
rect 25340 48132 25396 48142
rect 25004 41188 25060 41198
rect 25004 41094 25060 41132
rect 24668 40910 24670 40962
rect 24722 40910 24724 40962
rect 24668 40898 24724 40910
rect 25340 40852 25396 48076
rect 26124 48130 26180 48142
rect 26124 48078 26126 48130
rect 26178 48078 26180 48130
rect 26124 48020 26180 48078
rect 26124 47954 26180 47964
rect 25564 47796 25620 47806
rect 25564 47570 25620 47740
rect 25564 47518 25566 47570
rect 25618 47518 25620 47570
rect 25452 46676 25508 46686
rect 25564 46676 25620 47518
rect 26460 47570 26516 50316
rect 26796 49924 26852 49934
rect 27020 49924 27076 50428
rect 26852 49868 26964 49924
rect 26796 49830 26852 49868
rect 26572 49812 26628 49822
rect 26572 49718 26628 49756
rect 26684 49810 26740 49822
rect 26684 49758 26686 49810
rect 26738 49758 26740 49810
rect 26684 49700 26740 49758
rect 26684 48916 26740 49644
rect 26796 49140 26852 49150
rect 26796 49046 26852 49084
rect 26908 49026 26964 49868
rect 27020 49858 27076 49868
rect 27692 49810 27748 51214
rect 29036 51268 29092 51278
rect 28252 51156 28308 51166
rect 28140 49924 28196 49934
rect 28140 49830 28196 49868
rect 27692 49758 27694 49810
rect 27746 49758 27748 49810
rect 27692 49700 27748 49758
rect 28252 49810 28308 51100
rect 29036 50428 29092 51212
rect 29484 50708 29540 50718
rect 29036 50372 29316 50428
rect 28252 49758 28254 49810
rect 28306 49758 28308 49810
rect 28252 49746 28308 49758
rect 27692 49634 27748 49644
rect 27916 49698 27972 49710
rect 27916 49646 27918 49698
rect 27970 49646 27972 49698
rect 26908 48974 26910 49026
rect 26962 48974 26964 49026
rect 26908 48962 26964 48974
rect 27244 49586 27300 49598
rect 27244 49534 27246 49586
rect 27298 49534 27300 49586
rect 26684 48860 26852 48916
rect 26460 47518 26462 47570
rect 26514 47518 26516 47570
rect 26460 47506 26516 47518
rect 26684 48018 26740 48030
rect 26684 47966 26686 48018
rect 26738 47966 26740 48018
rect 26012 47460 26068 47470
rect 26684 47460 26740 47966
rect 26796 48020 26852 48860
rect 26908 48804 26964 48814
rect 26908 48242 26964 48748
rect 27132 48356 27188 48366
rect 27132 48262 27188 48300
rect 27244 48354 27300 49534
rect 27916 49140 27972 49646
rect 27916 49074 27972 49084
rect 27244 48302 27246 48354
rect 27298 48302 27300 48354
rect 27244 48290 27300 48302
rect 26908 48190 26910 48242
rect 26962 48190 26964 48242
rect 26908 48178 26964 48190
rect 27468 48020 27524 48030
rect 26796 47964 26964 48020
rect 26012 47458 26180 47460
rect 26012 47406 26014 47458
rect 26066 47406 26180 47458
rect 26012 47404 26180 47406
rect 26012 47394 26068 47404
rect 25900 46676 25956 46686
rect 25564 46674 25956 46676
rect 25564 46622 25902 46674
rect 25954 46622 25956 46674
rect 25564 46620 25956 46622
rect 25452 46114 25508 46620
rect 25900 46610 25956 46620
rect 26124 46674 26180 47404
rect 26684 47394 26740 47404
rect 26908 46786 26964 47964
rect 27468 47926 27524 47964
rect 26908 46734 26910 46786
rect 26962 46734 26964 46786
rect 26908 46722 26964 46734
rect 28476 47236 28532 47246
rect 26124 46622 26126 46674
rect 26178 46622 26180 46674
rect 26124 46564 26180 46622
rect 27244 46676 27300 46686
rect 27244 46582 27300 46620
rect 26124 46498 26180 46508
rect 26460 46562 26516 46574
rect 26460 46510 26462 46562
rect 26514 46510 26516 46562
rect 25452 46062 25454 46114
rect 25506 46062 25508 46114
rect 25452 46050 25508 46062
rect 26124 46004 26180 46014
rect 26124 45910 26180 45948
rect 26460 45332 26516 46510
rect 27356 46562 27412 46574
rect 27356 46510 27358 46562
rect 27410 46510 27412 46562
rect 27020 46004 27076 46014
rect 27020 45910 27076 45948
rect 26572 45892 26628 45902
rect 26572 45890 26740 45892
rect 26572 45838 26574 45890
rect 26626 45838 26740 45890
rect 26572 45836 26740 45838
rect 26572 45826 26628 45836
rect 26572 45332 26628 45342
rect 26460 45330 26628 45332
rect 26460 45278 26574 45330
rect 26626 45278 26628 45330
rect 26460 45276 26628 45278
rect 26572 45266 26628 45276
rect 25900 45218 25956 45230
rect 25900 45166 25902 45218
rect 25954 45166 25956 45218
rect 25676 44882 25732 44894
rect 25676 44830 25678 44882
rect 25730 44830 25732 44882
rect 25564 44436 25620 44446
rect 25564 44342 25620 44380
rect 25676 43540 25732 44830
rect 25900 44324 25956 45166
rect 26684 44994 26740 45836
rect 27356 45444 27412 46510
rect 28252 46228 28308 46238
rect 28252 45890 28308 46172
rect 28476 46116 28532 47180
rect 28476 46060 28644 46116
rect 28252 45838 28254 45890
rect 28306 45838 28308 45890
rect 28252 45826 28308 45838
rect 28476 45892 28532 45902
rect 28476 45798 28532 45836
rect 27356 45378 27412 45388
rect 28364 45666 28420 45678
rect 28588 45668 28644 46060
rect 28924 45890 28980 45902
rect 28924 45838 28926 45890
rect 28978 45838 28980 45890
rect 28364 45614 28366 45666
rect 28418 45614 28420 45666
rect 26684 44942 26686 44994
rect 26738 44942 26740 44994
rect 25788 44100 25844 44110
rect 25788 43650 25844 44044
rect 25900 43762 25956 44268
rect 26012 44882 26068 44894
rect 26012 44830 26014 44882
rect 26066 44830 26068 44882
rect 26012 44322 26068 44830
rect 26012 44270 26014 44322
rect 26066 44270 26068 44322
rect 26012 44258 26068 44270
rect 26124 44436 26180 44446
rect 25900 43710 25902 43762
rect 25954 43710 25956 43762
rect 25900 43698 25956 43710
rect 26124 43762 26180 44380
rect 26460 44324 26516 44334
rect 26684 44324 26740 44942
rect 26460 44322 26740 44324
rect 26460 44270 26462 44322
rect 26514 44270 26740 44322
rect 26460 44268 26740 44270
rect 26460 44258 26516 44268
rect 28364 44212 28420 45614
rect 26124 43710 26126 43762
rect 26178 43710 26180 43762
rect 26124 43698 26180 43710
rect 28252 44156 28420 44212
rect 28476 45612 28644 45668
rect 28700 45668 28756 45678
rect 25788 43598 25790 43650
rect 25842 43598 25844 43650
rect 25788 43586 25844 43598
rect 25676 43446 25732 43484
rect 26348 42868 26404 42878
rect 26348 42774 26404 42812
rect 26908 42868 26964 42878
rect 28252 42868 28308 44156
rect 28476 43650 28532 45612
rect 28476 43598 28478 43650
rect 28530 43598 28532 43650
rect 28476 43586 28532 43598
rect 28476 42980 28532 42990
rect 28364 42868 28420 42878
rect 28252 42866 28420 42868
rect 28252 42814 28366 42866
rect 28418 42814 28420 42866
rect 28252 42812 28420 42814
rect 26908 42754 26964 42812
rect 28364 42802 28420 42812
rect 26908 42702 26910 42754
rect 26962 42702 26964 42754
rect 26908 42690 26964 42702
rect 28140 42756 28196 42766
rect 28140 42662 28196 42700
rect 27244 42530 27300 42542
rect 27244 42478 27246 42530
rect 27298 42478 27300 42530
rect 27244 42420 27300 42478
rect 27244 42354 27300 42364
rect 26012 42196 26068 42234
rect 26012 42130 26068 42140
rect 25788 41970 25844 41982
rect 25788 41918 25790 41970
rect 25842 41918 25844 41970
rect 25788 40964 25844 41918
rect 26012 41970 26068 41982
rect 26012 41918 26014 41970
rect 26066 41918 26068 41970
rect 25228 40796 25396 40852
rect 25676 40908 25844 40964
rect 25900 41748 25956 41758
rect 25900 41074 25956 41692
rect 26012 41412 26068 41918
rect 26348 41972 26404 41982
rect 26684 41972 26740 41982
rect 26348 41970 26740 41972
rect 26348 41918 26350 41970
rect 26402 41918 26686 41970
rect 26738 41918 26740 41970
rect 26348 41916 26740 41918
rect 26348 41906 26404 41916
rect 26012 41346 26068 41356
rect 25900 41022 25902 41074
rect 25954 41022 25956 41074
rect 25900 40964 25956 41022
rect 24332 40404 24388 40414
rect 24332 40310 24388 40348
rect 24668 40290 24724 40302
rect 24668 40238 24670 40290
rect 24722 40238 24724 40290
rect 24668 39396 24724 40238
rect 24668 39330 24724 39340
rect 24780 39394 24836 39406
rect 24780 39342 24782 39394
rect 24834 39342 24836 39394
rect 24332 38946 24388 38958
rect 24332 38894 24334 38946
rect 24386 38894 24388 38946
rect 24332 38836 24388 38894
rect 24332 38770 24388 38780
rect 24444 38834 24500 38846
rect 24444 38782 24446 38834
rect 24498 38782 24500 38834
rect 24332 38610 24388 38622
rect 24332 38558 24334 38610
rect 24386 38558 24388 38610
rect 24332 37938 24388 38558
rect 24444 38612 24500 38782
rect 24444 38546 24500 38556
rect 24780 38612 24836 39342
rect 24780 38546 24836 38556
rect 25004 38722 25060 38734
rect 25004 38670 25006 38722
rect 25058 38670 25060 38722
rect 25004 38276 25060 38670
rect 24332 37886 24334 37938
rect 24386 37886 24388 37938
rect 24332 37874 24388 37886
rect 24556 38220 25060 38276
rect 25228 38274 25284 40796
rect 25676 40290 25732 40908
rect 25788 40628 25844 40638
rect 25900 40628 25956 40908
rect 25788 40626 25956 40628
rect 25788 40574 25790 40626
rect 25842 40574 25956 40626
rect 25788 40572 25956 40574
rect 26348 41298 26404 41310
rect 26348 41246 26350 41298
rect 26402 41246 26404 41298
rect 26348 41076 26404 41246
rect 25788 40562 25844 40572
rect 25676 40238 25678 40290
rect 25730 40238 25732 40290
rect 25676 40226 25732 40238
rect 26012 40180 26068 40190
rect 26348 40180 26404 41020
rect 26012 40178 26404 40180
rect 26012 40126 26014 40178
rect 26066 40126 26404 40178
rect 26012 40124 26404 40126
rect 26684 41188 26740 41916
rect 27244 41412 27300 41422
rect 27244 41318 27300 41356
rect 25228 38222 25230 38274
rect 25282 38222 25284 38274
rect 24556 37154 24612 38220
rect 25228 38210 25284 38222
rect 25340 39394 25396 39406
rect 25340 39342 25342 39394
rect 25394 39342 25396 39394
rect 25340 38276 25396 39342
rect 25788 39396 25844 39406
rect 25788 39302 25844 39340
rect 25788 38946 25844 38958
rect 25788 38894 25790 38946
rect 25842 38894 25844 38946
rect 25340 38210 25396 38220
rect 25452 38612 25508 38622
rect 24556 37102 24558 37154
rect 24610 37102 24612 37154
rect 24220 36764 24500 36820
rect 23884 36652 24388 36708
rect 24332 36594 24388 36652
rect 24332 36542 24334 36594
rect 24386 36542 24388 36594
rect 24332 36530 24388 36542
rect 24444 36372 24500 36764
rect 24220 36316 24500 36372
rect 24556 36372 24612 37102
rect 23660 36258 23828 36260
rect 23660 36206 23774 36258
rect 23826 36206 23828 36258
rect 23660 36204 23828 36206
rect 23660 34804 23716 36204
rect 23772 36194 23828 36204
rect 24108 36260 24164 36270
rect 24108 35698 24164 36204
rect 24108 35646 24110 35698
rect 24162 35646 24164 35698
rect 24108 35028 24164 35646
rect 24108 34962 24164 34972
rect 23772 34916 23828 34926
rect 23772 34822 23828 34860
rect 23660 34738 23716 34748
rect 23884 34802 23940 34814
rect 23884 34750 23886 34802
rect 23938 34750 23940 34802
rect 23548 33516 23828 33572
rect 22540 33460 22596 33470
rect 22540 33366 22596 33404
rect 23660 33348 23716 33358
rect 23548 33346 23716 33348
rect 23548 33294 23662 33346
rect 23714 33294 23716 33346
rect 23548 33292 23716 33294
rect 23100 33234 23156 33246
rect 23436 33236 23492 33246
rect 23100 33182 23102 33234
rect 23154 33182 23156 33234
rect 22988 33124 23044 33134
rect 22876 33012 22932 33022
rect 22876 32786 22932 32956
rect 22876 32734 22878 32786
rect 22930 32734 22932 32786
rect 22876 32722 22932 32734
rect 22652 32674 22708 32686
rect 22652 32622 22654 32674
rect 22706 32622 22708 32674
rect 22204 32002 22372 32004
rect 22204 31950 22206 32002
rect 22258 31950 22372 32002
rect 22204 31948 22372 31950
rect 22540 32562 22596 32574
rect 22540 32510 22542 32562
rect 22594 32510 22596 32562
rect 22204 31938 22260 31948
rect 22540 31892 22596 32510
rect 22652 32340 22708 32622
rect 22652 32274 22708 32284
rect 22540 31826 22596 31836
rect 22428 31780 22484 31790
rect 21756 30382 21758 30434
rect 21810 30382 21812 30434
rect 21756 30370 21812 30382
rect 21980 31164 22148 31220
rect 22204 31332 22260 31342
rect 21980 30324 22036 31164
rect 22092 30548 22148 30558
rect 22092 30434 22148 30492
rect 22092 30382 22094 30434
rect 22146 30382 22148 30434
rect 22092 30370 22148 30382
rect 21980 30098 22036 30268
rect 21980 30046 21982 30098
rect 22034 30046 22036 30098
rect 21980 30034 22036 30046
rect 21868 29652 21924 29662
rect 21532 29316 21588 29326
rect 21532 29222 21588 29260
rect 21868 29092 21924 29596
rect 21868 29026 21924 29036
rect 22204 28866 22260 31276
rect 22428 31218 22484 31724
rect 22988 31444 23044 33068
rect 23100 32340 23156 33182
rect 23100 32274 23156 32284
rect 23212 33234 23492 33236
rect 23212 33182 23438 33234
rect 23490 33182 23492 33234
rect 23212 33180 23492 33182
rect 23100 32116 23156 32126
rect 23100 32002 23156 32060
rect 23100 31950 23102 32002
rect 23154 31950 23156 32002
rect 23100 31938 23156 31950
rect 23212 31780 23268 33180
rect 23436 33170 23492 33180
rect 23324 32676 23380 32686
rect 23548 32676 23604 33292
rect 23660 33282 23716 33292
rect 23772 32788 23828 33516
rect 23884 33012 23940 34750
rect 24220 33348 24276 36316
rect 24556 36278 24612 36316
rect 24668 38052 24724 38062
rect 24668 37604 24724 37996
rect 25452 38050 25508 38556
rect 25452 37998 25454 38050
rect 25506 37998 25508 38050
rect 24668 37548 24948 37604
rect 24668 37266 24724 37548
rect 24668 37214 24670 37266
rect 24722 37214 24724 37266
rect 24668 35698 24724 37214
rect 24668 35646 24670 35698
rect 24722 35646 24724 35698
rect 24668 35634 24724 35646
rect 24780 37380 24836 37390
rect 24780 36370 24836 37324
rect 24780 36318 24782 36370
rect 24834 36318 24836 36370
rect 24332 35028 24388 35038
rect 24332 34934 24388 34972
rect 24780 34804 24836 36318
rect 24892 36370 24948 37548
rect 24892 36318 24894 36370
rect 24946 36318 24948 36370
rect 24892 36306 24948 36318
rect 25116 36260 25172 36270
rect 25004 36258 25172 36260
rect 25004 36206 25118 36258
rect 25170 36206 25172 36258
rect 25004 36204 25172 36206
rect 24780 34738 24836 34748
rect 24892 36148 24948 36158
rect 24892 35812 24948 36092
rect 24332 34354 24388 34366
rect 24332 34302 24334 34354
rect 24386 34302 24388 34354
rect 24332 33572 24388 34302
rect 24892 34354 24948 35756
rect 24892 34302 24894 34354
rect 24946 34302 24948 34354
rect 24892 34290 24948 34302
rect 24332 33506 24388 33516
rect 24556 34020 24612 34030
rect 24220 33292 24388 33348
rect 23884 32946 23940 32956
rect 23772 32732 23940 32788
rect 23324 32674 23604 32676
rect 23324 32622 23326 32674
rect 23378 32622 23604 32674
rect 23324 32620 23604 32622
rect 23324 32610 23380 32620
rect 23212 31714 23268 31724
rect 23548 31778 23604 32620
rect 23772 32564 23828 32574
rect 23772 32470 23828 32508
rect 23772 32340 23828 32350
rect 23548 31726 23550 31778
rect 23602 31726 23604 31778
rect 23548 31714 23604 31726
rect 23660 31892 23716 31902
rect 23660 31778 23716 31836
rect 23660 31726 23662 31778
rect 23714 31726 23716 31778
rect 23660 31714 23716 31726
rect 22988 31378 23044 31388
rect 23772 31666 23828 32284
rect 23772 31614 23774 31666
rect 23826 31614 23828 31666
rect 22428 31166 22430 31218
rect 22482 31166 22484 31218
rect 22428 31154 22484 31166
rect 23660 31332 23716 31342
rect 23660 31218 23716 31276
rect 23660 31166 23662 31218
rect 23714 31166 23716 31218
rect 23660 31154 23716 31166
rect 22764 31106 22820 31118
rect 22764 31054 22766 31106
rect 22818 31054 22820 31106
rect 22204 28814 22206 28866
rect 22258 28814 22260 28866
rect 22204 28802 22260 28814
rect 22316 30994 22372 31006
rect 22316 30942 22318 30994
rect 22370 30942 22372 30994
rect 21420 28354 21476 28364
rect 21532 28756 21588 28766
rect 21084 27916 21252 27972
rect 20636 27298 20692 27692
rect 20860 27858 20916 27870
rect 20860 27806 20862 27858
rect 20914 27806 20916 27858
rect 20860 27412 20916 27806
rect 20860 27346 20916 27356
rect 20636 27246 20638 27298
rect 20690 27246 20692 27298
rect 20636 27234 20692 27246
rect 20860 27076 20916 27086
rect 20300 27074 20580 27076
rect 20300 27022 20302 27074
rect 20354 27022 20580 27074
rect 20300 27020 20580 27022
rect 20300 27010 20356 27020
rect 19964 26852 20020 26862
rect 19292 26514 19460 26516
rect 19292 26462 19294 26514
rect 19346 26462 19460 26514
rect 19292 26460 19460 26462
rect 19628 26850 20020 26852
rect 19628 26798 19966 26850
rect 20018 26798 20020 26850
rect 19628 26796 20020 26798
rect 19292 26450 19348 26460
rect 19180 26290 19236 26302
rect 19180 26238 19182 26290
rect 19234 26238 19236 26290
rect 18956 26180 19012 26190
rect 18732 26066 18788 26078
rect 18732 26014 18734 26066
rect 18786 26014 18788 26066
rect 18732 25508 18788 26014
rect 18956 25620 19012 26124
rect 18956 25554 19012 25564
rect 18732 25442 18788 25452
rect 19068 25508 19124 25518
rect 18956 25282 19012 25294
rect 18956 25230 18958 25282
rect 19010 25230 19012 25282
rect 18956 24948 19012 25230
rect 18956 24882 19012 24892
rect 18956 24724 19012 24734
rect 18732 24612 18788 24622
rect 18732 24610 18900 24612
rect 18732 24558 18734 24610
rect 18786 24558 18900 24610
rect 18732 24556 18900 24558
rect 18732 24546 18788 24556
rect 18508 22540 18676 22596
rect 18844 24388 18900 24556
rect 18508 21924 18564 22540
rect 18732 22484 18788 22494
rect 18732 22390 18788 22428
rect 18620 22370 18676 22382
rect 18620 22318 18622 22370
rect 18674 22318 18676 22370
rect 18620 22148 18676 22318
rect 18732 22148 18788 22158
rect 18620 22092 18732 22148
rect 18732 22082 18788 22092
rect 18508 21868 18788 21924
rect 18284 21308 18452 21364
rect 18172 20972 18340 21028
rect 18172 20804 18228 20814
rect 18060 20802 18228 20804
rect 18060 20750 18174 20802
rect 18226 20750 18228 20802
rect 18060 20748 18228 20750
rect 18172 20738 18228 20748
rect 18284 20468 18340 20972
rect 18284 20402 18340 20412
rect 17724 20076 18004 20132
rect 18060 20356 18116 20366
rect 17612 19236 17668 19246
rect 17612 19142 17668 19180
rect 17276 17726 17278 17778
rect 17330 17726 17332 17778
rect 17276 17714 17332 17726
rect 17500 18676 17556 18686
rect 17388 17332 17444 17342
rect 17388 14754 17444 17276
rect 17500 17108 17556 18620
rect 17724 17892 17780 20076
rect 17948 19908 18004 19918
rect 17500 17042 17556 17052
rect 17612 17836 17780 17892
rect 17836 19122 17892 19134
rect 17836 19070 17838 19122
rect 17890 19070 17892 19122
rect 17500 16210 17556 16222
rect 17500 16158 17502 16210
rect 17554 16158 17556 16210
rect 17500 15540 17556 16158
rect 17500 15474 17556 15484
rect 17388 14702 17390 14754
rect 17442 14702 17444 14754
rect 17388 14690 17444 14702
rect 17388 14532 17444 14542
rect 17612 14532 17668 17836
rect 17724 17668 17780 17678
rect 17836 17668 17892 19070
rect 17948 19012 18004 19852
rect 18060 19346 18116 20300
rect 18060 19294 18062 19346
rect 18114 19294 18116 19346
rect 18060 19282 18116 19294
rect 18172 20244 18228 20254
rect 17948 18946 18004 18956
rect 18172 18900 18228 20188
rect 18172 18834 18228 18844
rect 18284 19234 18340 19246
rect 18284 19182 18286 19234
rect 18338 19182 18340 19234
rect 17948 18676 18004 18686
rect 17948 17890 18004 18620
rect 18284 18676 18340 19182
rect 18284 18610 18340 18620
rect 18060 18450 18116 18462
rect 18060 18398 18062 18450
rect 18114 18398 18116 18450
rect 18060 18116 18116 18398
rect 18284 18452 18340 18462
rect 18284 18358 18340 18396
rect 18060 18050 18116 18060
rect 18172 18338 18228 18350
rect 18172 18286 18174 18338
rect 18226 18286 18228 18338
rect 17948 17838 17950 17890
rect 18002 17838 18004 17890
rect 17948 17826 18004 17838
rect 18172 17892 18228 18286
rect 18284 17892 18340 17902
rect 18172 17890 18340 17892
rect 18172 17838 18286 17890
rect 18338 17838 18340 17890
rect 18172 17836 18340 17838
rect 18284 17826 18340 17836
rect 17780 17612 17892 17668
rect 17724 17574 17780 17612
rect 18172 17108 18228 17118
rect 18172 17014 18228 17052
rect 17724 16996 17780 17006
rect 17724 16902 17780 16940
rect 18060 16996 18116 17006
rect 17948 16884 18004 16894
rect 17948 16790 18004 16828
rect 17836 15988 17892 15998
rect 17836 15894 17892 15932
rect 17948 15876 18004 15886
rect 17164 14476 17332 14532
rect 16828 13840 16884 13916
rect 16828 13188 16884 13198
rect 16828 13094 16884 13132
rect 16604 12402 16772 12404
rect 16604 12350 16606 12402
rect 16658 12350 16772 12402
rect 16604 12348 16772 12350
rect 16940 12962 16996 12974
rect 16940 12910 16942 12962
rect 16994 12910 16996 12962
rect 16604 12338 16660 12348
rect 16156 9996 16324 10052
rect 15932 9940 15988 9950
rect 15932 9826 15988 9884
rect 15932 9774 15934 9826
rect 15986 9774 15988 9826
rect 15932 9762 15988 9774
rect 16044 9828 16100 9838
rect 15820 9426 15876 9436
rect 15932 9268 15988 9278
rect 16044 9268 16100 9772
rect 16156 9826 16212 9838
rect 16156 9774 16158 9826
rect 16210 9774 16212 9826
rect 16156 9604 16212 9774
rect 16268 9716 16324 9996
rect 16268 9650 16324 9660
rect 16156 9538 16212 9548
rect 16268 9492 16324 9502
rect 15932 9266 16100 9268
rect 15932 9214 15934 9266
rect 15986 9214 16100 9266
rect 15932 9212 16100 9214
rect 16156 9268 16212 9278
rect 15932 9202 15988 9212
rect 16156 9174 16212 9212
rect 15820 9156 15876 9166
rect 15820 9062 15876 9100
rect 16156 8596 16212 8606
rect 15820 8372 15876 8382
rect 15820 8278 15876 8316
rect 16156 8370 16212 8540
rect 16156 8318 16158 8370
rect 16210 8318 16212 8370
rect 16156 8306 16212 8318
rect 15708 8092 15876 8148
rect 15820 8036 15876 8092
rect 15708 7362 15764 7374
rect 15708 7310 15710 7362
rect 15762 7310 15764 7362
rect 15708 6692 15764 7310
rect 15820 7028 15876 7980
rect 15876 6972 15988 7028
rect 15820 6962 15876 6972
rect 15708 6626 15764 6636
rect 15708 6468 15764 6478
rect 15708 6466 15876 6468
rect 15708 6414 15710 6466
rect 15762 6414 15876 6466
rect 15708 6412 15876 6414
rect 15708 6402 15764 6412
rect 15708 6244 15764 6254
rect 15708 6130 15764 6188
rect 15708 6078 15710 6130
rect 15762 6078 15764 6130
rect 15708 6066 15764 6078
rect 15820 6132 15876 6412
rect 15820 5684 15876 6076
rect 15820 5618 15876 5628
rect 15820 5236 15876 5246
rect 15820 5142 15876 5180
rect 15596 4116 15652 4732
rect 15820 4564 15876 4574
rect 15932 4564 15988 6972
rect 16268 6130 16324 9436
rect 16380 8428 16436 11788
rect 16716 12180 16772 12190
rect 16492 10052 16548 10062
rect 16492 8930 16548 9996
rect 16492 8878 16494 8930
rect 16546 8878 16548 8930
rect 16492 8596 16548 8878
rect 16492 8530 16548 8540
rect 16380 8372 16548 8428
rect 16380 7476 16436 7486
rect 16380 7252 16436 7420
rect 16380 7186 16436 7196
rect 16268 6078 16270 6130
rect 16322 6078 16324 6130
rect 16268 6066 16324 6078
rect 16380 6692 16436 6702
rect 16380 6578 16436 6636
rect 16380 6526 16382 6578
rect 16434 6526 16436 6578
rect 16380 5460 16436 6526
rect 15876 4508 15988 4564
rect 16156 5404 16436 5460
rect 15820 4432 15876 4508
rect 15596 4050 15652 4060
rect 16156 4228 16212 5404
rect 16268 5236 16324 5246
rect 16492 5236 16548 8372
rect 16716 8370 16772 12124
rect 16828 12178 16884 12190
rect 16828 12126 16830 12178
rect 16882 12126 16884 12178
rect 16828 11396 16884 12126
rect 16940 11844 16996 12910
rect 16940 11788 17108 11844
rect 16940 11618 16996 11630
rect 16940 11566 16942 11618
rect 16994 11566 16996 11618
rect 16940 11508 16996 11566
rect 16940 11442 16996 11452
rect 16828 11330 16884 11340
rect 16940 10948 16996 10958
rect 16940 10610 16996 10892
rect 16940 10558 16942 10610
rect 16994 10558 16996 10610
rect 16940 9492 16996 10558
rect 17052 10612 17108 11788
rect 17276 11620 17332 14476
rect 17388 14530 17668 14532
rect 17388 14478 17390 14530
rect 17442 14478 17668 14530
rect 17388 14476 17668 14478
rect 17836 15764 17892 15774
rect 17388 13524 17444 14476
rect 17388 12628 17444 13468
rect 17612 13972 17668 13982
rect 17612 12850 17668 13916
rect 17612 12798 17614 12850
rect 17666 12798 17668 12850
rect 17612 12786 17668 12798
rect 17724 13636 17780 13646
rect 17388 12562 17444 12572
rect 17276 11564 17668 11620
rect 17276 11506 17332 11564
rect 17276 11454 17278 11506
rect 17330 11454 17332 11506
rect 17276 11442 17332 11454
rect 17500 11396 17556 11406
rect 17052 10546 17108 10556
rect 17388 11394 17556 11396
rect 17388 11342 17502 11394
rect 17554 11342 17556 11394
rect 17388 11340 17556 11342
rect 16940 9436 17220 9492
rect 17052 9268 17108 9278
rect 17052 9174 17108 9212
rect 16716 8318 16718 8370
rect 16770 8318 16772 8370
rect 16716 8306 16772 8318
rect 16828 8484 16884 8494
rect 16716 6804 16772 6814
rect 16604 6690 16660 6702
rect 16604 6638 16606 6690
rect 16658 6638 16660 6690
rect 16604 6468 16660 6638
rect 16604 6402 16660 6412
rect 16268 5234 16548 5236
rect 16268 5182 16270 5234
rect 16322 5182 16548 5234
rect 16268 5180 16548 5182
rect 16604 5348 16660 5358
rect 16268 5170 16324 5180
rect 16604 4788 16660 5292
rect 16716 5012 16772 6748
rect 16828 5236 16884 8428
rect 16940 7474 16996 7486
rect 16940 7422 16942 7474
rect 16994 7422 16996 7474
rect 16940 6692 16996 7422
rect 16940 6626 16996 6636
rect 16940 5794 16996 5806
rect 16940 5742 16942 5794
rect 16994 5742 16996 5794
rect 16940 5348 16996 5742
rect 16940 5282 16996 5292
rect 16828 5170 16884 5180
rect 17164 5124 17220 9436
rect 17388 8484 17444 11340
rect 17500 11330 17556 11340
rect 17500 9826 17556 9838
rect 17500 9774 17502 9826
rect 17554 9774 17556 9826
rect 17500 8484 17556 9774
rect 17612 9604 17668 11564
rect 17724 11060 17780 13580
rect 17836 13076 17892 15708
rect 17948 15426 18004 15820
rect 17948 15374 17950 15426
rect 18002 15374 18004 15426
rect 17948 14308 18004 15374
rect 18060 15090 18116 16940
rect 18284 16772 18340 16782
rect 18284 16678 18340 16716
rect 18396 16548 18452 21308
rect 18620 20916 18676 20926
rect 18620 20822 18676 20860
rect 18508 20468 18564 20478
rect 18508 20242 18564 20412
rect 18508 20190 18510 20242
rect 18562 20190 18564 20242
rect 18508 19460 18564 20190
rect 18508 19394 18564 19404
rect 18620 19010 18676 19022
rect 18620 18958 18622 19010
rect 18674 18958 18676 19010
rect 18620 18900 18676 18958
rect 18620 18834 18676 18844
rect 18732 18226 18788 21868
rect 18732 18174 18734 18226
rect 18786 18174 18788 18226
rect 18732 18162 18788 18174
rect 18844 21026 18900 24332
rect 18956 23492 19012 24668
rect 19068 24722 19124 25452
rect 19068 24670 19070 24722
rect 19122 24670 19124 24722
rect 19068 24658 19124 24670
rect 18956 23426 19012 23436
rect 19068 24500 19124 24510
rect 19068 23268 19124 24444
rect 19180 24164 19236 26238
rect 19404 26292 19460 26302
rect 19404 26198 19460 26236
rect 19516 25620 19572 25630
rect 19628 25620 19684 26796
rect 19964 26786 20020 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 20412 26404 20468 26414
rect 20412 26310 20468 26348
rect 20300 26290 20356 26302
rect 20300 26238 20302 26290
rect 20354 26238 20356 26290
rect 20188 26068 20244 26078
rect 19852 25844 19908 25854
rect 19852 25730 19908 25788
rect 19852 25678 19854 25730
rect 19906 25678 19908 25730
rect 19852 25666 19908 25678
rect 19516 25618 19684 25620
rect 19516 25566 19518 25618
rect 19570 25566 19684 25618
rect 19516 25564 19684 25566
rect 19740 25620 19796 25630
rect 19516 25554 19572 25564
rect 19740 25506 19796 25564
rect 19740 25454 19742 25506
rect 19794 25454 19796 25506
rect 19740 25442 19796 25454
rect 20076 25506 20132 25518
rect 20076 25454 20078 25506
rect 20130 25454 20132 25506
rect 19404 25394 19460 25406
rect 19404 25342 19406 25394
rect 19458 25342 19460 25394
rect 19292 25060 19348 25070
rect 19292 24946 19348 25004
rect 19292 24894 19294 24946
rect 19346 24894 19348 24946
rect 19292 24882 19348 24894
rect 19180 24098 19236 24108
rect 19292 23940 19348 23978
rect 19068 23202 19124 23212
rect 19180 23884 19292 23940
rect 19068 23042 19124 23054
rect 19068 22990 19070 23042
rect 19122 22990 19124 23042
rect 18956 22596 19012 22606
rect 18956 22482 19012 22540
rect 18956 22430 18958 22482
rect 19010 22430 19012 22482
rect 18956 22418 19012 22430
rect 19068 22484 19124 22990
rect 19068 22418 19124 22428
rect 19180 22370 19236 23884
rect 19292 23874 19348 23884
rect 19292 23716 19348 23726
rect 19404 23716 19460 25342
rect 20076 25284 20132 25454
rect 20076 25218 20132 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 20188 24722 20244 26012
rect 20188 24670 20190 24722
rect 20242 24670 20244 24722
rect 20188 24658 20244 24670
rect 19628 24610 19684 24622
rect 19628 24558 19630 24610
rect 19682 24558 19684 24610
rect 19292 23714 19460 23716
rect 19292 23662 19294 23714
rect 19346 23662 19460 23714
rect 19292 23660 19460 23662
rect 19516 24500 19572 24510
rect 19292 23650 19348 23660
rect 19516 23492 19572 24444
rect 19628 24500 19684 24558
rect 19628 24498 19796 24500
rect 19628 24446 19630 24498
rect 19682 24446 19796 24498
rect 19628 24444 19796 24446
rect 19628 24434 19684 24444
rect 19180 22318 19182 22370
rect 19234 22318 19236 22370
rect 19180 22306 19236 22318
rect 19292 23436 19572 23492
rect 19628 23938 19684 23950
rect 19628 23886 19630 23938
rect 19682 23886 19684 23938
rect 19180 22148 19236 22158
rect 19180 21810 19236 22092
rect 19292 22146 19348 23436
rect 19516 23268 19572 23278
rect 19516 23174 19572 23212
rect 19292 22094 19294 22146
rect 19346 22094 19348 22146
rect 19292 22082 19348 22094
rect 19404 23044 19460 23054
rect 19404 22484 19460 22988
rect 19628 22484 19684 23886
rect 19740 23938 19796 24444
rect 20300 24388 20356 26238
rect 20524 26292 20580 27020
rect 20860 26982 20916 27020
rect 20524 26226 20580 26236
rect 20860 25508 20916 25518
rect 20860 25414 20916 25452
rect 20300 24322 20356 24332
rect 20524 25284 20580 25294
rect 19740 23886 19742 23938
rect 19794 23886 19796 23938
rect 19740 23874 19796 23886
rect 20300 24164 20356 24174
rect 20076 23826 20132 23838
rect 20076 23774 20078 23826
rect 20130 23774 20132 23826
rect 20076 23716 20132 23774
rect 20076 23650 20132 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19404 21812 19460 22428
rect 19180 21758 19182 21810
rect 19234 21758 19236 21810
rect 19180 21746 19236 21758
rect 19292 21756 19460 21812
rect 19516 22428 19684 22484
rect 20076 23380 20132 23390
rect 19068 21476 19124 21486
rect 19068 21382 19124 21420
rect 18844 20974 18846 21026
rect 18898 20974 18900 21026
rect 18844 18116 18900 20974
rect 19292 20916 19348 21756
rect 19516 21700 19572 22428
rect 20076 22370 20132 23324
rect 20076 22318 20078 22370
rect 20130 22318 20132 22370
rect 20076 22306 20132 22318
rect 19628 22260 19684 22270
rect 19628 21812 19684 22204
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 21812 20132 21822
rect 20300 21812 20356 24108
rect 20524 23938 20580 25228
rect 21196 24946 21252 27916
rect 21196 24894 21198 24946
rect 21250 24894 21252 24946
rect 21196 24882 21252 24894
rect 21420 27076 21476 27086
rect 21084 24834 21140 24846
rect 21084 24782 21086 24834
rect 21138 24782 21140 24834
rect 20524 23886 20526 23938
rect 20578 23886 20580 23938
rect 20524 23874 20580 23886
rect 20860 24724 20916 24734
rect 20860 23938 20916 24668
rect 20860 23886 20862 23938
rect 20914 23886 20916 23938
rect 20748 23828 20804 23838
rect 20748 23734 20804 23772
rect 20860 23378 20916 23886
rect 20860 23326 20862 23378
rect 20914 23326 20916 23378
rect 20860 23314 20916 23326
rect 20412 23266 20468 23278
rect 20412 23214 20414 23266
rect 20466 23214 20468 23266
rect 20412 23044 20468 23214
rect 20636 23266 20692 23278
rect 20636 23214 20638 23266
rect 20690 23214 20692 23266
rect 20636 23156 20692 23214
rect 20636 23090 20692 23100
rect 20412 22978 20468 22988
rect 20860 22708 20916 22718
rect 20636 22484 20692 22494
rect 20636 22370 20692 22428
rect 20636 22318 20638 22370
rect 20690 22318 20692 22370
rect 20636 22260 20692 22318
rect 20636 22194 20692 22204
rect 19628 21756 20076 21812
rect 19516 21644 19684 21700
rect 20076 21680 20132 21756
rect 20188 21756 20356 21812
rect 19404 21588 19460 21598
rect 19404 21494 19460 21532
rect 19292 20850 19348 20860
rect 19180 20692 19236 20702
rect 19180 20598 19236 20636
rect 19516 20692 19572 20702
rect 19516 20598 19572 20636
rect 19068 20020 19124 20030
rect 19628 20020 19684 21644
rect 19852 21028 19908 21038
rect 20076 21028 20132 21038
rect 19852 21026 20132 21028
rect 19852 20974 19854 21026
rect 19906 20974 20078 21026
rect 20130 20974 20132 21026
rect 19852 20972 20132 20974
rect 19852 20962 19908 20972
rect 20076 20962 20132 20972
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20242 20244 21756
rect 20860 21698 20916 22652
rect 21084 22484 21140 24782
rect 21308 24052 21364 24062
rect 21196 23154 21252 23166
rect 21196 23102 21198 23154
rect 21250 23102 21252 23154
rect 21196 22820 21252 23102
rect 21196 22754 21252 22764
rect 21084 22418 21140 22428
rect 21308 22372 21364 23996
rect 20860 21646 20862 21698
rect 20914 21646 20916 21698
rect 20860 21634 20916 21646
rect 21196 22316 21364 22372
rect 20524 21588 20580 21598
rect 20524 21494 20580 21532
rect 21084 21362 21140 21374
rect 21084 21310 21086 21362
rect 21138 21310 21140 21362
rect 20748 21252 20804 21262
rect 20636 20916 20692 20926
rect 20636 20822 20692 20860
rect 20188 20190 20190 20242
rect 20242 20190 20244 20242
rect 19852 20130 19908 20142
rect 19852 20078 19854 20130
rect 19906 20078 19908 20130
rect 19740 20020 19796 20030
rect 19628 20018 19796 20020
rect 19628 19966 19742 20018
rect 19794 19966 19796 20018
rect 19628 19964 19796 19966
rect 19068 19926 19124 19964
rect 19740 19684 19796 19964
rect 19740 19618 19796 19628
rect 19404 19572 19460 19582
rect 19404 19348 19460 19516
rect 19404 19282 19460 19292
rect 19628 19348 19684 19358
rect 19628 19254 19684 19292
rect 19516 19234 19572 19246
rect 19516 19182 19518 19234
rect 19570 19182 19572 19234
rect 19292 19122 19348 19134
rect 19292 19070 19294 19122
rect 19346 19070 19348 19122
rect 19180 18452 19236 18462
rect 18844 18050 18900 18060
rect 18956 18450 19236 18452
rect 18956 18398 19182 18450
rect 19234 18398 19236 18450
rect 18956 18396 19236 18398
rect 18844 17442 18900 17454
rect 18844 17390 18846 17442
rect 18898 17390 18900 17442
rect 18844 17108 18900 17390
rect 18844 17042 18900 17052
rect 18844 16884 18900 16894
rect 18844 16790 18900 16828
rect 18172 16492 18452 16548
rect 18172 16210 18228 16492
rect 18172 16158 18174 16210
rect 18226 16158 18228 16210
rect 18172 16146 18228 16158
rect 18284 16212 18340 16222
rect 18284 16098 18340 16156
rect 18284 16046 18286 16098
rect 18338 16046 18340 16098
rect 18284 16034 18340 16046
rect 18396 15988 18452 15998
rect 18284 15764 18340 15774
rect 18172 15540 18228 15550
rect 18172 15446 18228 15484
rect 18060 15038 18062 15090
rect 18114 15038 18116 15090
rect 18060 15026 18116 15038
rect 18284 14756 18340 15708
rect 18396 15316 18452 15932
rect 18620 15540 18676 15550
rect 18956 15540 19012 18396
rect 19180 18386 19236 18396
rect 19292 18340 19348 19070
rect 19404 18452 19460 18462
rect 19404 18358 19460 18396
rect 19180 17556 19236 17566
rect 19180 17462 19236 17500
rect 19292 17108 19348 18284
rect 19292 17042 19348 17052
rect 19404 16884 19460 16894
rect 19292 16882 19460 16884
rect 19292 16830 19406 16882
rect 19458 16830 19460 16882
rect 19292 16828 19460 16830
rect 19292 16548 19348 16828
rect 19404 16818 19460 16828
rect 19516 16660 19572 19182
rect 19628 19124 19684 19134
rect 19628 18676 19684 19068
rect 19852 19012 19908 20078
rect 20188 19236 20244 20190
rect 20300 20802 20356 20814
rect 20300 20750 20302 20802
rect 20354 20750 20356 20802
rect 20300 19460 20356 20750
rect 20524 20580 20580 20590
rect 20524 20578 20692 20580
rect 20524 20526 20526 20578
rect 20578 20526 20692 20578
rect 20524 20524 20692 20526
rect 20524 20514 20580 20524
rect 20524 20356 20580 20366
rect 20524 19906 20580 20300
rect 20636 20020 20692 20524
rect 20748 20578 20804 21196
rect 20748 20526 20750 20578
rect 20802 20526 20804 20578
rect 20748 20468 20804 20526
rect 20748 20402 20804 20412
rect 20972 20020 21028 20030
rect 20636 20018 21028 20020
rect 20636 19966 20974 20018
rect 21026 19966 21028 20018
rect 20636 19964 21028 19966
rect 20524 19854 20526 19906
rect 20578 19854 20580 19906
rect 20300 19404 20468 19460
rect 20300 19236 20356 19246
rect 20188 19234 20356 19236
rect 20188 19182 20302 19234
rect 20354 19182 20356 19234
rect 20188 19180 20356 19182
rect 20300 19170 20356 19180
rect 19852 18946 19908 18956
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19628 18620 19908 18676
rect 19628 18452 19684 18462
rect 19628 17668 19684 18396
rect 19628 16884 19684 17612
rect 19740 17892 19796 17902
rect 19740 17666 19796 17836
rect 19740 17614 19742 17666
rect 19794 17614 19796 17666
rect 19740 17602 19796 17614
rect 19852 17554 19908 18620
rect 20412 18564 20468 19404
rect 20412 18498 20468 18508
rect 20412 17780 20468 17790
rect 20412 17686 20468 17724
rect 20524 17556 20580 19854
rect 20860 19684 20916 19694
rect 20748 19346 20804 19358
rect 20748 19294 20750 19346
rect 20802 19294 20804 19346
rect 20748 18674 20804 19294
rect 20748 18622 20750 18674
rect 20802 18622 20804 18674
rect 20748 18610 20804 18622
rect 20860 18676 20916 19628
rect 20972 19236 21028 19964
rect 21084 19908 21140 21310
rect 21084 19842 21140 19852
rect 20972 19180 21140 19236
rect 20860 18674 21028 18676
rect 20860 18622 20862 18674
rect 20914 18622 21028 18674
rect 20860 18620 21028 18622
rect 20860 18610 20916 18620
rect 19852 17502 19854 17554
rect 19906 17502 19908 17554
rect 19852 17490 19908 17502
rect 20412 17500 20580 17556
rect 20636 18450 20692 18462
rect 20636 18398 20638 18450
rect 20690 18398 20692 18450
rect 20076 17444 20132 17454
rect 20076 17442 20244 17444
rect 20076 17390 20078 17442
rect 20130 17390 20244 17442
rect 20076 17388 20244 17390
rect 20076 17378 20132 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 20188 17106 20244 17388
rect 20188 17054 20190 17106
rect 20242 17054 20244 17106
rect 20188 17042 20244 17054
rect 19964 16994 20020 17006
rect 19964 16942 19966 16994
rect 20018 16942 20020 16994
rect 19740 16884 19796 16894
rect 19684 16882 19796 16884
rect 19684 16830 19742 16882
rect 19794 16830 19796 16882
rect 19684 16828 19796 16830
rect 19628 16752 19684 16828
rect 19740 16818 19796 16828
rect 19964 16884 20020 16942
rect 19852 16770 19908 16782
rect 19292 16482 19348 16492
rect 19404 16604 19572 16660
rect 19852 16718 19854 16770
rect 19906 16718 19908 16770
rect 19852 16660 19908 16718
rect 19068 16100 19124 16138
rect 19068 16034 19124 16044
rect 19180 15874 19236 15886
rect 19180 15822 19182 15874
rect 19234 15822 19236 15874
rect 19180 15652 19236 15822
rect 19180 15586 19236 15596
rect 19292 15874 19348 15886
rect 19292 15822 19294 15874
rect 19346 15822 19348 15874
rect 18396 15222 18452 15260
rect 18508 15314 18564 15326
rect 18508 15262 18510 15314
rect 18562 15262 18564 15314
rect 18508 14980 18564 15262
rect 18620 15092 18676 15484
rect 18844 15484 19012 15540
rect 18620 15036 18788 15092
rect 18508 14756 18564 14924
rect 18172 14700 18340 14756
rect 18396 14700 18564 14756
rect 18060 14644 18116 14654
rect 18060 14550 18116 14588
rect 17948 14242 18004 14252
rect 18172 13970 18228 14700
rect 18172 13918 18174 13970
rect 18226 13918 18228 13970
rect 17836 12404 17892 13020
rect 17948 13412 18004 13422
rect 17948 12962 18004 13356
rect 17948 12910 17950 12962
rect 18002 12910 18004 12962
rect 17948 12898 18004 12910
rect 18060 12516 18116 12526
rect 17948 12404 18004 12414
rect 17836 12402 18004 12404
rect 17836 12350 17950 12402
rect 18002 12350 18004 12402
rect 17836 12348 18004 12350
rect 17948 12338 18004 12348
rect 17724 10994 17780 11004
rect 17948 10836 18004 10846
rect 17948 10742 18004 10780
rect 18060 10052 18116 12460
rect 18172 10836 18228 13918
rect 18284 14420 18340 14430
rect 18284 13636 18340 14364
rect 18284 13570 18340 13580
rect 18396 12180 18452 14700
rect 18732 14418 18788 15036
rect 18732 14366 18734 14418
rect 18786 14366 18788 14418
rect 18732 14354 18788 14366
rect 18508 14308 18564 14318
rect 18508 12404 18564 14252
rect 18844 14196 18900 15484
rect 19292 14980 19348 15822
rect 19404 15148 19460 16604
rect 19852 16594 19908 16604
rect 19516 15876 19572 15886
rect 19964 15876 20020 16828
rect 19516 15782 19572 15820
rect 19628 15820 20020 15876
rect 20188 16548 20244 16558
rect 19628 15764 19684 15820
rect 19628 15698 19684 15708
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19516 15428 19572 15438
rect 19516 15314 19572 15372
rect 20188 15428 20244 16492
rect 20188 15362 20244 15372
rect 19516 15262 19518 15314
rect 19570 15262 19572 15314
rect 19516 15250 19572 15262
rect 19852 15314 19908 15326
rect 19852 15262 19854 15314
rect 19906 15262 19908 15314
rect 19852 15148 19908 15262
rect 19404 15092 19796 15148
rect 19852 15092 20020 15148
rect 19292 14914 19348 14924
rect 19068 14644 19124 14654
rect 19068 14550 19124 14588
rect 19628 14530 19684 14542
rect 19628 14478 19630 14530
rect 19682 14478 19684 14530
rect 18956 14308 19012 14318
rect 18956 14214 19012 14252
rect 19180 14308 19236 14318
rect 19180 14214 19236 14252
rect 18620 14140 18900 14196
rect 19068 14196 19124 14206
rect 18620 13074 18676 14140
rect 18732 13860 18788 13870
rect 18732 13766 18788 13804
rect 18620 13022 18622 13074
rect 18674 13022 18676 13074
rect 18620 13010 18676 13022
rect 18732 13188 18788 13198
rect 19068 13188 19124 14140
rect 19628 14196 19684 14478
rect 19740 14532 19796 15092
rect 19852 14756 19908 14766
rect 19852 14642 19908 14700
rect 19852 14590 19854 14642
rect 19906 14590 19908 14642
rect 19852 14578 19908 14590
rect 19740 14466 19796 14476
rect 19964 14532 20020 15092
rect 20412 14754 20468 17500
rect 20636 17332 20692 18398
rect 20636 17266 20692 17276
rect 20748 18228 20804 18238
rect 20748 16882 20804 18172
rect 20860 17444 20916 17454
rect 20860 17350 20916 17388
rect 20748 16830 20750 16882
rect 20802 16830 20804 16882
rect 20524 16100 20580 16110
rect 20524 16006 20580 16044
rect 20524 15540 20580 15550
rect 20524 15314 20580 15484
rect 20524 15262 20526 15314
rect 20578 15262 20580 15314
rect 20524 15250 20580 15262
rect 20412 14702 20414 14754
rect 20466 14702 20468 14754
rect 20412 14690 20468 14702
rect 19964 14466 20020 14476
rect 20076 14418 20132 14430
rect 20076 14366 20078 14418
rect 20130 14366 20132 14418
rect 20076 14308 20132 14366
rect 20300 14420 20356 14430
rect 20356 14364 20468 14420
rect 20300 14326 20356 14364
rect 20076 14242 20132 14252
rect 19628 14130 19684 14140
rect 19836 14140 20100 14150
rect 19516 14084 19572 14094
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19516 13970 19572 14028
rect 19516 13918 19518 13970
rect 19570 13918 19572 13970
rect 19516 13906 19572 13918
rect 19740 13972 19796 13982
rect 19180 13636 19236 13646
rect 19180 13542 19236 13580
rect 19068 13132 19236 13188
rect 18732 12962 18788 13132
rect 19068 12964 19124 12974
rect 18732 12910 18734 12962
rect 18786 12910 18788 12962
rect 18732 12898 18788 12910
rect 18844 12962 19124 12964
rect 18844 12910 19070 12962
rect 19122 12910 19124 12962
rect 18844 12908 19124 12910
rect 18620 12738 18676 12750
rect 18620 12686 18622 12738
rect 18674 12686 18676 12738
rect 18620 12628 18676 12686
rect 18620 12562 18676 12572
rect 18732 12740 18788 12750
rect 18508 12348 18676 12404
rect 18508 12180 18564 12190
rect 18396 12178 18564 12180
rect 18396 12126 18510 12178
rect 18562 12126 18564 12178
rect 18396 12124 18564 12126
rect 18620 12180 18676 12348
rect 18732 12402 18788 12684
rect 18732 12350 18734 12402
rect 18786 12350 18788 12402
rect 18732 12338 18788 12350
rect 18620 12124 18788 12180
rect 18396 11396 18452 11406
rect 18284 10836 18340 10846
rect 18172 10834 18340 10836
rect 18172 10782 18286 10834
rect 18338 10782 18340 10834
rect 18172 10780 18340 10782
rect 18284 10770 18340 10780
rect 18284 10612 18340 10622
rect 18060 9996 18228 10052
rect 17836 9828 17892 9838
rect 17836 9826 18116 9828
rect 17836 9774 17838 9826
rect 17890 9774 18116 9826
rect 17836 9772 18116 9774
rect 17836 9762 17892 9772
rect 17948 9604 18004 9614
rect 17612 9602 18004 9604
rect 17612 9550 17950 9602
rect 18002 9550 18004 9602
rect 17612 9548 18004 9550
rect 17612 8484 17668 8494
rect 17500 8428 17612 8484
rect 17388 8418 17444 8428
rect 17612 8418 17668 8428
rect 17500 8258 17556 8270
rect 17500 8206 17502 8258
rect 17554 8206 17556 8258
rect 17500 7476 17556 8206
rect 17836 8260 17892 9548
rect 17948 9538 18004 9548
rect 18060 9042 18116 9772
rect 18172 9154 18228 9996
rect 18172 9102 18174 9154
rect 18226 9102 18228 9154
rect 18172 9090 18228 9102
rect 18060 8990 18062 9042
rect 18114 8990 18116 9042
rect 17948 8484 18004 8494
rect 17948 8370 18004 8428
rect 17948 8318 17950 8370
rect 18002 8318 18004 8370
rect 17948 8306 18004 8318
rect 17836 8194 17892 8204
rect 17276 6804 17332 6814
rect 17276 6710 17332 6748
rect 16940 5068 17220 5124
rect 17276 5122 17332 5134
rect 17276 5070 17278 5122
rect 17330 5070 17332 5122
rect 16940 5012 16996 5068
rect 16716 4946 16772 4956
rect 16828 4956 16996 5012
rect 16828 4898 16884 4956
rect 16828 4846 16830 4898
rect 16882 4846 16884 4898
rect 16828 4788 16884 4846
rect 16604 4732 16884 4788
rect 17276 4788 17332 5070
rect 17276 4722 17332 4732
rect 16492 4564 16548 4574
rect 16492 4340 16548 4508
rect 16940 4564 16996 4574
rect 16940 4470 16996 4508
rect 16492 4274 16548 4284
rect 15372 3938 15428 3948
rect 15596 3668 15652 3678
rect 15260 3666 15652 3668
rect 15260 3614 15598 3666
rect 15650 3614 15652 3666
rect 15260 3612 15652 3614
rect 15596 3602 15652 3612
rect 16156 3666 16212 4172
rect 16156 3614 16158 3666
rect 16210 3614 16212 3666
rect 16156 3602 16212 3614
rect 16828 3668 16884 3678
rect 17500 3668 17556 7420
rect 17836 7700 17892 7710
rect 17836 6690 17892 7644
rect 18060 6804 18116 8990
rect 18284 8930 18340 10556
rect 18284 8878 18286 8930
rect 18338 8878 18340 8930
rect 18172 7476 18228 7486
rect 18172 7382 18228 7420
rect 18060 6748 18228 6804
rect 17836 6638 17838 6690
rect 17890 6638 17892 6690
rect 17836 6626 17892 6638
rect 18060 6580 18116 6590
rect 18060 6486 18116 6524
rect 18060 6356 18116 6366
rect 17836 5908 17892 5918
rect 17836 5234 17892 5852
rect 17836 5182 17838 5234
rect 17890 5182 17892 5234
rect 17836 5170 17892 5182
rect 17948 5794 18004 5806
rect 17948 5742 17950 5794
rect 18002 5742 18004 5794
rect 17724 4452 17780 4462
rect 17724 4358 17780 4396
rect 17948 4004 18004 5742
rect 18060 5348 18116 6300
rect 18060 5282 18116 5292
rect 18172 4564 18228 6748
rect 18284 6356 18340 8878
rect 18396 8370 18452 11340
rect 18508 10724 18564 12124
rect 18732 11060 18788 12124
rect 18844 12066 18900 12908
rect 19068 12898 19124 12908
rect 18956 12740 19012 12750
rect 19180 12740 19236 13132
rect 18956 12738 19124 12740
rect 18956 12686 18958 12738
rect 19010 12686 19124 12738
rect 18956 12684 19124 12686
rect 18956 12674 19012 12684
rect 19068 12516 19124 12684
rect 19180 12674 19236 12684
rect 19740 12962 19796 13916
rect 20300 13634 20356 13646
rect 20300 13582 20302 13634
rect 20354 13582 20356 13634
rect 20300 13412 20356 13582
rect 20300 13346 20356 13356
rect 20188 13076 20244 13086
rect 20188 12982 20244 13020
rect 19740 12910 19742 12962
rect 19794 12910 19796 12962
rect 19740 12740 19796 12910
rect 19740 12674 19796 12684
rect 19836 12572 20100 12582
rect 19516 12516 19572 12526
rect 19068 12460 19460 12516
rect 19404 12404 19460 12460
rect 19404 12338 19460 12348
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 18956 12292 19012 12302
rect 19180 12292 19236 12302
rect 18956 12290 19124 12292
rect 18956 12238 18958 12290
rect 19010 12238 19124 12290
rect 18956 12236 19124 12238
rect 18956 12226 19012 12236
rect 18844 12014 18846 12066
rect 18898 12014 18900 12066
rect 18844 12002 18900 12014
rect 19068 12180 19124 12236
rect 18956 11508 19012 11518
rect 18956 11394 19012 11452
rect 18956 11342 18958 11394
rect 19010 11342 19012 11394
rect 18956 11330 19012 11342
rect 18732 11004 19012 11060
rect 18844 10724 18900 10734
rect 18508 10722 18900 10724
rect 18508 10670 18846 10722
rect 18898 10670 18900 10722
rect 18508 10668 18900 10670
rect 18844 10658 18900 10668
rect 18956 10164 19012 11004
rect 18620 10108 19012 10164
rect 19068 10164 19124 12124
rect 19180 11788 19236 12236
rect 19516 12290 19572 12460
rect 19852 12404 19908 12442
rect 20412 12404 20468 14364
rect 19852 12338 19908 12348
rect 19964 12348 20468 12404
rect 20636 14308 20692 14318
rect 20636 12402 20692 14252
rect 20748 13412 20804 16830
rect 20972 16884 21028 18620
rect 20972 16818 21028 16828
rect 21084 18340 21140 19180
rect 20972 16660 21028 16670
rect 20972 16210 21028 16604
rect 21084 16548 21140 18284
rect 21084 16482 21140 16492
rect 20972 16158 20974 16210
rect 21026 16158 21028 16210
rect 20972 16146 21028 16158
rect 21084 16212 21140 16222
rect 21084 15988 21140 16156
rect 20972 15932 21140 15988
rect 20972 15202 21028 15932
rect 21084 15316 21140 15326
rect 21084 15222 21140 15260
rect 20972 15150 20974 15202
rect 21026 15150 21028 15202
rect 20972 15138 21028 15150
rect 21084 14980 21140 14990
rect 20972 14754 21028 14766
rect 20972 14702 20974 14754
rect 21026 14702 21028 14754
rect 20748 13346 20804 13356
rect 20860 14308 20916 14318
rect 20972 14308 21028 14702
rect 20860 14306 21028 14308
rect 20860 14254 20862 14306
rect 20914 14254 21028 14306
rect 20860 14252 21028 14254
rect 20860 12964 20916 14252
rect 21084 13634 21140 14924
rect 21196 13970 21252 22316
rect 21308 22148 21364 22158
rect 21308 21700 21364 22092
rect 21308 21586 21364 21644
rect 21308 21534 21310 21586
rect 21362 21534 21364 21586
rect 21308 21522 21364 21534
rect 21308 19460 21364 19470
rect 21308 18450 21364 19404
rect 21308 18398 21310 18450
rect 21362 18398 21364 18450
rect 21308 18386 21364 18398
rect 21196 13918 21198 13970
rect 21250 13918 21252 13970
rect 21196 13906 21252 13918
rect 21308 17220 21364 17230
rect 21308 16882 21364 17164
rect 21420 16996 21476 27020
rect 21532 25730 21588 28700
rect 21756 28756 21812 28766
rect 21756 28662 21812 28700
rect 22204 28642 22260 28654
rect 22204 28590 22206 28642
rect 22258 28590 22260 28642
rect 22092 28532 22148 28542
rect 21980 27970 22036 27982
rect 21980 27918 21982 27970
rect 22034 27918 22036 27970
rect 21644 27860 21700 27870
rect 21644 27300 21700 27804
rect 21980 27636 22036 27918
rect 21644 27186 21700 27244
rect 21644 27134 21646 27186
rect 21698 27134 21700 27186
rect 21644 27122 21700 27134
rect 21756 27580 22036 27636
rect 21532 25678 21534 25730
rect 21586 25678 21588 25730
rect 21532 25666 21588 25678
rect 21644 25282 21700 25294
rect 21644 25230 21646 25282
rect 21698 25230 21700 25282
rect 21644 24948 21700 25230
rect 21644 24882 21700 24892
rect 21644 24500 21700 24510
rect 21644 24050 21700 24444
rect 21644 23998 21646 24050
rect 21698 23998 21700 24050
rect 21644 23986 21700 23998
rect 21756 23492 21812 27580
rect 22092 27412 22148 28476
rect 22204 28308 22260 28590
rect 22204 28242 22260 28252
rect 22092 27186 22148 27356
rect 22092 27134 22094 27186
rect 22146 27134 22148 27186
rect 22092 27122 22148 27134
rect 22204 27860 22260 27870
rect 22316 27860 22372 30942
rect 22540 30996 22596 31006
rect 22540 30902 22596 30940
rect 22540 30772 22596 30782
rect 22428 29316 22484 29326
rect 22428 29222 22484 29260
rect 22540 29092 22596 30716
rect 22764 30548 22820 31054
rect 23548 30772 23604 30782
rect 22764 30482 22820 30492
rect 23436 30770 23604 30772
rect 23436 30718 23550 30770
rect 23602 30718 23604 30770
rect 23436 30716 23604 30718
rect 23212 30324 23268 30334
rect 23212 30210 23268 30268
rect 23212 30158 23214 30210
rect 23266 30158 23268 30210
rect 23212 30146 23268 30158
rect 23436 29988 23492 30716
rect 23548 30706 23604 30716
rect 23772 30770 23828 31614
rect 23884 31332 23940 32732
rect 24220 32676 24276 32686
rect 24220 32562 24276 32620
rect 24220 32510 24222 32562
rect 24274 32510 24276 32562
rect 24220 32498 24276 32510
rect 23884 31266 23940 31276
rect 23996 31780 24052 31790
rect 23772 30718 23774 30770
rect 23826 30718 23828 30770
rect 23772 30706 23828 30718
rect 23212 29932 23492 29988
rect 23660 30322 23716 30334
rect 23660 30270 23662 30322
rect 23714 30270 23716 30322
rect 22204 27858 22372 27860
rect 22204 27806 22206 27858
rect 22258 27806 22372 27858
rect 22204 27804 22372 27806
rect 22428 29036 22596 29092
rect 22652 29538 22708 29550
rect 22652 29486 22654 29538
rect 22706 29486 22708 29538
rect 22204 26402 22260 27804
rect 22204 26350 22206 26402
rect 22258 26350 22260 26402
rect 22204 26338 22260 26350
rect 22092 25394 22148 25406
rect 22092 25342 22094 25394
rect 22146 25342 22148 25394
rect 21868 25284 21924 25294
rect 21868 25190 21924 25228
rect 21980 25172 22036 25182
rect 21980 24722 22036 25116
rect 21980 24670 21982 24722
rect 22034 24670 22036 24722
rect 21980 24658 22036 24670
rect 21756 23426 21812 23436
rect 21756 23266 21812 23278
rect 21756 23214 21758 23266
rect 21810 23214 21812 23266
rect 21644 22484 21700 22494
rect 21644 22390 21700 22428
rect 21756 22260 21812 23214
rect 21980 23156 22036 23166
rect 21868 23154 22036 23156
rect 21868 23102 21982 23154
rect 22034 23102 22036 23154
rect 21868 23100 22036 23102
rect 21868 22372 21924 23100
rect 21980 23090 22036 23100
rect 22092 23042 22148 25342
rect 22316 23826 22372 23838
rect 22316 23774 22318 23826
rect 22370 23774 22372 23826
rect 22316 23268 22372 23774
rect 22428 23714 22484 29036
rect 22652 28868 22708 29486
rect 22764 29316 22820 29326
rect 22764 29222 22820 29260
rect 22652 28802 22708 28812
rect 22764 28866 22820 28878
rect 22764 28814 22766 28866
rect 22818 28814 22820 28866
rect 22652 28644 22708 28654
rect 22764 28644 22820 28814
rect 22652 28642 22820 28644
rect 22652 28590 22654 28642
rect 22706 28590 22820 28642
rect 22652 28588 22820 28590
rect 23100 28644 23156 28654
rect 22652 28578 22708 28588
rect 23100 28550 23156 28588
rect 22540 28532 22596 28542
rect 22540 27972 22596 28476
rect 22652 27972 22708 27982
rect 22540 27970 22708 27972
rect 22540 27918 22654 27970
rect 22706 27918 22708 27970
rect 22540 27916 22708 27918
rect 22652 27906 22708 27916
rect 22764 27972 22820 27982
rect 22764 27858 22820 27916
rect 22764 27806 22766 27858
rect 22818 27806 22820 27858
rect 22764 27794 22820 27806
rect 23100 27636 23156 27646
rect 22652 27300 22708 27310
rect 22652 27186 22708 27244
rect 22652 27134 22654 27186
rect 22706 27134 22708 27186
rect 22652 27122 22708 27134
rect 22652 26292 22708 26302
rect 22652 26198 22708 26236
rect 22652 25732 22708 25742
rect 22428 23662 22430 23714
rect 22482 23662 22484 23714
rect 22428 23650 22484 23662
rect 22540 25620 22596 25630
rect 22540 23380 22596 25564
rect 22652 25618 22708 25676
rect 23100 25620 23156 27580
rect 22652 25566 22654 25618
rect 22706 25566 22708 25618
rect 22652 25554 22708 25566
rect 22988 25564 23156 25620
rect 23212 25620 23268 29932
rect 23548 29652 23604 29662
rect 23548 29426 23604 29596
rect 23548 29374 23550 29426
rect 23602 29374 23604 29426
rect 23548 28868 23604 29374
rect 23660 29428 23716 30270
rect 23660 29362 23716 29372
rect 23772 29538 23828 29550
rect 23772 29486 23774 29538
rect 23826 29486 23828 29538
rect 23772 28980 23828 29486
rect 23996 29314 24052 31724
rect 24220 31332 24276 31342
rect 24108 30882 24164 30894
rect 24108 30830 24110 30882
rect 24162 30830 24164 30882
rect 24108 30770 24164 30830
rect 24108 30718 24110 30770
rect 24162 30718 24164 30770
rect 24108 30706 24164 30718
rect 24220 30322 24276 31276
rect 24332 30434 24388 33292
rect 24444 33236 24500 33246
rect 24444 33142 24500 33180
rect 24444 31892 24500 31902
rect 24444 31666 24500 31836
rect 24444 31614 24446 31666
rect 24498 31614 24500 31666
rect 24444 31602 24500 31614
rect 24556 31556 24612 33964
rect 24780 32450 24836 32462
rect 24780 32398 24782 32450
rect 24834 32398 24836 32450
rect 24780 32340 24836 32398
rect 24780 32274 24836 32284
rect 24668 31780 24724 31790
rect 24668 31686 24724 31724
rect 24556 31500 24724 31556
rect 24556 30996 24612 31006
rect 24556 30902 24612 30940
rect 24332 30382 24334 30434
rect 24386 30382 24388 30434
rect 24332 30370 24388 30382
rect 24220 30270 24222 30322
rect 24274 30270 24276 30322
rect 24220 30258 24276 30270
rect 24444 30212 24500 30222
rect 24444 30118 24500 30156
rect 24668 29988 24724 31500
rect 24780 31332 24836 31342
rect 24780 31218 24836 31276
rect 24780 31166 24782 31218
rect 24834 31166 24836 31218
rect 24780 31154 24836 31166
rect 24892 31108 24948 31118
rect 24892 31014 24948 31052
rect 24444 29932 24724 29988
rect 24780 30212 24836 30222
rect 24332 29428 24388 29438
rect 24220 29372 24332 29428
rect 23996 29262 23998 29314
rect 24050 29262 24052 29314
rect 23996 29250 24052 29262
rect 24108 29316 24164 29326
rect 24108 29222 24164 29260
rect 23772 28924 24052 28980
rect 23436 28812 23604 28868
rect 23660 28868 23716 28878
rect 23324 27074 23380 27086
rect 23324 27022 23326 27074
rect 23378 27022 23380 27074
rect 23324 26964 23380 27022
rect 23436 26964 23492 28812
rect 23660 28756 23716 28812
rect 23548 28700 23716 28756
rect 23772 28756 23828 28766
rect 23548 28642 23604 28700
rect 23772 28662 23828 28700
rect 23548 28590 23550 28642
rect 23602 28590 23604 28642
rect 23548 27186 23604 28590
rect 23660 28308 23716 28318
rect 23660 28082 23716 28252
rect 23660 28030 23662 28082
rect 23714 28030 23716 28082
rect 23660 27300 23716 28030
rect 23996 28084 24052 28924
rect 24108 28868 24164 28878
rect 24220 28868 24276 29372
rect 24332 29334 24388 29372
rect 24108 28866 24276 28868
rect 24108 28814 24110 28866
rect 24162 28814 24276 28866
rect 24108 28812 24276 28814
rect 24108 28802 24164 28812
rect 23996 28082 24164 28084
rect 23996 28030 23998 28082
rect 24050 28030 24164 28082
rect 23996 28028 24164 28030
rect 23996 28018 24052 28028
rect 23772 27300 23828 27310
rect 23660 27298 23828 27300
rect 23660 27246 23774 27298
rect 23826 27246 23828 27298
rect 23660 27244 23828 27246
rect 23548 27134 23550 27186
rect 23602 27134 23604 27186
rect 23548 27122 23604 27134
rect 23772 27076 23828 27244
rect 23772 27020 24052 27076
rect 23436 26908 23604 26964
rect 23324 26898 23380 26908
rect 23548 26852 23828 26908
rect 23436 26404 23492 26414
rect 22876 23828 22932 23838
rect 22316 23202 22372 23212
rect 22428 23324 22596 23380
rect 22652 23826 22932 23828
rect 22652 23774 22878 23826
rect 22930 23774 22932 23826
rect 22652 23772 22932 23774
rect 22092 22990 22094 23042
rect 22146 22990 22148 23042
rect 22092 22978 22148 22990
rect 22204 23154 22260 23166
rect 22204 23102 22206 23154
rect 22258 23102 22260 23154
rect 22204 23044 22260 23102
rect 21868 22306 21924 22316
rect 21756 22194 21812 22204
rect 21980 22258 22036 22270
rect 22204 22260 22260 22988
rect 21980 22206 21982 22258
rect 22034 22206 22036 22258
rect 21980 22148 22036 22206
rect 21980 22082 22036 22092
rect 22092 22204 22260 22260
rect 21868 22036 21924 22046
rect 21644 21810 21700 21822
rect 21644 21758 21646 21810
rect 21698 21758 21700 21810
rect 21644 21700 21700 21758
rect 21644 21634 21700 21644
rect 21532 21586 21588 21598
rect 21532 21534 21534 21586
rect 21586 21534 21588 21586
rect 21532 20692 21588 21534
rect 21532 18228 21588 20636
rect 21756 21476 21812 21486
rect 21644 20580 21700 20590
rect 21644 19458 21700 20524
rect 21756 20356 21812 21420
rect 21756 20290 21812 20300
rect 21868 20578 21924 21980
rect 22092 21924 22148 22204
rect 21980 21868 22148 21924
rect 21980 20804 22036 21868
rect 22092 21700 22148 21710
rect 22092 21606 22148 21644
rect 22316 21700 22372 21710
rect 22316 21140 22372 21644
rect 22316 21074 22372 21084
rect 21980 20748 22260 20804
rect 21868 20526 21870 20578
rect 21922 20526 21924 20578
rect 21868 20132 21924 20526
rect 21868 20066 21924 20076
rect 21868 19906 21924 19918
rect 21868 19854 21870 19906
rect 21922 19854 21924 19906
rect 21868 19684 21924 19854
rect 21868 19618 21924 19628
rect 21980 19908 22036 19918
rect 21644 19406 21646 19458
rect 21698 19406 21700 19458
rect 21644 19394 21700 19406
rect 21980 19458 22036 19852
rect 21980 19406 21982 19458
rect 22034 19406 22036 19458
rect 21980 19394 22036 19406
rect 21532 18162 21588 18172
rect 21756 19012 21812 19022
rect 21756 17780 21812 18956
rect 21980 18676 22036 18686
rect 21980 18582 22036 18620
rect 21868 18562 21924 18574
rect 21868 18510 21870 18562
rect 21922 18510 21924 18562
rect 21868 18340 21924 18510
rect 21868 18274 21924 18284
rect 21980 18452 22036 18462
rect 21756 17714 21812 17724
rect 21980 17666 22036 18396
rect 22092 18228 22148 18238
rect 22092 18134 22148 18172
rect 21980 17614 21982 17666
rect 22034 17614 22036 17666
rect 21980 17602 22036 17614
rect 21644 17554 21700 17566
rect 21644 17502 21646 17554
rect 21698 17502 21700 17554
rect 21644 17220 21700 17502
rect 21644 17154 21700 17164
rect 21756 17442 21812 17454
rect 21756 17390 21758 17442
rect 21810 17390 21812 17442
rect 21756 17332 21812 17390
rect 21420 16940 21588 16996
rect 21308 16830 21310 16882
rect 21362 16830 21364 16882
rect 21084 13582 21086 13634
rect 21138 13582 21140 13634
rect 21084 13570 21140 13582
rect 21196 13746 21252 13758
rect 21196 13694 21198 13746
rect 21250 13694 21252 13746
rect 21196 13636 21252 13694
rect 20860 12962 21028 12964
rect 20860 12910 20862 12962
rect 20914 12910 21028 12962
rect 20860 12908 21028 12910
rect 20860 12898 20916 12908
rect 20748 12852 20804 12862
rect 20748 12758 20804 12796
rect 20636 12350 20638 12402
rect 20690 12350 20692 12402
rect 19516 12238 19518 12290
rect 19570 12238 19572 12290
rect 19516 12226 19572 12238
rect 19852 12180 19908 12190
rect 19964 12180 20020 12348
rect 20636 12338 20692 12350
rect 19628 12178 20020 12180
rect 19628 12126 19854 12178
rect 19906 12126 20020 12178
rect 19628 12124 20020 12126
rect 20076 12178 20132 12190
rect 20076 12126 20078 12178
rect 20130 12126 20132 12178
rect 19628 11788 19684 12124
rect 19852 12114 19908 12124
rect 19180 11732 19460 11788
rect 19180 11394 19236 11406
rect 19180 11342 19182 11394
rect 19234 11342 19236 11394
rect 19180 11284 19236 11342
rect 19180 11218 19236 11228
rect 19180 10612 19236 10622
rect 19180 10518 19236 10556
rect 18620 9714 18676 10108
rect 18956 9828 19012 9838
rect 18956 9734 19012 9772
rect 18620 9662 18622 9714
rect 18674 9662 18676 9714
rect 18620 9268 18676 9662
rect 18620 9202 18676 9212
rect 18620 8932 18676 8942
rect 18396 8318 18398 8370
rect 18450 8318 18452 8370
rect 18396 8306 18452 8318
rect 18508 8484 18564 8494
rect 18284 6290 18340 6300
rect 18396 6916 18452 6926
rect 18396 6130 18452 6860
rect 18396 6078 18398 6130
rect 18450 6078 18452 6130
rect 18396 6066 18452 6078
rect 18284 5796 18340 5806
rect 18284 5234 18340 5740
rect 18284 5182 18286 5234
rect 18338 5182 18340 5234
rect 18284 5170 18340 5182
rect 18172 4498 18228 4508
rect 18396 4564 18452 4574
rect 18508 4564 18564 8428
rect 18620 8258 18676 8876
rect 19068 8820 19124 10108
rect 19180 9042 19236 9054
rect 19180 8990 19182 9042
rect 19234 8990 19236 9042
rect 19180 8932 19236 8990
rect 19404 9044 19460 11732
rect 19516 11732 19684 11788
rect 19852 11844 19908 11854
rect 19516 9268 19572 11732
rect 19628 11396 19684 11406
rect 19628 11302 19684 11340
rect 19852 11172 19908 11788
rect 19628 11116 19908 11172
rect 20076 11172 20132 12126
rect 20860 12178 20916 12190
rect 20860 12126 20862 12178
rect 20914 12126 20916 12178
rect 20076 11116 20244 11172
rect 19628 9492 19684 11116
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 20188 10836 20244 11116
rect 20076 10780 20244 10836
rect 19964 10610 20020 10622
rect 19964 10558 19966 10610
rect 20018 10558 20020 10610
rect 19852 10388 19908 10398
rect 19852 9938 19908 10332
rect 19852 9886 19854 9938
rect 19906 9886 19908 9938
rect 19852 9874 19908 9886
rect 19964 9940 20020 10558
rect 19964 9604 20020 9884
rect 20076 9604 20132 10780
rect 20412 10724 20468 10734
rect 20300 10612 20356 10622
rect 20300 10518 20356 10556
rect 20188 10500 20244 10510
rect 20188 10406 20244 10444
rect 20412 9940 20468 10668
rect 20860 10724 20916 12126
rect 20860 10658 20916 10668
rect 20972 11620 21028 12908
rect 21196 11732 21252 13580
rect 21308 13076 21364 16830
rect 21420 16772 21476 16782
rect 21420 16678 21476 16716
rect 21532 16548 21588 16940
rect 21420 16492 21588 16548
rect 21644 16884 21700 16894
rect 21756 16884 21812 17276
rect 21644 16882 21812 16884
rect 21644 16830 21646 16882
rect 21698 16830 21812 16882
rect 21644 16828 21812 16830
rect 21868 16884 21924 16894
rect 21868 16882 22148 16884
rect 21868 16830 21870 16882
rect 21922 16830 22148 16882
rect 21868 16828 22148 16830
rect 21420 15540 21476 16492
rect 21644 16436 21700 16828
rect 21868 16818 21924 16828
rect 21420 15474 21476 15484
rect 21532 16380 21700 16436
rect 21868 16548 21924 16558
rect 21532 14644 21588 16380
rect 21756 15988 21812 15998
rect 21756 15894 21812 15932
rect 21644 15540 21700 15550
rect 21644 15426 21700 15484
rect 21644 15374 21646 15426
rect 21698 15374 21700 15426
rect 21644 14756 21700 15374
rect 21868 15316 21924 16492
rect 21700 14700 21812 14756
rect 21644 14690 21700 14700
rect 21532 14578 21588 14588
rect 21532 14308 21588 14318
rect 21532 13746 21588 14252
rect 21532 13694 21534 13746
rect 21586 13694 21588 13746
rect 21532 13682 21588 13694
rect 21308 13010 21364 13020
rect 21532 13300 21588 13310
rect 21532 13074 21588 13244
rect 21532 13022 21534 13074
rect 21586 13022 21588 13074
rect 21532 13010 21588 13022
rect 21644 13076 21700 13086
rect 21420 12740 21476 12750
rect 21420 12402 21476 12684
rect 21420 12350 21422 12402
rect 21474 12350 21476 12402
rect 21420 12338 21476 12350
rect 21252 11676 21476 11732
rect 21196 11666 21252 11676
rect 20636 10612 20692 10622
rect 20412 9938 20580 9940
rect 20412 9886 20414 9938
rect 20466 9886 20580 9938
rect 20412 9884 20580 9886
rect 20412 9874 20468 9884
rect 20076 9548 20244 9604
rect 19964 9538 20020 9548
rect 19628 9426 19684 9436
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19964 9268 20020 9278
rect 20188 9268 20244 9548
rect 19516 9212 19796 9268
rect 19404 8988 19572 9044
rect 19180 8866 19236 8876
rect 19068 8754 19124 8764
rect 19516 8708 19572 8988
rect 19628 9042 19684 9054
rect 19628 8990 19630 9042
rect 19682 8990 19684 9042
rect 19628 8932 19684 8990
rect 19628 8866 19684 8876
rect 19404 8652 19572 8708
rect 18620 8206 18622 8258
rect 18674 8206 18676 8258
rect 18620 7700 18676 8206
rect 18620 7634 18676 7644
rect 18956 8596 19012 8606
rect 18844 7364 18900 7374
rect 18732 7250 18788 7262
rect 18732 7198 18734 7250
rect 18786 7198 18788 7250
rect 18732 7140 18788 7198
rect 18732 7074 18788 7084
rect 18732 6916 18788 6926
rect 18732 5796 18788 6860
rect 18844 6020 18900 7308
rect 18956 7252 19012 8540
rect 19292 8372 19348 8382
rect 19292 8260 19348 8316
rect 19068 8258 19348 8260
rect 19068 8206 19294 8258
rect 19346 8206 19348 8258
rect 19068 8204 19348 8206
rect 19068 7476 19124 8204
rect 19292 8194 19348 8204
rect 19292 7476 19348 7486
rect 19068 7474 19236 7476
rect 19068 7422 19070 7474
rect 19122 7422 19236 7474
rect 19068 7420 19236 7422
rect 19068 7410 19124 7420
rect 18956 7196 19124 7252
rect 18956 6580 19012 6590
rect 18956 6466 19012 6524
rect 18956 6414 18958 6466
rect 19010 6414 19012 6466
rect 18956 6402 19012 6414
rect 18844 5964 19012 6020
rect 18844 5796 18900 5806
rect 18732 5794 18900 5796
rect 18732 5742 18846 5794
rect 18898 5742 18900 5794
rect 18732 5740 18900 5742
rect 18844 5730 18900 5740
rect 18844 4564 18900 4574
rect 18396 4562 18900 4564
rect 18396 4510 18398 4562
rect 18450 4510 18846 4562
rect 18898 4510 18900 4562
rect 18396 4508 18900 4510
rect 18396 4498 18452 4508
rect 18844 4498 18900 4508
rect 17948 3938 18004 3948
rect 16884 3612 17556 3668
rect 18732 3892 18788 3902
rect 16828 3536 16884 3612
rect 18732 3554 18788 3836
rect 18956 3778 19012 5964
rect 19068 5234 19124 7196
rect 19180 6916 19236 7420
rect 19292 7382 19348 7420
rect 19292 6916 19348 6926
rect 19180 6914 19348 6916
rect 19180 6862 19294 6914
rect 19346 6862 19348 6914
rect 19180 6860 19348 6862
rect 19292 6132 19348 6860
rect 19404 6468 19460 8652
rect 19740 8596 19796 9212
rect 19740 8530 19796 8540
rect 19516 8484 19572 8494
rect 19516 8034 19572 8428
rect 19516 7982 19518 8034
rect 19570 7982 19572 8034
rect 19516 7970 19572 7982
rect 19740 8372 19796 8382
rect 19740 8036 19796 8316
rect 19964 8372 20020 9212
rect 20076 9212 20244 9268
rect 20076 8428 20132 9212
rect 20412 8596 20468 8606
rect 20076 8372 20244 8428
rect 19964 8306 20020 8316
rect 20076 8036 20132 8046
rect 19740 8034 20132 8036
rect 19740 7982 20078 8034
rect 20130 7982 20132 8034
rect 19740 7980 20132 7982
rect 20076 7970 20132 7980
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19852 7700 19908 7710
rect 19852 7606 19908 7644
rect 20188 7252 20244 8372
rect 20300 8372 20356 8382
rect 20300 7700 20356 8316
rect 20300 7634 20356 7644
rect 20188 7186 20244 7196
rect 20300 7362 20356 7374
rect 20300 7310 20302 7362
rect 20354 7310 20356 7362
rect 19628 7140 19684 7150
rect 19516 6692 19572 6702
rect 19516 6598 19572 6636
rect 19404 6412 19572 6468
rect 19404 6132 19460 6142
rect 19292 6130 19460 6132
rect 19292 6078 19406 6130
rect 19458 6078 19460 6130
rect 19292 6076 19460 6078
rect 19404 6066 19460 6076
rect 19068 5182 19070 5234
rect 19122 5182 19124 5234
rect 19068 5170 19124 5182
rect 19516 5234 19572 6412
rect 19628 6132 19684 7084
rect 20076 6580 20132 6590
rect 20076 6486 20132 6524
rect 20300 6468 20356 7310
rect 20412 6578 20468 8540
rect 20412 6526 20414 6578
rect 20466 6526 20468 6578
rect 20412 6514 20468 6526
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19628 6066 19684 6076
rect 19516 5182 19518 5234
rect 19570 5182 19572 5234
rect 19516 5170 19572 5182
rect 19628 5906 19684 5918
rect 19628 5854 19630 5906
rect 19682 5854 19684 5906
rect 19628 5572 19684 5854
rect 19292 5124 19348 5134
rect 19292 4562 19348 5068
rect 19292 4510 19294 4562
rect 19346 4510 19348 4562
rect 19292 4498 19348 4510
rect 19628 4564 19684 5516
rect 19964 5236 20020 5246
rect 19964 5142 20020 5180
rect 20300 5124 20356 6412
rect 20300 5058 20356 5068
rect 20300 4900 20356 4910
rect 20524 4900 20580 9884
rect 20636 8370 20692 10556
rect 20748 9940 20804 9950
rect 20748 8932 20804 9884
rect 20748 8838 20804 8876
rect 20860 9602 20916 9614
rect 20860 9550 20862 9602
rect 20914 9550 20916 9602
rect 20636 8318 20638 8370
rect 20690 8318 20692 8370
rect 20636 8306 20692 8318
rect 20860 8372 20916 9550
rect 20860 7698 20916 8316
rect 20860 7646 20862 7698
rect 20914 7646 20916 7698
rect 20860 7634 20916 7646
rect 20860 7252 20916 7262
rect 20636 6132 20692 6142
rect 20636 6038 20692 6076
rect 20860 5234 20916 7196
rect 20972 6802 21028 11564
rect 21308 10500 21364 10510
rect 21420 10500 21476 11676
rect 21644 11506 21700 13020
rect 21644 11454 21646 11506
rect 21698 11454 21700 11506
rect 21644 11442 21700 11454
rect 21532 11396 21588 11406
rect 21532 10724 21588 11340
rect 21532 10668 21700 10724
rect 21532 10500 21588 10510
rect 21420 10498 21588 10500
rect 21420 10446 21534 10498
rect 21586 10446 21588 10498
rect 21420 10444 21588 10446
rect 21308 9266 21364 10444
rect 21532 9380 21588 10444
rect 21308 9214 21310 9266
rect 21362 9214 21364 9266
rect 21308 9202 21364 9214
rect 21420 9324 21532 9380
rect 20972 6750 20974 6802
rect 21026 6750 21028 6802
rect 20972 6738 21028 6750
rect 21084 7700 21140 7710
rect 21084 6130 21140 7644
rect 21084 6078 21086 6130
rect 21138 6078 21140 6130
rect 21084 6066 21140 6078
rect 21420 6132 21476 9324
rect 21532 9314 21588 9324
rect 21644 8372 21700 10668
rect 21756 10052 21812 14700
rect 21868 14642 21924 15260
rect 21868 14590 21870 14642
rect 21922 14590 21924 14642
rect 21868 14578 21924 14590
rect 21980 15986 22036 15998
rect 21980 15934 21982 15986
rect 22034 15934 22036 15986
rect 21980 14868 22036 15934
rect 22092 15988 22148 16828
rect 22204 15988 22260 20748
rect 22316 20578 22372 20590
rect 22316 20526 22318 20578
rect 22370 20526 22372 20578
rect 22316 20244 22372 20526
rect 22316 20178 22372 20188
rect 22428 20130 22484 23324
rect 22540 21812 22596 21822
rect 22652 21812 22708 23772
rect 22876 23762 22932 23772
rect 22764 23044 22820 23054
rect 22764 22950 22820 22988
rect 22876 22372 22932 22382
rect 22876 22278 22932 22316
rect 22540 21810 22708 21812
rect 22540 21758 22542 21810
rect 22594 21758 22708 21810
rect 22540 21756 22708 21758
rect 22764 22258 22820 22270
rect 22764 22206 22766 22258
rect 22818 22206 22820 22258
rect 22540 21746 22596 21756
rect 22652 21586 22708 21598
rect 22652 21534 22654 21586
rect 22706 21534 22708 21586
rect 22652 20916 22708 21534
rect 22652 20850 22708 20860
rect 22764 21588 22820 22206
rect 22764 20356 22820 21532
rect 22876 20802 22932 20814
rect 22876 20750 22878 20802
rect 22930 20750 22932 20802
rect 22876 20580 22932 20750
rect 22876 20514 22932 20524
rect 22428 20078 22430 20130
rect 22482 20078 22484 20130
rect 22428 20066 22484 20078
rect 22540 20300 22820 20356
rect 22428 19572 22484 19582
rect 22316 15988 22372 15998
rect 22204 15986 22372 15988
rect 22204 15934 22318 15986
rect 22370 15934 22372 15986
rect 22204 15932 22372 15934
rect 22092 15874 22148 15932
rect 22092 15822 22094 15874
rect 22146 15822 22148 15874
rect 22092 15810 22148 15822
rect 22316 15652 22372 15932
rect 22316 15586 22372 15596
rect 22428 15540 22484 19516
rect 22540 17444 22596 20300
rect 22652 20132 22708 20142
rect 22988 20132 23044 25564
rect 23212 25554 23268 25564
rect 23324 25956 23380 25966
rect 23100 25394 23156 25406
rect 23100 25342 23102 25394
rect 23154 25342 23156 25394
rect 23100 25172 23156 25342
rect 23212 25396 23268 25406
rect 23212 25302 23268 25340
rect 23100 25106 23156 25116
rect 23100 24836 23156 24846
rect 23100 23380 23156 24780
rect 23212 23940 23268 23950
rect 23212 23846 23268 23884
rect 23212 23380 23268 23390
rect 23100 23378 23268 23380
rect 23100 23326 23214 23378
rect 23266 23326 23268 23378
rect 23100 23324 23268 23326
rect 23212 23314 23268 23324
rect 23212 23044 23268 23054
rect 23100 21028 23156 21038
rect 23100 20934 23156 20972
rect 22652 18340 22708 20076
rect 22876 20076 23044 20132
rect 22764 19796 22820 19806
rect 22764 19702 22820 19740
rect 22876 19348 22932 20076
rect 22988 19906 23044 19918
rect 22988 19854 22990 19906
rect 23042 19854 23044 19906
rect 22988 19572 23044 19854
rect 22988 19506 23044 19516
rect 22988 19348 23044 19358
rect 22876 19346 23044 19348
rect 22876 19294 22990 19346
rect 23042 19294 23044 19346
rect 22876 19292 23044 19294
rect 22988 19282 23044 19292
rect 22876 19012 22932 19022
rect 23100 19012 23156 19022
rect 22876 19010 23044 19012
rect 22876 18958 22878 19010
rect 22930 18958 23044 19010
rect 22876 18956 23044 18958
rect 22876 18946 22932 18956
rect 22876 18340 22932 18350
rect 22652 18338 22932 18340
rect 22652 18286 22878 18338
rect 22930 18286 22932 18338
rect 22652 18284 22932 18286
rect 22876 18274 22932 18284
rect 22988 18340 23044 18956
rect 23100 18918 23156 18956
rect 23212 18788 23268 22988
rect 23324 21924 23380 25900
rect 23436 25508 23492 26348
rect 23436 25376 23492 25452
rect 23548 26402 23604 26414
rect 23548 26350 23550 26402
rect 23602 26350 23604 26402
rect 23548 24724 23604 26350
rect 23548 24658 23604 24668
rect 23660 25394 23716 25406
rect 23660 25342 23662 25394
rect 23714 25342 23716 25394
rect 23660 24500 23716 25342
rect 23660 24434 23716 24444
rect 23772 24052 23828 26852
rect 23996 25060 24052 27020
rect 24108 26852 24164 28028
rect 24108 26516 24164 26796
rect 24108 26450 24164 26460
rect 24332 27074 24388 27086
rect 24332 27022 24334 27074
rect 24386 27022 24388 27074
rect 24332 26404 24388 27022
rect 24332 26338 24388 26348
rect 24220 26290 24276 26302
rect 24220 26238 24222 26290
rect 24274 26238 24276 26290
rect 24220 26068 24276 26238
rect 24444 26068 24500 29932
rect 24556 29428 24612 29438
rect 24556 28868 24612 29372
rect 24780 29428 24836 30156
rect 24668 28868 24724 28878
rect 24556 28866 24724 28868
rect 24556 28814 24670 28866
rect 24722 28814 24724 28866
rect 24556 28812 24724 28814
rect 24668 28802 24724 28812
rect 24780 28754 24836 29372
rect 24780 28702 24782 28754
rect 24834 28702 24836 28754
rect 24780 28690 24836 28702
rect 24892 29316 24948 29326
rect 24668 28644 24724 28654
rect 24668 28082 24724 28588
rect 24892 28530 24948 29260
rect 24892 28478 24894 28530
rect 24946 28478 24948 28530
rect 24892 28466 24948 28478
rect 24668 28030 24670 28082
rect 24722 28030 24724 28082
rect 24556 27860 24612 27870
rect 24556 27766 24612 27804
rect 24220 26002 24276 26012
rect 24332 26012 24500 26068
rect 24556 26850 24612 26862
rect 24556 26798 24558 26850
rect 24610 26798 24612 26850
rect 24332 25618 24388 26012
rect 24332 25566 24334 25618
rect 24386 25566 24388 25618
rect 24332 25554 24388 25566
rect 24444 25508 24500 25518
rect 24556 25508 24612 26798
rect 24444 25506 24612 25508
rect 24444 25454 24446 25506
rect 24498 25454 24612 25506
rect 24444 25452 24612 25454
rect 24444 25442 24500 25452
rect 24220 25284 24276 25294
rect 24220 25190 24276 25228
rect 23996 25004 24500 25060
rect 24332 24836 24388 24846
rect 24332 24742 24388 24780
rect 23660 23996 23828 24052
rect 23996 24722 24052 24734
rect 23996 24670 23998 24722
rect 24050 24670 24052 24722
rect 23548 23828 23604 23838
rect 23436 23268 23492 23278
rect 23436 21924 23492 23212
rect 23548 22258 23604 23772
rect 23660 23604 23716 23996
rect 23772 23828 23828 23838
rect 23772 23734 23828 23772
rect 23660 23548 23828 23604
rect 23548 22206 23550 22258
rect 23602 22206 23604 22258
rect 23548 22194 23604 22206
rect 23660 23154 23716 23166
rect 23660 23102 23662 23154
rect 23714 23102 23716 23154
rect 23660 22036 23716 23102
rect 23660 21970 23716 21980
rect 23436 21868 23604 21924
rect 23324 21858 23380 21868
rect 23436 21698 23492 21710
rect 23436 21646 23438 21698
rect 23490 21646 23492 21698
rect 23324 21588 23380 21598
rect 23324 21494 23380 21532
rect 23324 20804 23380 20814
rect 23436 20804 23492 21646
rect 23324 20802 23492 20804
rect 23324 20750 23326 20802
rect 23378 20750 23492 20802
rect 23324 20748 23492 20750
rect 23324 20692 23380 20748
rect 23324 20626 23380 20636
rect 23548 20244 23604 21868
rect 23660 21700 23716 21710
rect 23660 21606 23716 21644
rect 23772 21026 23828 23548
rect 23996 22708 24052 24670
rect 24332 24500 24388 24510
rect 24108 24050 24164 24062
rect 24108 23998 24110 24050
rect 24162 23998 24164 24050
rect 24108 23940 24164 23998
rect 24108 23874 24164 23884
rect 24220 23938 24276 23950
rect 24220 23886 24222 23938
rect 24274 23886 24276 23938
rect 24220 23044 24276 23886
rect 24220 22950 24276 22988
rect 23996 22652 24164 22708
rect 24108 22260 24164 22652
rect 23996 22204 24164 22260
rect 23772 20974 23774 21026
rect 23826 20974 23828 21026
rect 23772 20962 23828 20974
rect 23884 22146 23940 22158
rect 23884 22094 23886 22146
rect 23938 22094 23940 22146
rect 23884 21812 23940 22094
rect 23884 20356 23940 21756
rect 23884 20290 23940 20300
rect 23996 21474 24052 22204
rect 23996 21422 23998 21474
rect 24050 21422 24052 21474
rect 23660 20244 23716 20254
rect 23548 20242 23716 20244
rect 23548 20190 23662 20242
rect 23714 20190 23716 20242
rect 23548 20188 23716 20190
rect 23660 20178 23716 20188
rect 23772 20132 23828 20142
rect 23772 20038 23828 20076
rect 23548 20018 23604 20030
rect 23548 19966 23550 20018
rect 23602 19966 23604 20018
rect 23548 19796 23604 19966
rect 23996 19908 24052 21422
rect 23436 19740 23548 19796
rect 23324 19236 23380 19246
rect 23324 19142 23380 19180
rect 22988 18274 23044 18284
rect 23100 18732 23268 18788
rect 22764 17892 22820 17902
rect 22540 17350 22596 17388
rect 22652 17780 22708 17790
rect 22652 17220 22708 17724
rect 22428 15408 22484 15484
rect 22540 17164 22708 17220
rect 22204 15204 22260 15214
rect 22204 15092 22372 15148
rect 21980 14532 22036 14812
rect 21980 14476 22260 14532
rect 22092 14308 22148 14318
rect 21980 12964 22036 12974
rect 21868 12292 21924 12302
rect 21868 12198 21924 12236
rect 21980 11956 22036 12908
rect 22092 12962 22148 14252
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 22092 12898 22148 12910
rect 22204 12740 22260 14476
rect 22092 12684 22260 12740
rect 22316 13074 22372 15092
rect 22428 14420 22484 14430
rect 22428 14306 22484 14364
rect 22428 14254 22430 14306
rect 22482 14254 22484 14306
rect 22428 13748 22484 14254
rect 22540 13972 22596 17164
rect 22652 16996 22708 17006
rect 22652 16882 22708 16940
rect 22652 16830 22654 16882
rect 22706 16830 22708 16882
rect 22652 16818 22708 16830
rect 22652 13972 22708 13982
rect 22540 13970 22708 13972
rect 22540 13918 22654 13970
rect 22706 13918 22708 13970
rect 22540 13916 22708 13918
rect 22652 13906 22708 13916
rect 22428 13682 22484 13692
rect 22540 13412 22596 13422
rect 22428 13300 22484 13310
rect 22428 13186 22484 13244
rect 22428 13134 22430 13186
rect 22482 13134 22484 13186
rect 22428 13122 22484 13134
rect 22316 13022 22318 13074
rect 22370 13022 22372 13074
rect 22092 12290 22148 12684
rect 22316 12404 22372 13022
rect 22316 12348 22484 12404
rect 22092 12238 22094 12290
rect 22146 12238 22148 12290
rect 22092 12180 22148 12238
rect 22204 12292 22260 12302
rect 22204 12198 22260 12236
rect 22092 12114 22148 12124
rect 21756 9996 21924 10052
rect 21756 9828 21812 9838
rect 21756 9266 21812 9772
rect 21756 9214 21758 9266
rect 21810 9214 21812 9266
rect 21756 9202 21812 9214
rect 21868 9268 21924 9996
rect 21868 9202 21924 9212
rect 21980 8596 22036 11900
rect 22092 11732 22148 11742
rect 22092 11172 22148 11676
rect 22092 11078 22148 11116
rect 22204 10836 22260 10846
rect 22204 10722 22260 10780
rect 22204 10670 22206 10722
rect 22258 10670 22260 10722
rect 22204 10658 22260 10670
rect 22092 10612 22148 10622
rect 22092 9940 22148 10556
rect 22204 9940 22260 9950
rect 22092 9938 22260 9940
rect 22092 9886 22206 9938
rect 22258 9886 22260 9938
rect 22092 9884 22260 9886
rect 22204 9874 22260 9884
rect 22316 9826 22372 9838
rect 22316 9774 22318 9826
rect 22370 9774 22372 9826
rect 22316 9492 22372 9774
rect 22316 9426 22372 9436
rect 22428 9156 22484 12348
rect 22540 10498 22596 13356
rect 22540 10446 22542 10498
rect 22594 10446 22596 10498
rect 22540 10434 22596 10446
rect 22652 11282 22708 11294
rect 22652 11230 22654 11282
rect 22706 11230 22708 11282
rect 22652 11172 22708 11230
rect 22540 9828 22596 9838
rect 22540 9734 22596 9772
rect 22540 9268 22596 9278
rect 22540 9174 22596 9212
rect 22316 9100 22484 9156
rect 21980 8530 22036 8540
rect 22092 9042 22148 9054
rect 22092 8990 22094 9042
rect 22146 8990 22148 9042
rect 21756 8372 21812 8382
rect 21644 8370 21812 8372
rect 21644 8318 21758 8370
rect 21810 8318 21812 8370
rect 21644 8316 21812 8318
rect 21756 8306 21812 8316
rect 22092 8372 22148 8990
rect 22092 8306 22148 8316
rect 21420 6066 21476 6076
rect 21532 8260 21588 8270
rect 20860 5182 20862 5234
rect 20914 5182 20916 5234
rect 20860 5170 20916 5182
rect 21532 5234 21588 8204
rect 22204 8148 22260 8158
rect 22204 8034 22260 8092
rect 22204 7982 22206 8034
rect 22258 7982 22260 8034
rect 21868 7586 21924 7598
rect 21868 7534 21870 7586
rect 21922 7534 21924 7586
rect 21644 7476 21700 7486
rect 21868 7476 21924 7534
rect 21644 7474 21812 7476
rect 21644 7422 21646 7474
rect 21698 7422 21812 7474
rect 21644 7420 21812 7422
rect 21644 7410 21700 7420
rect 21756 6804 21812 7420
rect 21868 7410 21924 7420
rect 22204 7476 22260 7982
rect 22204 7410 22260 7420
rect 22316 7140 22372 9100
rect 22316 7074 22372 7084
rect 22428 8932 22484 8942
rect 22652 8932 22708 11116
rect 22764 11060 22820 17836
rect 23100 17332 23156 18732
rect 23436 18676 23492 19740
rect 23548 19664 23604 19740
rect 23772 19852 24052 19908
rect 24108 21924 24164 21934
rect 23548 19348 23604 19358
rect 23548 19254 23604 19292
rect 23436 18610 23492 18620
rect 23548 18452 23604 18462
rect 23492 18450 23604 18452
rect 23492 18398 23550 18450
rect 23602 18398 23604 18450
rect 23492 18386 23604 18398
rect 23772 18452 23828 19852
rect 23996 19458 24052 19470
rect 23996 19406 23998 19458
rect 24050 19406 24052 19458
rect 23996 18788 24052 19406
rect 23996 18674 24052 18732
rect 23996 18622 23998 18674
rect 24050 18622 24052 18674
rect 23996 18610 24052 18622
rect 24108 18674 24164 21868
rect 24332 21252 24388 24444
rect 24444 21812 24500 25004
rect 24444 21746 24500 21756
rect 24444 21588 24500 21598
rect 24444 21494 24500 21532
rect 24332 21196 24500 21252
rect 24332 20804 24388 20814
rect 24220 20802 24388 20804
rect 24220 20750 24334 20802
rect 24386 20750 24388 20802
rect 24220 20748 24388 20750
rect 24220 19458 24276 20748
rect 24332 20738 24388 20748
rect 24444 20580 24500 21196
rect 24668 21140 24724 28030
rect 24892 28084 24948 28094
rect 25004 28084 25060 36204
rect 25116 36194 25172 36204
rect 25116 34690 25172 34702
rect 25116 34638 25118 34690
rect 25170 34638 25172 34690
rect 25116 33572 25172 34638
rect 25116 33506 25172 33516
rect 25340 32004 25396 32014
rect 25340 30322 25396 31948
rect 25340 30270 25342 30322
rect 25394 30270 25396 30322
rect 24892 28082 25060 28084
rect 24892 28030 24894 28082
rect 24946 28030 25060 28082
rect 24892 28028 25060 28030
rect 25116 28980 25172 28990
rect 24892 28018 24948 28028
rect 25004 27748 25060 27758
rect 24780 27300 24836 27310
rect 24780 27074 24836 27244
rect 24780 27022 24782 27074
rect 24834 27022 24836 27074
rect 24780 27010 24836 27022
rect 24892 27188 24948 27198
rect 24892 26908 24948 27132
rect 25004 27074 25060 27692
rect 25004 27022 25006 27074
rect 25058 27022 25060 27074
rect 25004 27010 25060 27022
rect 24780 26852 24948 26908
rect 24780 25506 24836 26852
rect 25116 26516 25172 28924
rect 25116 26450 25172 26460
rect 25228 28420 25284 28430
rect 24892 26292 24948 26302
rect 24892 26180 24948 26236
rect 25228 26180 25284 28364
rect 25340 28196 25396 30270
rect 25340 28130 25396 28140
rect 24892 26178 25284 26180
rect 24892 26126 24894 26178
rect 24946 26126 25284 26178
rect 24892 26124 25284 26126
rect 25340 27748 25396 27758
rect 24892 26114 24948 26124
rect 24780 25454 24782 25506
rect 24834 25454 24836 25506
rect 24780 25442 24836 25454
rect 24892 25732 24948 25742
rect 24892 25284 24948 25676
rect 24892 24610 24948 25228
rect 24892 24558 24894 24610
rect 24946 24558 24948 24610
rect 24780 23940 24836 23950
rect 24780 23846 24836 23884
rect 24892 23156 24948 24558
rect 25004 23378 25060 26124
rect 25004 23326 25006 23378
rect 25058 23326 25060 23378
rect 25004 23314 25060 23326
rect 25228 25284 25284 25294
rect 24892 23090 24948 23100
rect 24892 21476 24948 21486
rect 24892 21382 24948 21420
rect 24668 21084 25060 21140
rect 24668 20914 24724 20926
rect 24668 20862 24670 20914
rect 24722 20862 24724 20914
rect 24668 20692 24724 20862
rect 24668 20626 24724 20636
rect 24556 20580 24612 20590
rect 24444 20578 24612 20580
rect 24444 20526 24558 20578
rect 24610 20526 24612 20578
rect 24444 20524 24612 20526
rect 24444 20244 24500 20254
rect 24332 20130 24388 20142
rect 24332 20078 24334 20130
rect 24386 20078 24388 20130
rect 24332 20020 24388 20078
rect 24332 19572 24388 19964
rect 24332 19506 24388 19516
rect 24220 19406 24222 19458
rect 24274 19406 24276 19458
rect 24220 19394 24276 19406
rect 24332 19236 24388 19246
rect 24220 19012 24276 19022
rect 24220 18918 24276 18956
rect 24108 18622 24110 18674
rect 24162 18622 24164 18674
rect 24108 18610 24164 18622
rect 24220 18564 24276 18574
rect 24220 18470 24276 18508
rect 23772 18386 23828 18396
rect 23884 18450 23940 18462
rect 23884 18398 23886 18450
rect 23938 18398 23940 18450
rect 23492 18350 23548 18386
rect 23436 18340 23548 18350
rect 23492 18284 23548 18340
rect 23324 18226 23380 18238
rect 23324 18174 23326 18226
rect 23378 18174 23380 18226
rect 23324 17892 23380 18174
rect 23324 17826 23380 17836
rect 23436 17780 23492 18284
rect 23884 17892 23940 18398
rect 24332 18004 24388 19180
rect 24444 18788 24500 20188
rect 24556 19796 24612 20524
rect 24892 20356 24948 20366
rect 24556 19730 24612 19740
rect 24668 20132 24724 20142
rect 24444 18732 24612 18788
rect 23436 17714 23492 17724
rect 23772 17836 23884 17892
rect 23324 17668 23380 17678
rect 23324 17574 23380 17612
rect 23212 17556 23268 17566
rect 23212 17462 23268 17500
rect 23436 17554 23492 17566
rect 23436 17502 23438 17554
rect 23490 17502 23492 17554
rect 23324 17444 23380 17454
rect 23436 17444 23492 17502
rect 23380 17388 23492 17444
rect 23100 17276 23268 17332
rect 23100 16882 23156 16894
rect 23100 16830 23102 16882
rect 23154 16830 23156 16882
rect 23100 16212 23156 16830
rect 23212 16436 23268 17276
rect 23212 16370 23268 16380
rect 23212 16212 23268 16222
rect 23100 16210 23268 16212
rect 23100 16158 23214 16210
rect 23266 16158 23268 16210
rect 23100 16156 23268 16158
rect 23212 16146 23268 16156
rect 23324 16100 23380 17388
rect 23660 16884 23716 16894
rect 23660 16770 23716 16828
rect 23772 16882 23828 17836
rect 23884 17826 23940 17836
rect 23996 17948 24388 18004
rect 24444 18228 24500 18238
rect 23772 16830 23774 16882
rect 23826 16830 23828 16882
rect 23772 16818 23828 16830
rect 23884 17668 23940 17678
rect 23996 17668 24052 17948
rect 24444 17778 24500 18172
rect 24444 17726 24446 17778
rect 24498 17726 24500 17778
rect 24444 17714 24500 17726
rect 23884 17666 24052 17668
rect 23884 17614 23886 17666
rect 23938 17614 24052 17666
rect 23884 17612 24052 17614
rect 23660 16718 23662 16770
rect 23714 16718 23716 16770
rect 23660 16706 23716 16718
rect 23436 16660 23492 16670
rect 23436 16566 23492 16604
rect 23884 16548 23940 17612
rect 23548 16492 23940 16548
rect 23996 16548 24052 16558
rect 23548 16436 23604 16492
rect 23996 16436 24052 16492
rect 24556 16548 24612 18732
rect 24556 16482 24612 16492
rect 23324 16034 23380 16044
rect 23436 16380 23604 16436
rect 23772 16380 24052 16436
rect 23436 16098 23492 16380
rect 23772 16322 23828 16380
rect 23772 16270 23774 16322
rect 23826 16270 23828 16322
rect 23772 16258 23828 16270
rect 23436 16046 23438 16098
rect 23490 16046 23492 16098
rect 23436 16034 23492 16046
rect 23548 16100 23604 16110
rect 22988 15988 23044 15998
rect 23044 15932 23156 15988
rect 22988 15922 23044 15932
rect 23100 15874 23156 15932
rect 23100 15822 23102 15874
rect 23154 15822 23156 15874
rect 23100 15810 23156 15822
rect 23324 15874 23380 15886
rect 23324 15822 23326 15874
rect 23378 15822 23380 15874
rect 23324 15764 23380 15822
rect 23324 15698 23380 15708
rect 22988 15540 23044 15550
rect 23548 15540 23604 16044
rect 23772 15540 23828 15550
rect 22988 15446 23044 15484
rect 23436 15538 23828 15540
rect 23436 15486 23774 15538
rect 23826 15486 23828 15538
rect 23436 15484 23828 15486
rect 23324 15314 23380 15326
rect 23324 15262 23326 15314
rect 23378 15262 23380 15314
rect 23324 15204 23380 15262
rect 23324 15138 23380 15148
rect 23436 15148 23492 15484
rect 23772 15474 23828 15484
rect 23884 15428 23940 16380
rect 23884 15362 23940 15372
rect 24220 16324 24276 16334
rect 24220 15764 24276 16268
rect 24556 16100 24612 16110
rect 24556 16006 24612 16044
rect 23660 15204 23716 15214
rect 23436 15092 23604 15148
rect 23100 14644 23156 14654
rect 23100 14550 23156 14588
rect 23324 14418 23380 14430
rect 23324 14366 23326 14418
rect 23378 14366 23380 14418
rect 22988 14306 23044 14318
rect 22988 14254 22990 14306
rect 23042 14254 23044 14306
rect 22988 14084 23044 14254
rect 23212 14308 23268 14318
rect 23212 14214 23268 14252
rect 23324 14196 23380 14366
rect 23324 14130 23380 14140
rect 22988 14018 23044 14028
rect 23436 14084 23492 14094
rect 23436 13858 23492 14028
rect 23436 13806 23438 13858
rect 23490 13806 23492 13858
rect 22876 13300 22932 13310
rect 22876 12402 22932 13244
rect 23436 13300 23492 13806
rect 23436 13234 23492 13244
rect 22988 13188 23044 13198
rect 22988 13074 23044 13132
rect 22988 13022 22990 13074
rect 23042 13022 23044 13074
rect 22988 13010 23044 13022
rect 22876 12350 22878 12402
rect 22930 12350 22932 12402
rect 22876 12292 22932 12350
rect 22876 12226 22932 12236
rect 23100 12740 23156 12750
rect 23100 11396 23156 12684
rect 23548 12404 23604 15092
rect 23660 12850 23716 15148
rect 23772 14532 23828 14542
rect 23772 14530 24164 14532
rect 23772 14478 23774 14530
rect 23826 14478 24164 14530
rect 23772 14476 24164 14478
rect 23772 14466 23828 14476
rect 23660 12798 23662 12850
rect 23714 12798 23716 12850
rect 23660 12786 23716 12798
rect 23772 13746 23828 13758
rect 23772 13694 23774 13746
rect 23826 13694 23828 13746
rect 23772 12852 23828 13694
rect 24108 13746 24164 14476
rect 24220 13970 24276 15708
rect 24556 15540 24612 15550
rect 24556 15446 24612 15484
rect 24668 14418 24724 20076
rect 24780 19348 24836 19358
rect 24780 16772 24836 19292
rect 24892 19346 24948 20300
rect 24892 19294 24894 19346
rect 24946 19294 24948 19346
rect 24892 19282 24948 19294
rect 24892 18788 24948 18798
rect 24892 18674 24948 18732
rect 24892 18622 24894 18674
rect 24946 18622 24948 18674
rect 24892 16996 24948 18622
rect 25004 17666 25060 21084
rect 25116 20802 25172 20814
rect 25116 20750 25118 20802
rect 25170 20750 25172 20802
rect 25116 20692 25172 20750
rect 25116 20626 25172 20636
rect 25004 17614 25006 17666
rect 25058 17614 25060 17666
rect 25004 17556 25060 17614
rect 25004 17490 25060 17500
rect 25116 17668 25172 17678
rect 25116 17554 25172 17612
rect 25116 17502 25118 17554
rect 25170 17502 25172 17554
rect 25116 17444 25172 17502
rect 24892 16940 25060 16996
rect 24892 16772 24948 16782
rect 24836 16770 24948 16772
rect 24836 16718 24894 16770
rect 24946 16718 24948 16770
rect 24836 16716 24948 16718
rect 24780 16706 24836 16716
rect 24892 16706 24948 16716
rect 24780 16548 24836 16558
rect 25004 16548 25060 16940
rect 25116 16772 25172 17388
rect 25228 16884 25284 25228
rect 25340 25060 25396 27692
rect 25452 27634 25508 37998
rect 25788 37828 25844 38894
rect 25900 38834 25956 38846
rect 25900 38782 25902 38834
rect 25954 38782 25956 38834
rect 25900 38276 25956 38782
rect 26012 38722 26068 40124
rect 26012 38670 26014 38722
rect 26066 38670 26068 38722
rect 26012 38658 26068 38670
rect 26348 38724 26404 38734
rect 26684 38668 26740 41132
rect 27804 41188 27860 41198
rect 27804 41094 27860 41132
rect 27356 41076 27412 41086
rect 27356 40982 27412 41020
rect 27244 40964 27300 40974
rect 27244 40870 27300 40908
rect 26796 40628 26852 40638
rect 26796 40514 26852 40572
rect 26796 40462 26798 40514
rect 26850 40462 26852 40514
rect 26796 40450 26852 40462
rect 27468 40404 27524 40414
rect 27468 40310 27524 40348
rect 28364 40404 28420 40414
rect 28364 40310 28420 40348
rect 27692 40292 27748 40302
rect 27692 40198 27748 40236
rect 27916 39396 27972 39406
rect 25900 38210 25956 38220
rect 25900 38052 25956 38062
rect 25900 37958 25956 37996
rect 25564 37772 25844 37828
rect 25564 37490 25620 37772
rect 26348 37492 26404 38668
rect 25564 37438 25566 37490
rect 25618 37438 25620 37490
rect 25564 37426 25620 37438
rect 25900 37490 26404 37492
rect 25900 37438 26350 37490
rect 26402 37438 26404 37490
rect 25900 37436 26404 37438
rect 25788 37380 25844 37390
rect 25788 37286 25844 37324
rect 25900 37378 25956 37436
rect 26348 37426 26404 37436
rect 26460 38612 26740 38668
rect 26908 38834 26964 38846
rect 26908 38782 26910 38834
rect 26962 38782 26964 38834
rect 25900 37326 25902 37378
rect 25954 37326 25956 37378
rect 25900 37314 25956 37326
rect 25676 36260 25732 36270
rect 25676 36166 25732 36204
rect 26012 36260 26068 36270
rect 26012 36166 26068 36204
rect 26460 35812 26516 38612
rect 26908 38052 26964 38782
rect 27020 38724 27076 38762
rect 27020 38658 27076 38668
rect 27804 38722 27860 38734
rect 27804 38670 27806 38722
rect 27858 38670 27860 38722
rect 27804 38612 27860 38670
rect 27804 38546 27860 38556
rect 26908 37986 26964 37996
rect 27804 38050 27860 38062
rect 27804 37998 27806 38050
rect 27858 37998 27860 38050
rect 27692 37940 27748 37950
rect 27132 37938 27748 37940
rect 27132 37886 27694 37938
rect 27746 37886 27748 37938
rect 27132 37884 27748 37886
rect 27132 36482 27188 37884
rect 27692 37874 27748 37884
rect 27804 37604 27860 37998
rect 27468 37548 27860 37604
rect 27356 37492 27412 37502
rect 27356 37398 27412 37436
rect 27468 37490 27524 37548
rect 27468 37438 27470 37490
rect 27522 37438 27524 37490
rect 27468 37426 27524 37438
rect 27580 37380 27636 37390
rect 27916 37380 27972 39340
rect 28140 38948 28196 38958
rect 27580 37378 27972 37380
rect 27580 37326 27582 37378
rect 27634 37326 27972 37378
rect 27580 37324 27972 37326
rect 28028 37380 28084 37390
rect 27580 37314 27636 37324
rect 28028 37286 28084 37324
rect 27132 36430 27134 36482
rect 27186 36430 27188 36482
rect 27132 36418 27188 36430
rect 26012 35756 26516 35812
rect 26684 36260 26740 36270
rect 25564 35586 25620 35598
rect 25564 35534 25566 35586
rect 25618 35534 25620 35586
rect 25564 34916 25620 35534
rect 25564 34850 25620 34860
rect 25900 34130 25956 34142
rect 25900 34078 25902 34130
rect 25954 34078 25956 34130
rect 25788 32788 25844 32798
rect 25900 32788 25956 34078
rect 26012 33796 26068 35756
rect 26124 35586 26180 35598
rect 26124 35534 26126 35586
rect 26178 35534 26180 35586
rect 26124 34132 26180 35534
rect 26348 34244 26404 34254
rect 26348 34150 26404 34188
rect 26124 34066 26180 34076
rect 26572 34130 26628 34142
rect 26572 34078 26574 34130
rect 26626 34078 26628 34130
rect 26460 34018 26516 34030
rect 26460 33966 26462 34018
rect 26514 33966 26516 34018
rect 26012 33740 26180 33796
rect 25788 32786 25956 32788
rect 25788 32734 25790 32786
rect 25842 32734 25956 32786
rect 25788 32732 25956 32734
rect 26012 33012 26068 33022
rect 26012 32786 26068 32956
rect 26012 32734 26014 32786
rect 26066 32734 26068 32786
rect 25788 32722 25844 32732
rect 26012 32722 26068 32734
rect 26124 32788 26180 33740
rect 26124 32732 26292 32788
rect 26124 32564 26180 32574
rect 26124 32470 26180 32508
rect 26236 32340 26292 32732
rect 26124 32284 26292 32340
rect 26012 32004 26068 32014
rect 26012 31218 26068 31948
rect 26012 31166 26014 31218
rect 26066 31166 26068 31218
rect 26012 31154 26068 31166
rect 26124 31218 26180 32284
rect 26460 31666 26516 33966
rect 26572 33348 26628 34078
rect 26572 33012 26628 33292
rect 26572 32946 26628 32956
rect 26684 32788 26740 36204
rect 26796 36258 26852 36270
rect 26796 36206 26798 36258
rect 26850 36206 26852 36258
rect 26796 35924 26852 36206
rect 26796 35858 26852 35868
rect 27356 35812 27412 35822
rect 27356 34914 27412 35756
rect 27356 34862 27358 34914
rect 27410 34862 27412 34914
rect 27356 34850 27412 34862
rect 27468 35700 27524 35710
rect 27020 34244 27076 34254
rect 27020 34150 27076 34188
rect 26908 33572 26964 33582
rect 26908 33478 26964 33516
rect 27020 33460 27076 33470
rect 26460 31614 26462 31666
rect 26514 31614 26516 31666
rect 26460 31602 26516 31614
rect 26572 32732 26740 32788
rect 26908 32788 26964 32798
rect 27020 32788 27076 33404
rect 27356 33460 27412 33470
rect 27356 33366 27412 33404
rect 26908 32786 27076 32788
rect 26908 32734 26910 32786
rect 26962 32734 27076 32786
rect 26908 32732 27076 32734
rect 26124 31166 26126 31218
rect 26178 31166 26180 31218
rect 26124 31154 26180 31166
rect 26236 31108 26292 31118
rect 25564 30996 25620 31006
rect 25564 30902 25620 30940
rect 26236 30212 26292 31052
rect 26124 30156 26292 30212
rect 25900 29986 25956 29998
rect 25900 29934 25902 29986
rect 25954 29934 25956 29986
rect 25900 29652 25956 29934
rect 25900 29586 25956 29596
rect 26124 29650 26180 30156
rect 26124 29598 26126 29650
rect 26178 29598 26180 29650
rect 26124 29586 26180 29598
rect 26236 29986 26292 29998
rect 26236 29934 26238 29986
rect 26290 29934 26292 29986
rect 26236 29652 26292 29934
rect 26236 29558 26292 29596
rect 25564 29428 25620 29438
rect 25564 29334 25620 29372
rect 26012 29428 26068 29438
rect 26012 29334 26068 29372
rect 26348 28532 26404 28542
rect 26236 28476 26348 28532
rect 25900 28420 25956 28430
rect 25900 28326 25956 28364
rect 25900 28196 25956 28206
rect 25452 27582 25454 27634
rect 25506 27582 25508 27634
rect 25452 27570 25508 27582
rect 25564 27746 25620 27758
rect 25564 27694 25566 27746
rect 25618 27694 25620 27746
rect 25452 26964 25508 26974
rect 25452 25730 25508 26908
rect 25564 26908 25620 27694
rect 25676 27412 25732 27422
rect 25900 27412 25956 28140
rect 26124 27972 26180 27982
rect 26012 27970 26180 27972
rect 26012 27918 26126 27970
rect 26178 27918 26180 27970
rect 26012 27916 26180 27918
rect 26012 27634 26068 27916
rect 26124 27906 26180 27916
rect 26012 27582 26014 27634
rect 26066 27582 26068 27634
rect 26012 27570 26068 27582
rect 26236 27412 26292 28476
rect 26348 28438 26404 28476
rect 26460 28420 26516 28430
rect 26460 27858 26516 28364
rect 26460 27806 26462 27858
rect 26514 27806 26516 27858
rect 26460 27794 26516 27806
rect 26460 27636 26516 27646
rect 25900 27356 26068 27412
rect 26236 27356 26404 27412
rect 25676 27186 25732 27356
rect 25676 27134 25678 27186
rect 25730 27134 25732 27186
rect 25676 27122 25732 27134
rect 25900 27076 25956 27086
rect 25564 26852 25844 26908
rect 25676 26292 25732 26302
rect 25676 26198 25732 26236
rect 25452 25678 25454 25730
rect 25506 25678 25508 25730
rect 25452 25666 25508 25678
rect 25564 25396 25620 25406
rect 25564 25302 25620 25340
rect 25452 25282 25508 25294
rect 25452 25230 25454 25282
rect 25506 25230 25508 25282
rect 25452 25172 25508 25230
rect 25452 25116 25620 25172
rect 25340 25004 25508 25060
rect 25340 24276 25396 24286
rect 25340 23938 25396 24220
rect 25340 23886 25342 23938
rect 25394 23886 25396 23938
rect 25340 23828 25396 23886
rect 25452 23938 25508 25004
rect 25564 24836 25620 25116
rect 25564 24770 25620 24780
rect 25452 23886 25454 23938
rect 25506 23886 25508 23938
rect 25452 23874 25508 23886
rect 25788 24722 25844 26796
rect 25900 26514 25956 27020
rect 26012 26908 26068 27356
rect 26124 27188 26180 27198
rect 26124 27074 26180 27132
rect 26124 27022 26126 27074
rect 26178 27022 26180 27074
rect 26124 27010 26180 27022
rect 26348 26908 26404 27356
rect 26460 27076 26516 27580
rect 26572 27186 26628 32732
rect 26908 32722 26964 32732
rect 27356 32676 27412 32686
rect 26684 32562 26740 32574
rect 26684 32510 26686 32562
rect 26738 32510 26740 32562
rect 26684 32004 26740 32510
rect 26796 32564 26852 32574
rect 26796 32470 26852 32508
rect 27356 32562 27412 32620
rect 27356 32510 27358 32562
rect 27410 32510 27412 32562
rect 26684 31938 26740 31948
rect 27020 31444 27076 31454
rect 26796 30884 26852 30894
rect 26684 29428 26740 29438
rect 26684 28644 26740 29372
rect 26796 28868 26852 30828
rect 26796 28812 26964 28868
rect 26684 28512 26740 28588
rect 26908 28420 26964 28812
rect 26572 27134 26574 27186
rect 26626 27134 26628 27186
rect 26572 27122 26628 27134
rect 26684 28364 26964 28420
rect 26460 27010 26516 27020
rect 26572 26964 26628 27002
rect 26012 26852 26180 26908
rect 26348 26852 26516 26908
rect 26572 26898 26628 26908
rect 25900 26462 25902 26514
rect 25954 26462 25956 26514
rect 25900 26450 25956 26462
rect 25900 26290 25956 26302
rect 25900 26238 25902 26290
rect 25954 26238 25956 26290
rect 25900 25732 25956 26238
rect 25900 25666 25956 25676
rect 26012 25396 26068 25406
rect 26012 25302 26068 25340
rect 26012 24836 26068 24846
rect 26012 24742 26068 24780
rect 25788 24670 25790 24722
rect 25842 24670 25844 24722
rect 25788 24276 25844 24670
rect 26124 24500 26180 26852
rect 26236 26404 26292 26414
rect 26236 26290 26292 26348
rect 26236 26238 26238 26290
rect 26290 26238 26292 26290
rect 26236 26180 26292 26238
rect 26236 26114 26292 26124
rect 26348 26292 26404 26302
rect 26124 24434 26180 24444
rect 26236 25620 26292 25630
rect 26236 25394 26292 25564
rect 26236 25342 26238 25394
rect 26290 25342 26292 25394
rect 25788 23940 25844 24220
rect 25844 23884 25956 23940
rect 25788 23874 25844 23884
rect 25340 23762 25396 23772
rect 25676 23492 25732 23502
rect 25676 23266 25732 23436
rect 25676 23214 25678 23266
rect 25730 23214 25732 23266
rect 25676 23202 25732 23214
rect 25788 23380 25844 23390
rect 25788 22932 25844 23324
rect 25788 22838 25844 22876
rect 25564 22820 25620 22830
rect 25564 22482 25620 22764
rect 25564 22430 25566 22482
rect 25618 22430 25620 22482
rect 25340 20916 25396 20926
rect 25340 20822 25396 20860
rect 25564 20802 25620 22430
rect 25676 22370 25732 22382
rect 25676 22318 25678 22370
rect 25730 22318 25732 22370
rect 25676 22036 25732 22318
rect 25900 22260 25956 23884
rect 26124 23828 26180 23838
rect 25900 22194 25956 22204
rect 26012 23604 26068 23614
rect 26012 22930 26068 23548
rect 26012 22878 26014 22930
rect 26066 22878 26068 22930
rect 26012 22036 26068 22878
rect 26124 22596 26180 23772
rect 26236 23716 26292 25342
rect 26236 23650 26292 23660
rect 26348 25394 26404 26236
rect 26348 25342 26350 25394
rect 26402 25342 26404 25394
rect 26124 22530 26180 22540
rect 26236 23154 26292 23166
rect 26236 23102 26238 23154
rect 26290 23102 26292 23154
rect 25676 21970 25732 21980
rect 25788 21980 26068 22036
rect 25788 21812 25844 21980
rect 25564 20750 25566 20802
rect 25618 20750 25620 20802
rect 25564 20738 25620 20750
rect 25676 21756 25844 21812
rect 26012 21812 26068 21822
rect 25676 20244 25732 21756
rect 26012 21718 26068 21756
rect 25788 20692 25844 20702
rect 25788 20690 26180 20692
rect 25788 20638 25790 20690
rect 25842 20638 26180 20690
rect 25788 20636 26180 20638
rect 25788 20626 25844 20636
rect 26012 20468 26068 20478
rect 25900 20356 25956 20366
rect 25340 20188 25732 20244
rect 25788 20244 25844 20254
rect 25340 19346 25396 20188
rect 25564 20020 25620 20030
rect 25340 19294 25342 19346
rect 25394 19294 25396 19346
rect 25340 19282 25396 19294
rect 25452 19796 25508 19806
rect 25340 18004 25396 18014
rect 25340 17666 25396 17948
rect 25452 17890 25508 19740
rect 25452 17838 25454 17890
rect 25506 17838 25508 17890
rect 25452 17826 25508 17838
rect 25340 17614 25342 17666
rect 25394 17614 25396 17666
rect 25340 17602 25396 17614
rect 25564 17108 25620 19964
rect 25788 19346 25844 20188
rect 25788 19294 25790 19346
rect 25842 19294 25844 19346
rect 25788 19282 25844 19294
rect 25900 20018 25956 20300
rect 25900 19966 25902 20018
rect 25954 19966 25956 20018
rect 25900 18788 25956 19966
rect 26012 20244 26068 20412
rect 26012 20018 26068 20188
rect 26012 19966 26014 20018
rect 26066 19966 26068 20018
rect 26012 19954 26068 19966
rect 25900 18722 25956 18732
rect 25676 18340 25732 18350
rect 25676 18246 25732 18284
rect 25564 16976 25620 17052
rect 25676 17890 25732 17902
rect 25676 17838 25678 17890
rect 25730 17838 25732 17890
rect 25676 17442 25732 17838
rect 25676 17390 25678 17442
rect 25730 17390 25732 17442
rect 25228 16828 25620 16884
rect 25116 16716 25284 16772
rect 24836 16492 24948 16548
rect 24780 16482 24836 16492
rect 24780 16100 24836 16110
rect 24780 15876 24836 16044
rect 24780 15538 24836 15820
rect 24892 15764 24948 16492
rect 25004 15876 25060 16492
rect 25116 16100 25172 16110
rect 25116 16006 25172 16044
rect 25004 15820 25172 15876
rect 24892 15708 25060 15764
rect 24780 15486 24782 15538
rect 24834 15486 24836 15538
rect 24780 15148 24836 15486
rect 24892 15316 24948 15326
rect 24892 15222 24948 15260
rect 24780 15092 24948 15148
rect 24668 14366 24670 14418
rect 24722 14366 24724 14418
rect 24668 14354 24724 14366
rect 24332 14308 24388 14346
rect 24332 14242 24388 14252
rect 24220 13918 24222 13970
rect 24274 13918 24276 13970
rect 24220 13906 24276 13918
rect 24332 14084 24388 14094
rect 24108 13694 24110 13746
rect 24162 13694 24164 13746
rect 23996 12852 24052 12862
rect 23772 12850 24052 12852
rect 23772 12798 23998 12850
rect 24050 12798 24052 12850
rect 23772 12796 24052 12798
rect 23660 12404 23716 12414
rect 23548 12402 23716 12404
rect 23548 12350 23662 12402
rect 23714 12350 23716 12402
rect 23548 12348 23716 12350
rect 23212 12180 23268 12190
rect 23212 12178 23380 12180
rect 23212 12126 23214 12178
rect 23266 12126 23380 12178
rect 23212 12124 23380 12126
rect 23212 12114 23268 12124
rect 22988 11340 23156 11396
rect 23212 11396 23268 11406
rect 22764 10994 22820 11004
rect 22876 11282 22932 11294
rect 22876 11230 22878 11282
rect 22930 11230 22932 11282
rect 22484 8876 22708 8932
rect 22764 10052 22820 10062
rect 22316 6804 22372 6814
rect 21756 6748 21924 6804
rect 21756 6578 21812 6590
rect 21756 6526 21758 6578
rect 21810 6526 21812 6578
rect 21756 6020 21812 6526
rect 21756 5954 21812 5964
rect 21644 5796 21700 5806
rect 21644 5702 21700 5740
rect 21532 5182 21534 5234
rect 21586 5182 21588 5234
rect 21532 5170 21588 5182
rect 21868 5236 21924 6748
rect 22092 6692 22148 6702
rect 22092 6578 22148 6636
rect 22092 6526 22094 6578
rect 22146 6526 22148 6578
rect 22092 6514 22148 6526
rect 22316 6130 22372 6748
rect 22316 6078 22318 6130
rect 22370 6078 22372 6130
rect 22316 6066 22372 6078
rect 21868 5170 21924 5180
rect 22092 5460 22148 5470
rect 22092 5234 22148 5404
rect 22092 5182 22094 5234
rect 22146 5182 22148 5234
rect 22092 5170 22148 5182
rect 22428 5124 22484 8876
rect 22764 8484 22820 9996
rect 22540 8036 22596 8046
rect 22540 7942 22596 7980
rect 22764 7700 22820 8428
rect 22652 7644 22820 7700
rect 22540 7362 22596 7374
rect 22540 7310 22542 7362
rect 22594 7310 22596 7362
rect 22540 6692 22596 7310
rect 22540 6626 22596 6636
rect 22540 6468 22596 6478
rect 22652 6468 22708 7644
rect 22876 7588 22932 11230
rect 22988 9156 23044 11340
rect 23100 11170 23156 11182
rect 23100 11118 23102 11170
rect 23154 11118 23156 11170
rect 23100 11060 23156 11118
rect 23100 10994 23156 11004
rect 23212 10948 23268 11340
rect 23212 10882 23268 10892
rect 22988 9090 23044 9100
rect 23100 10610 23156 10622
rect 23100 10558 23102 10610
rect 23154 10558 23156 10610
rect 23100 9940 23156 10558
rect 23324 10052 23380 12124
rect 23548 12068 23604 12348
rect 23660 12338 23716 12348
rect 23324 9986 23380 9996
rect 23436 12012 23604 12068
rect 23100 9492 23156 9884
rect 23212 9604 23268 9614
rect 23436 9604 23492 12012
rect 23660 11732 23716 11742
rect 23212 9602 23492 9604
rect 23212 9550 23214 9602
rect 23266 9550 23492 9602
rect 23212 9548 23492 9550
rect 23548 10388 23604 10398
rect 23212 9538 23268 9548
rect 22988 8930 23044 8942
rect 22988 8878 22990 8930
rect 23042 8878 23044 8930
rect 22988 8596 23044 8878
rect 22988 8530 23044 8540
rect 23100 8372 23156 9436
rect 22764 7474 22820 7486
rect 22764 7422 22766 7474
rect 22818 7422 22820 7474
rect 22764 7364 22820 7422
rect 22764 7298 22820 7308
rect 22876 6804 22932 7532
rect 22876 6738 22932 6748
rect 22988 8316 23156 8372
rect 23212 9156 23268 9166
rect 22988 6690 23044 8316
rect 23100 8148 23156 8158
rect 23100 8054 23156 8092
rect 22988 6638 22990 6690
rect 23042 6638 23044 6690
rect 22988 6626 23044 6638
rect 22540 6466 22708 6468
rect 22540 6414 22542 6466
rect 22594 6414 22708 6466
rect 22540 6412 22708 6414
rect 22764 6580 22820 6590
rect 22540 6402 22596 6412
rect 22764 6130 22820 6524
rect 22764 6078 22766 6130
rect 22818 6078 22820 6130
rect 22764 6066 22820 6078
rect 22316 5122 22484 5124
rect 22316 5070 22430 5122
rect 22482 5070 22484 5122
rect 22316 5068 22484 5070
rect 20300 4898 20804 4900
rect 20300 4846 20302 4898
rect 20354 4846 20804 4898
rect 20300 4844 20804 4846
rect 20300 4834 20356 4844
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20748 4676 20804 4844
rect 20748 4620 21364 4676
rect 19964 4564 20020 4574
rect 20412 4564 20468 4574
rect 19628 4562 20468 4564
rect 19628 4510 19966 4562
rect 20018 4510 20414 4562
rect 20466 4510 20468 4562
rect 19628 4508 20468 4510
rect 19964 4498 20020 4508
rect 20412 4498 20468 4508
rect 21308 4562 21364 4620
rect 21308 4510 21310 4562
rect 21362 4510 21364 4562
rect 21308 4498 21364 4510
rect 22316 4452 22372 5068
rect 22428 5058 22484 5068
rect 22540 6020 22596 6030
rect 22428 4564 22484 4574
rect 22540 4564 22596 5964
rect 22988 5236 23044 5246
rect 22988 5142 23044 5180
rect 22428 4562 22596 4564
rect 22428 4510 22430 4562
rect 22482 4510 22596 4562
rect 22428 4508 22596 4510
rect 22428 4498 22484 4508
rect 22316 4386 22372 4396
rect 20188 4004 20244 4014
rect 18956 3726 18958 3778
rect 19010 3726 19012 3778
rect 18956 3714 19012 3726
rect 19292 3892 19348 3902
rect 19292 3666 19348 3836
rect 19292 3614 19294 3666
rect 19346 3614 19348 3666
rect 19292 3602 19348 3614
rect 19740 3778 19796 3790
rect 19740 3726 19742 3778
rect 19794 3726 19796 3778
rect 19740 3666 19796 3726
rect 19740 3614 19742 3666
rect 19794 3614 19796 3666
rect 19740 3602 19796 3614
rect 20188 3666 20244 3948
rect 23212 3780 23268 9100
rect 23436 8932 23492 8942
rect 23548 8932 23604 10332
rect 23324 8930 23604 8932
rect 23324 8878 23438 8930
rect 23490 8878 23604 8930
rect 23324 8876 23604 8878
rect 23660 8930 23716 11676
rect 23772 11172 23828 11182
rect 23772 10052 23828 11116
rect 23996 10948 24052 12796
rect 24108 11732 24164 13694
rect 24332 13188 24388 14028
rect 24780 13972 24836 13982
rect 24780 13878 24836 13916
rect 24332 13132 24612 13188
rect 24220 12852 24276 12862
rect 24220 12404 24276 12796
rect 24220 12402 24500 12404
rect 24220 12350 24222 12402
rect 24274 12350 24500 12402
rect 24220 12348 24500 12350
rect 24220 12338 24276 12348
rect 24108 11282 24164 11676
rect 24108 11230 24110 11282
rect 24162 11230 24164 11282
rect 24108 11218 24164 11230
rect 24220 12180 24276 12190
rect 23996 10892 24164 10948
rect 24108 10724 24164 10892
rect 24220 10834 24276 12124
rect 24220 10782 24222 10834
rect 24274 10782 24276 10834
rect 24220 10770 24276 10782
rect 23884 10612 23940 10622
rect 23884 10518 23940 10556
rect 23996 10610 24052 10622
rect 23996 10558 23998 10610
rect 24050 10558 24052 10610
rect 23996 10164 24052 10558
rect 24108 10612 24164 10668
rect 24332 10612 24388 10622
rect 24108 10610 24388 10612
rect 24108 10558 24334 10610
rect 24386 10558 24388 10610
rect 24108 10556 24388 10558
rect 24332 10388 24388 10556
rect 24332 10322 24388 10332
rect 23996 10108 24276 10164
rect 24220 10052 24276 10108
rect 23772 9996 24164 10052
rect 23660 8878 23662 8930
rect 23714 8878 23716 8930
rect 23324 7364 23380 8876
rect 23436 8866 23492 8876
rect 23660 8866 23716 8878
rect 23772 9828 23828 9838
rect 23772 9602 23828 9772
rect 24108 9714 24164 9996
rect 24108 9662 24110 9714
rect 24162 9662 24164 9714
rect 24108 9650 24164 9662
rect 23772 9550 23774 9602
rect 23826 9550 23828 9602
rect 23772 8708 23828 9550
rect 23996 9380 24052 9390
rect 23996 9266 24052 9324
rect 23996 9214 23998 9266
rect 24050 9214 24052 9266
rect 23996 9202 24052 9214
rect 24220 9268 24276 9996
rect 24220 9202 24276 9212
rect 23436 8652 23828 8708
rect 23436 8146 23492 8652
rect 23436 8094 23438 8146
rect 23490 8094 23492 8146
rect 23436 8082 23492 8094
rect 23884 8036 23940 8046
rect 23772 8034 23940 8036
rect 23772 7982 23886 8034
rect 23938 7982 23940 8034
rect 23772 7980 23940 7982
rect 23436 7364 23492 7374
rect 23324 7362 23492 7364
rect 23324 7310 23438 7362
rect 23490 7310 23492 7362
rect 23324 7308 23492 7310
rect 23436 7252 23492 7308
rect 23436 7186 23492 7196
rect 23548 7364 23604 7374
rect 23548 6916 23604 7308
rect 23772 7252 23828 7980
rect 23884 7970 23940 7980
rect 23772 7186 23828 7196
rect 23884 7700 23940 7710
rect 23884 7028 23940 7644
rect 24444 7700 24500 12348
rect 24556 12402 24612 13132
rect 24556 12350 24558 12402
rect 24610 12350 24612 12402
rect 24556 12338 24612 12350
rect 24668 13186 24724 13198
rect 24668 13134 24670 13186
rect 24722 13134 24724 13186
rect 24668 12738 24724 13134
rect 24892 13186 24948 15092
rect 25004 14420 25060 15708
rect 25116 14980 25172 15820
rect 25228 15148 25284 16716
rect 25452 16436 25508 16446
rect 25452 15986 25508 16380
rect 25452 15934 25454 15986
rect 25506 15934 25508 15986
rect 25452 15428 25508 15934
rect 25452 15362 25508 15372
rect 25228 15092 25508 15148
rect 25116 14924 25284 14980
rect 25228 14642 25284 14924
rect 25452 14868 25508 15092
rect 25564 15090 25620 16828
rect 25564 15038 25566 15090
rect 25618 15038 25620 15090
rect 25564 15026 25620 15038
rect 25452 14812 25620 14868
rect 25228 14590 25230 14642
rect 25282 14590 25284 14642
rect 25228 14578 25284 14590
rect 25564 14420 25620 14812
rect 25004 14364 25508 14420
rect 24892 13134 24894 13186
rect 24946 13134 24948 13186
rect 24892 13122 24948 13134
rect 25228 13300 25284 13310
rect 24668 12686 24670 12738
rect 24722 12686 24724 12738
rect 24668 11844 24724 12686
rect 24668 11788 24836 11844
rect 24668 11396 24724 11406
rect 24668 11282 24724 11340
rect 24668 11230 24670 11282
rect 24722 11230 24724 11282
rect 24668 10276 24724 11230
rect 24780 10500 24836 11788
rect 24780 10406 24836 10444
rect 24892 11394 24948 11406
rect 24892 11342 24894 11394
rect 24946 11342 24948 11394
rect 24556 9602 24612 9614
rect 24556 9550 24558 9602
rect 24610 9550 24612 9602
rect 24556 9156 24612 9550
rect 24556 9090 24612 9100
rect 24556 8930 24612 8942
rect 24556 8878 24558 8930
rect 24610 8878 24612 8930
rect 24556 8818 24612 8878
rect 24556 8766 24558 8818
rect 24610 8766 24612 8818
rect 24556 8754 24612 8766
rect 24668 8370 24724 10220
rect 24668 8318 24670 8370
rect 24722 8318 24724 8370
rect 24668 8306 24724 8318
rect 24892 9044 24948 11342
rect 25228 11284 25284 13244
rect 25340 12964 25396 12974
rect 25340 12870 25396 12908
rect 25452 12404 25508 14364
rect 25564 14326 25620 14364
rect 25564 13634 25620 13646
rect 25564 13582 25566 13634
rect 25618 13582 25620 13634
rect 25564 12850 25620 13582
rect 25564 12798 25566 12850
rect 25618 12798 25620 12850
rect 25564 12786 25620 12798
rect 25564 12404 25620 12414
rect 25452 12402 25620 12404
rect 25452 12350 25566 12402
rect 25618 12350 25620 12402
rect 25452 12348 25620 12350
rect 25564 12338 25620 12348
rect 25452 11956 25508 11966
rect 25228 11218 25284 11228
rect 25340 11954 25508 11956
rect 25340 11902 25454 11954
rect 25506 11902 25508 11954
rect 25340 11900 25508 11902
rect 24444 7634 24500 7644
rect 24892 7698 24948 8988
rect 24892 7646 24894 7698
rect 24946 7646 24948 7698
rect 24892 7634 24948 7646
rect 25228 8034 25284 8046
rect 25228 7982 25230 8034
rect 25282 7982 25284 8034
rect 23884 6962 23940 6972
rect 24556 7474 24612 7486
rect 24556 7422 24558 7474
rect 24610 7422 24612 7474
rect 23548 6690 23604 6860
rect 24332 6804 24388 6814
rect 24332 6710 24388 6748
rect 23548 6638 23550 6690
rect 23602 6638 23604 6690
rect 23436 6580 23492 6590
rect 23436 6130 23492 6524
rect 23436 6078 23438 6130
rect 23490 6078 23492 6130
rect 23436 5012 23492 6078
rect 23548 5236 23604 6638
rect 23772 6692 23828 6702
rect 23772 6598 23828 6636
rect 23884 6580 23940 6590
rect 23884 6486 23940 6524
rect 24556 6580 24612 7422
rect 24332 6020 24388 6030
rect 24556 6020 24612 6524
rect 24892 7476 24948 7486
rect 24892 6578 24948 7420
rect 25228 6916 25284 7982
rect 25340 8036 25396 11900
rect 25452 11890 25508 11900
rect 25564 11282 25620 11294
rect 25564 11230 25566 11282
rect 25618 11230 25620 11282
rect 25564 11172 25620 11230
rect 25564 10836 25620 11116
rect 25564 10770 25620 10780
rect 25676 10612 25732 17390
rect 25788 17556 25844 17566
rect 25788 15538 25844 17500
rect 26124 16210 26180 20636
rect 26236 20242 26292 23102
rect 26348 23044 26404 25342
rect 26460 25284 26516 26852
rect 26460 25218 26516 25228
rect 26572 26068 26628 26078
rect 26348 22370 26404 22988
rect 26460 24836 26516 24846
rect 26460 22708 26516 24780
rect 26572 22820 26628 26012
rect 26572 22754 26628 22764
rect 26460 22642 26516 22652
rect 26684 22596 26740 28364
rect 27020 28308 27076 31388
rect 27356 31218 27412 32510
rect 27356 31166 27358 31218
rect 27410 31166 27412 31218
rect 27356 31154 27412 31166
rect 27356 29426 27412 29438
rect 27356 29374 27358 29426
rect 27410 29374 27412 29426
rect 27356 28868 27412 29374
rect 27356 28802 27412 28812
rect 27356 28532 27412 28542
rect 27356 28438 27412 28476
rect 27132 28420 27188 28430
rect 27132 28326 27188 28364
rect 27244 28418 27300 28430
rect 27244 28366 27246 28418
rect 27298 28366 27300 28418
rect 26908 28252 27076 28308
rect 26796 27746 26852 27758
rect 26796 27694 26798 27746
rect 26850 27694 26852 27746
rect 26796 27636 26852 27694
rect 26796 27570 26852 27580
rect 26796 25284 26852 25294
rect 26796 25190 26852 25228
rect 26908 24948 26964 28252
rect 27244 27972 27300 28366
rect 27244 27906 27300 27916
rect 27132 27858 27188 27870
rect 27132 27806 27134 27858
rect 27186 27806 27188 27858
rect 27020 27076 27076 27086
rect 27132 27076 27188 27806
rect 27020 27074 27188 27076
rect 27020 27022 27022 27074
rect 27074 27022 27188 27074
rect 27020 27020 27188 27022
rect 27020 27010 27076 27020
rect 27132 26964 27188 27020
rect 27132 26898 27188 26908
rect 27244 27300 27300 27310
rect 27132 26516 27188 26526
rect 27132 26422 27188 26460
rect 27244 25060 27300 27244
rect 27468 26292 27524 35644
rect 27804 34916 27860 34926
rect 27804 34822 27860 34860
rect 27916 34130 27972 34142
rect 27916 34078 27918 34130
rect 27970 34078 27972 34130
rect 27916 33570 27972 34078
rect 27916 33518 27918 33570
rect 27970 33518 27972 33570
rect 27916 33506 27972 33518
rect 27580 33348 27636 33358
rect 27580 33254 27636 33292
rect 28028 33348 28084 33358
rect 27692 32450 27748 32462
rect 27692 32398 27694 32450
rect 27746 32398 27748 32450
rect 27692 32004 27748 32398
rect 27692 31938 27748 31948
rect 28028 32452 28084 33292
rect 28140 32676 28196 38892
rect 28252 38724 28308 38762
rect 28252 32788 28308 38668
rect 28364 38052 28420 38062
rect 28364 37958 28420 37996
rect 28364 35812 28420 35822
rect 28364 35026 28420 35756
rect 28364 34974 28366 35026
rect 28418 34974 28420 35026
rect 28364 34962 28420 34974
rect 28476 33348 28532 42924
rect 28700 42420 28756 45612
rect 28924 45332 28980 45838
rect 28924 45266 28980 45276
rect 29036 43426 29092 43438
rect 29036 43374 29038 43426
rect 29090 43374 29092 43426
rect 28812 42644 28868 42654
rect 28812 42550 28868 42588
rect 28700 42364 28868 42420
rect 28588 42084 28644 42094
rect 28588 41186 28644 42028
rect 28588 41134 28590 41186
rect 28642 41134 28644 41186
rect 28588 41122 28644 41134
rect 28700 41076 28756 41086
rect 28700 40982 28756 41020
rect 28812 40852 28868 42364
rect 28700 40796 28868 40852
rect 28924 40962 28980 40974
rect 28924 40910 28926 40962
rect 28978 40910 28980 40962
rect 28700 38668 28756 40796
rect 28812 40404 28868 40414
rect 28812 38946 28868 40348
rect 28924 40402 28980 40910
rect 28924 40350 28926 40402
rect 28978 40350 28980 40402
rect 28924 40338 28980 40350
rect 29036 40292 29092 43374
rect 29036 40226 29092 40236
rect 29148 40404 29204 40414
rect 29148 40290 29204 40348
rect 29148 40238 29150 40290
rect 29202 40238 29204 40290
rect 29148 40226 29204 40238
rect 28812 38894 28814 38946
rect 28866 38894 28868 38946
rect 28812 38882 28868 38894
rect 28700 38612 28980 38668
rect 28812 38052 28868 38062
rect 28812 37378 28868 37996
rect 28812 37326 28814 37378
rect 28866 37326 28868 37378
rect 28812 37314 28868 37326
rect 28476 33216 28532 33292
rect 28812 33460 28868 33470
rect 28812 33234 28868 33404
rect 28812 33182 28814 33234
rect 28866 33182 28868 33234
rect 28812 33170 28868 33182
rect 28252 32732 28532 32788
rect 28140 32620 28420 32676
rect 28140 32452 28196 32462
rect 28028 32450 28308 32452
rect 28028 32398 28142 32450
rect 28194 32398 28308 32450
rect 28028 32396 28308 32398
rect 28028 31668 28084 32396
rect 28140 32386 28196 32396
rect 27580 31612 28084 31668
rect 27580 31218 27636 31612
rect 28140 31556 28196 31566
rect 27580 31166 27582 31218
rect 27634 31166 27636 31218
rect 27580 31154 27636 31166
rect 27692 31554 28196 31556
rect 27692 31502 28142 31554
rect 28194 31502 28196 31554
rect 27692 31500 28196 31502
rect 27692 31106 27748 31500
rect 28140 31490 28196 31500
rect 28252 31218 28308 32396
rect 28252 31166 28254 31218
rect 28306 31166 28308 31218
rect 28252 31154 28308 31166
rect 27692 31054 27694 31106
rect 27746 31054 27748 31106
rect 27692 31042 27748 31054
rect 28140 30212 28196 30222
rect 28140 30118 28196 30156
rect 27580 29540 27636 29550
rect 27580 29446 27636 29484
rect 27916 29540 27972 29550
rect 27916 28756 27972 29484
rect 27916 28642 27972 28700
rect 27916 28590 27918 28642
rect 27970 28590 27972 28642
rect 27916 28578 27972 28590
rect 28028 29314 28084 29326
rect 28028 29262 28030 29314
rect 28082 29262 28084 29314
rect 28028 28644 28084 29262
rect 28028 28196 28084 28588
rect 28252 28418 28308 28430
rect 28252 28366 28254 28418
rect 28306 28366 28308 28418
rect 28252 28196 28308 28366
rect 27916 28140 28308 28196
rect 27916 27412 27972 28140
rect 28140 27972 28196 27982
rect 27916 27346 27972 27356
rect 28028 27970 28196 27972
rect 28028 27918 28142 27970
rect 28194 27918 28196 27970
rect 28028 27916 28196 27918
rect 27692 27188 27748 27198
rect 28028 27188 28084 27916
rect 28140 27906 28196 27916
rect 28252 27972 28308 27982
rect 28252 27878 28308 27916
rect 28140 27636 28196 27646
rect 28364 27636 28420 32620
rect 28476 30212 28532 32732
rect 28700 30212 28756 30222
rect 28476 30156 28644 30212
rect 28476 29988 28532 29998
rect 28476 29894 28532 29932
rect 28588 29764 28644 30156
rect 28700 30098 28756 30156
rect 28700 30046 28702 30098
rect 28754 30046 28756 30098
rect 28700 30034 28756 30046
rect 28812 30098 28868 30110
rect 28812 30046 28814 30098
rect 28866 30046 28868 30098
rect 28140 27634 28420 27636
rect 28140 27582 28142 27634
rect 28194 27582 28420 27634
rect 28140 27580 28420 27582
rect 28476 29708 28644 29764
rect 28812 29764 28868 30046
rect 28140 27570 28196 27580
rect 28476 27524 28532 29708
rect 28812 29698 28868 29708
rect 28364 27468 28532 27524
rect 28588 28868 28644 28878
rect 28252 27412 28308 27422
rect 27692 27186 28084 27188
rect 27692 27134 27694 27186
rect 27746 27134 28084 27186
rect 27692 27132 28084 27134
rect 27692 27122 27748 27132
rect 27468 26226 27524 26236
rect 27580 26964 27636 26974
rect 27468 26068 27524 26078
rect 27356 26066 27524 26068
rect 27356 26014 27470 26066
rect 27522 26014 27524 26066
rect 27356 26012 27524 26014
rect 27356 25284 27412 26012
rect 27468 26002 27524 26012
rect 27580 25396 27636 26908
rect 27804 26740 27860 26750
rect 27692 26178 27748 26190
rect 27692 26126 27694 26178
rect 27746 26126 27748 26178
rect 27692 25956 27748 26126
rect 27692 25890 27748 25900
rect 27692 25732 27748 25742
rect 27804 25732 27860 26684
rect 28028 26292 28084 27132
rect 28140 27188 28196 27198
rect 28140 27094 28196 27132
rect 28252 26852 28308 27356
rect 28252 26786 28308 26796
rect 28364 26740 28420 27468
rect 28588 27412 28644 28812
rect 28700 28756 28756 28766
rect 28700 28662 28756 28700
rect 28700 27746 28756 27758
rect 28700 27694 28702 27746
rect 28754 27694 28756 27746
rect 28700 27636 28756 27694
rect 28700 27570 28756 27580
rect 28364 26674 28420 26684
rect 28476 27356 28644 27412
rect 28252 26516 28308 26526
rect 28476 26516 28532 27356
rect 28700 27188 28756 27198
rect 28588 27076 28644 27086
rect 28588 26982 28644 27020
rect 28252 26514 28532 26516
rect 28252 26462 28254 26514
rect 28306 26462 28532 26514
rect 28252 26460 28532 26462
rect 28700 26516 28756 27132
rect 28924 26908 28980 38612
rect 29036 38610 29092 38622
rect 29036 38558 29038 38610
rect 29090 38558 29092 38610
rect 29036 38052 29092 38558
rect 29036 37986 29092 37996
rect 29260 28308 29316 50372
rect 29484 48356 29540 50652
rect 30044 49924 30100 49934
rect 30044 49830 30100 49868
rect 30268 49810 30324 49822
rect 30268 49758 30270 49810
rect 30322 49758 30324 49810
rect 30268 49140 30324 49758
rect 30268 49026 30324 49084
rect 30268 48974 30270 49026
rect 30322 48974 30324 49026
rect 30268 48962 30324 48974
rect 30604 49028 30660 49038
rect 30604 48934 30660 48972
rect 29596 48916 29652 48926
rect 29596 48822 29652 48860
rect 30044 48916 30100 48926
rect 30044 48822 30100 48860
rect 30492 48916 30548 48926
rect 29484 48290 29540 48300
rect 30268 48802 30324 48814
rect 30268 48750 30270 48802
rect 30322 48750 30324 48802
rect 29708 48244 29764 48254
rect 29708 48150 29764 48188
rect 29932 48132 29988 48142
rect 29932 48038 29988 48076
rect 29372 48018 29428 48030
rect 29372 47966 29374 48018
rect 29426 47966 29428 48018
rect 29372 46228 29428 47966
rect 30044 47460 30100 47470
rect 29932 47458 30100 47460
rect 29932 47406 30046 47458
rect 30098 47406 30100 47458
rect 29932 47404 30100 47406
rect 29372 46162 29428 46172
rect 29708 46676 29764 46686
rect 29708 45218 29764 46620
rect 29932 46450 29988 47404
rect 30044 47394 30100 47404
rect 30156 47236 30212 47246
rect 30156 47142 30212 47180
rect 30268 46676 30324 48750
rect 29932 46398 29934 46450
rect 29986 46398 29988 46450
rect 29820 46228 29876 46238
rect 29820 46002 29876 46172
rect 29820 45950 29822 46002
rect 29874 45950 29876 46002
rect 29820 45938 29876 45950
rect 29932 45892 29988 46398
rect 29932 45760 29988 45836
rect 30044 46562 30100 46574
rect 30044 46510 30046 46562
rect 30098 46510 30100 46562
rect 30268 46544 30324 46620
rect 30492 48242 30548 48860
rect 30492 48190 30494 48242
rect 30546 48190 30548 48242
rect 29708 45166 29710 45218
rect 29762 45166 29764 45218
rect 29708 45154 29764 45166
rect 29932 45108 29988 45118
rect 30044 45108 30100 46510
rect 30268 45332 30324 45342
rect 30268 45238 30324 45276
rect 29988 45052 30100 45108
rect 29932 45014 29988 45052
rect 29932 44324 29988 44334
rect 29820 44322 29988 44324
rect 29820 44270 29934 44322
rect 29986 44270 29988 44322
rect 29820 44268 29988 44270
rect 29596 44210 29652 44222
rect 29596 44158 29598 44210
rect 29650 44158 29652 44210
rect 29596 43538 29652 44158
rect 29596 43486 29598 43538
rect 29650 43486 29652 43538
rect 29596 42756 29652 43486
rect 29820 43540 29876 44268
rect 29932 44258 29988 44268
rect 30380 44322 30436 44334
rect 30380 44270 30382 44322
rect 30434 44270 30436 44322
rect 30380 44212 30436 44270
rect 30380 44146 30436 44156
rect 29820 42978 29876 43484
rect 29820 42926 29822 42978
rect 29874 42926 29876 42978
rect 29820 42914 29876 42926
rect 29596 42690 29652 42700
rect 30380 42756 30436 42766
rect 29372 42644 29428 42654
rect 29372 29876 29428 42588
rect 30268 42644 30324 42654
rect 30268 42550 30324 42588
rect 29596 42084 29652 42094
rect 29596 41186 29652 42028
rect 30380 42084 30436 42700
rect 30492 42532 30548 48190
rect 30828 48354 30884 48366
rect 30828 48302 30830 48354
rect 30882 48302 30884 48354
rect 30828 48020 30884 48302
rect 30828 47954 30884 47964
rect 30940 48132 30996 48142
rect 30940 47348 30996 48076
rect 30940 47254 30996 47292
rect 30604 45778 30660 45790
rect 30604 45726 30606 45778
rect 30658 45726 30660 45778
rect 30604 44324 30660 45726
rect 30716 45332 30772 45342
rect 30716 45108 30772 45276
rect 31052 45220 31108 55468
rect 31388 55412 31668 55468
rect 33628 56308 33684 56318
rect 31388 55410 31444 55412
rect 31388 55358 31390 55410
rect 31442 55358 31444 55410
rect 31388 55346 31444 55358
rect 31612 55356 32004 55412
rect 31948 55186 32004 55356
rect 31948 55134 31950 55186
rect 32002 55134 32004 55186
rect 31948 55122 32004 55134
rect 33628 55188 33684 56252
rect 37212 56082 37268 56094
rect 37212 56030 37214 56082
rect 37266 56030 37268 56082
rect 36428 55970 36484 55982
rect 36428 55918 36430 55970
rect 36482 55918 36484 55970
rect 36428 55860 36484 55918
rect 36428 55794 36484 55804
rect 36876 55972 36932 55982
rect 35196 55692 35460 55702
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35196 55626 35460 55636
rect 36876 55300 36932 55916
rect 37212 55860 37268 56030
rect 37884 55970 37940 56590
rect 37884 55918 37886 55970
rect 37938 55918 37940 55970
rect 37884 55906 37940 55918
rect 40012 56084 40068 56094
rect 37212 55794 37268 55804
rect 37772 55300 37828 55310
rect 39788 55300 39844 55310
rect 40012 55300 40068 56028
rect 40908 56082 40964 56094
rect 40908 56030 40910 56082
rect 40962 56030 40964 56082
rect 40908 55468 40964 56030
rect 41244 56084 41300 56094
rect 41244 55990 41300 56028
rect 41580 56082 41636 56094
rect 41580 56030 41582 56082
rect 41634 56030 41636 56082
rect 40572 55412 40964 55468
rect 41132 55970 41188 55982
rect 41132 55918 41134 55970
rect 41186 55918 41188 55970
rect 36876 55234 36932 55244
rect 37660 55298 37828 55300
rect 37660 55246 37774 55298
rect 37826 55246 37828 55298
rect 37660 55244 37828 55246
rect 33628 55122 33684 55132
rect 37548 55188 37604 55198
rect 37548 55094 37604 55132
rect 34412 55074 34468 55086
rect 34412 55022 34414 55074
rect 34466 55022 34468 55074
rect 33628 52946 33684 52958
rect 33628 52894 33630 52946
rect 33682 52894 33684 52946
rect 32284 52836 32340 52846
rect 31948 51940 32004 51950
rect 31612 51380 31668 51390
rect 31164 50372 31220 50382
rect 31164 49810 31220 50316
rect 31612 49922 31668 51324
rect 31948 50428 32004 51884
rect 32284 51266 32340 52780
rect 32732 52388 32788 52398
rect 32508 52162 32564 52174
rect 32508 52110 32510 52162
rect 32562 52110 32564 52162
rect 32284 51214 32286 51266
rect 32338 51214 32340 51266
rect 32396 51380 32452 51390
rect 32508 51380 32564 52110
rect 32732 52050 32788 52332
rect 33180 52164 33236 52174
rect 33180 52070 33236 52108
rect 32732 51998 32734 52050
rect 32786 51998 32788 52050
rect 32732 51986 32788 51998
rect 33628 52052 33684 52894
rect 33964 52946 34020 52958
rect 33964 52894 33966 52946
rect 34018 52894 34020 52946
rect 33740 52836 33796 52846
rect 33740 52742 33796 52780
rect 33852 52276 33908 52286
rect 33852 52162 33908 52220
rect 33852 52110 33854 52162
rect 33906 52110 33908 52162
rect 33852 52098 33908 52110
rect 33964 52164 34020 52894
rect 34188 52946 34244 52958
rect 34188 52894 34190 52946
rect 34242 52894 34244 52946
rect 34188 52388 34244 52894
rect 33964 52098 34020 52108
rect 34076 52332 34244 52388
rect 34300 52724 34356 52734
rect 32452 51324 32564 51380
rect 32620 51938 32676 51950
rect 32620 51886 32622 51938
rect 32674 51886 32676 51938
rect 32396 51248 32452 51324
rect 32284 51202 32340 51214
rect 31836 50372 31892 50382
rect 31948 50372 32340 50428
rect 31836 50278 31892 50316
rect 31612 49870 31614 49922
rect 31666 49870 31668 49922
rect 31612 49858 31668 49870
rect 31164 49758 31166 49810
rect 31218 49758 31220 49810
rect 31164 48916 31220 49758
rect 32060 49700 32116 49710
rect 32172 49700 32228 49710
rect 32060 49698 32172 49700
rect 32060 49646 32062 49698
rect 32114 49646 32172 49698
rect 32060 49644 32172 49646
rect 32060 49634 32116 49644
rect 31276 49140 31332 49150
rect 31276 49046 31332 49084
rect 31500 49140 31556 49150
rect 31276 48916 31332 48926
rect 31164 48860 31276 48916
rect 31164 48244 31220 48254
rect 31276 48244 31332 48860
rect 31388 48804 31444 48814
rect 31388 48710 31444 48748
rect 31388 48468 31444 48478
rect 31500 48468 31556 49084
rect 31612 48916 31668 48926
rect 31612 48822 31668 48860
rect 32172 48914 32228 49644
rect 32172 48862 32174 48914
rect 32226 48862 32228 48914
rect 31388 48466 31556 48468
rect 31388 48414 31390 48466
rect 31442 48414 31556 48466
rect 31388 48412 31556 48414
rect 32172 48804 32228 48862
rect 31388 48402 31444 48412
rect 31724 48244 31780 48254
rect 31276 48242 31780 48244
rect 31276 48190 31726 48242
rect 31778 48190 31780 48242
rect 31276 48188 31780 48190
rect 31164 47458 31220 48188
rect 31724 48178 31780 48188
rect 32172 48132 32228 48748
rect 32172 48066 32228 48076
rect 31164 47406 31166 47458
rect 31218 47406 31220 47458
rect 31164 47394 31220 47406
rect 32060 47684 32116 47694
rect 31836 46450 31892 46462
rect 31836 46398 31838 46450
rect 31890 46398 31892 46450
rect 31836 46116 31892 46398
rect 31836 46050 31892 46060
rect 30940 45164 31108 45220
rect 30828 45108 30884 45118
rect 30716 45106 30884 45108
rect 30716 45054 30830 45106
rect 30882 45054 30884 45106
rect 30716 45052 30884 45054
rect 30828 45042 30884 45052
rect 30940 44772 30996 45164
rect 31724 45108 31780 45118
rect 31052 45052 31332 45108
rect 31052 44994 31108 45052
rect 31052 44942 31054 44994
rect 31106 44942 31108 44994
rect 31052 44930 31108 44942
rect 31276 44996 31332 45052
rect 31724 45014 31780 45052
rect 31276 44940 31444 44996
rect 31164 44882 31220 44894
rect 31164 44830 31166 44882
rect 31218 44830 31220 44882
rect 30940 44716 31108 44772
rect 30604 44268 30884 44324
rect 30604 44100 30660 44110
rect 30604 42754 30660 44044
rect 30604 42702 30606 42754
rect 30658 42702 30660 42754
rect 30604 42690 30660 42702
rect 30492 42476 30660 42532
rect 30380 42018 30436 42028
rect 29596 41134 29598 41186
rect 29650 41134 29652 41186
rect 29596 41122 29652 41134
rect 29932 41076 29988 41086
rect 29932 40982 29988 41020
rect 30156 41074 30212 41086
rect 30156 41022 30158 41074
rect 30210 41022 30212 41074
rect 29820 40962 29876 40974
rect 29820 40910 29822 40962
rect 29874 40910 29876 40962
rect 29708 40516 29764 40526
rect 29596 40292 29652 40302
rect 29596 39842 29652 40236
rect 29596 39790 29598 39842
rect 29650 39790 29652 39842
rect 29484 39284 29540 39294
rect 29484 38668 29540 39228
rect 29596 38836 29652 39790
rect 29708 39732 29764 40460
rect 29820 39844 29876 40910
rect 30044 40402 30100 40414
rect 30044 40350 30046 40402
rect 30098 40350 30100 40402
rect 29820 39788 29988 39844
rect 29708 39676 29876 39732
rect 29820 39506 29876 39676
rect 29820 39454 29822 39506
rect 29874 39454 29876 39506
rect 29820 39442 29876 39454
rect 29708 39396 29764 39406
rect 29708 39302 29764 39340
rect 29820 38836 29876 38846
rect 29596 38834 29876 38836
rect 29596 38782 29822 38834
rect 29874 38782 29876 38834
rect 29596 38780 29876 38782
rect 29820 38770 29876 38780
rect 29484 38612 29652 38668
rect 29484 37156 29540 37166
rect 29484 37062 29540 37100
rect 29484 34018 29540 34030
rect 29484 33966 29486 34018
rect 29538 33966 29540 34018
rect 29484 33572 29540 33966
rect 29484 33506 29540 33516
rect 29596 30436 29652 38612
rect 29708 37828 29764 37838
rect 29708 37734 29764 37772
rect 29932 37826 29988 39788
rect 30044 39284 30100 40350
rect 30156 40404 30212 41022
rect 30156 40338 30212 40348
rect 30492 40404 30548 40414
rect 30492 40310 30548 40348
rect 30604 40180 30660 42476
rect 30044 39218 30100 39228
rect 30492 40124 30660 40180
rect 30268 39172 30324 39182
rect 30268 38946 30324 39116
rect 30268 38894 30270 38946
rect 30322 38894 30324 38946
rect 30268 38882 30324 38894
rect 30044 38836 30100 38846
rect 30044 38162 30100 38780
rect 30380 38836 30436 38846
rect 30380 38742 30436 38780
rect 30492 38668 30548 40124
rect 30604 39394 30660 39406
rect 30604 39342 30606 39394
rect 30658 39342 30660 39394
rect 30604 39284 30660 39342
rect 30604 39218 30660 39228
rect 30044 38110 30046 38162
rect 30098 38110 30100 38162
rect 30044 38098 30100 38110
rect 30380 38612 30548 38668
rect 30828 38668 30884 44268
rect 30940 44210 30996 44222
rect 30940 44158 30942 44210
rect 30994 44158 30996 44210
rect 30940 42644 30996 44158
rect 31052 43316 31108 44716
rect 31164 44212 31220 44830
rect 31164 44098 31220 44156
rect 31164 44046 31166 44098
rect 31218 44046 31220 44098
rect 31164 44034 31220 44046
rect 31276 44210 31332 44222
rect 31276 44158 31278 44210
rect 31330 44158 31332 44210
rect 31276 43764 31332 44158
rect 31052 43250 31108 43260
rect 31164 43708 31332 43764
rect 31052 42980 31108 42990
rect 31164 42980 31220 43708
rect 31276 43540 31332 43550
rect 31388 43540 31444 44940
rect 31500 44210 31556 44222
rect 31500 44158 31502 44210
rect 31554 44158 31556 44210
rect 31500 44100 31556 44158
rect 31500 44034 31556 44044
rect 31724 43540 31780 43550
rect 31388 43538 31780 43540
rect 31388 43486 31726 43538
rect 31778 43486 31780 43538
rect 31388 43484 31780 43486
rect 31276 43446 31332 43484
rect 31724 43474 31780 43484
rect 31948 43428 32004 43438
rect 31052 42978 31220 42980
rect 31052 42926 31054 42978
rect 31106 42926 31220 42978
rect 31052 42924 31220 42926
rect 31276 43204 31332 43214
rect 31052 42756 31108 42924
rect 31052 42690 31108 42700
rect 30940 42578 30996 42588
rect 31164 40290 31220 40302
rect 31164 40238 31166 40290
rect 31218 40238 31220 40290
rect 31164 39618 31220 40238
rect 31164 39566 31166 39618
rect 31218 39566 31220 39618
rect 31164 39284 31220 39566
rect 31164 39218 31220 39228
rect 31276 38668 31332 43148
rect 31948 42866 32004 43372
rect 31948 42814 31950 42866
rect 32002 42814 32004 42866
rect 31948 42802 32004 42814
rect 31500 42756 31556 42766
rect 31388 42754 31556 42756
rect 31388 42702 31502 42754
rect 31554 42702 31556 42754
rect 31388 42700 31556 42702
rect 31388 42532 31444 42700
rect 31500 42690 31556 42700
rect 31724 42756 31780 42766
rect 31724 42662 31780 42700
rect 31388 40852 31444 42476
rect 31612 42196 31668 42206
rect 31612 41858 31668 42140
rect 31836 42084 31892 42094
rect 31836 41972 31892 42028
rect 31612 41806 31614 41858
rect 31666 41806 31668 41858
rect 31500 41076 31556 41086
rect 31500 40982 31556 41020
rect 31612 40852 31668 41806
rect 31724 41970 31892 41972
rect 31724 41918 31838 41970
rect 31890 41918 31892 41970
rect 31724 41916 31892 41918
rect 31724 41074 31780 41916
rect 31836 41906 31892 41916
rect 31724 41022 31726 41074
rect 31778 41022 31780 41074
rect 31724 41010 31780 41022
rect 31836 41074 31892 41086
rect 31836 41022 31838 41074
rect 31890 41022 31892 41074
rect 31836 40852 31892 41022
rect 31388 40796 31556 40852
rect 31612 40796 31892 40852
rect 31388 40402 31444 40414
rect 31388 40350 31390 40402
rect 31442 40350 31444 40402
rect 31388 39508 31444 40350
rect 31388 39442 31444 39452
rect 31500 38668 31556 40796
rect 31724 39730 31780 39742
rect 31724 39678 31726 39730
rect 31778 39678 31780 39730
rect 31612 39508 31668 39518
rect 31612 39414 31668 39452
rect 30828 38612 30996 38668
rect 31276 38612 31444 38668
rect 31500 38612 31668 38668
rect 30156 38052 30212 38062
rect 30156 37958 30212 37996
rect 29932 37774 29934 37826
rect 29986 37774 29988 37826
rect 29932 37492 29988 37774
rect 29932 37426 29988 37436
rect 29708 37268 29764 37278
rect 29708 37174 29764 37212
rect 30044 35700 30100 35710
rect 29820 35698 30100 35700
rect 29820 35646 30046 35698
rect 30098 35646 30100 35698
rect 29820 35644 30100 35646
rect 29708 35476 29764 35486
rect 29708 33684 29764 35420
rect 29820 34354 29876 35644
rect 30044 35634 30100 35644
rect 30044 35364 30100 35374
rect 30044 34802 30100 35308
rect 30044 34750 30046 34802
rect 30098 34750 30100 34802
rect 30044 34738 30100 34750
rect 29820 34302 29822 34354
rect 29874 34302 29876 34354
rect 29820 34290 29876 34302
rect 30044 34244 30100 34254
rect 29932 34242 30100 34244
rect 29932 34190 30046 34242
rect 30098 34190 30100 34242
rect 29932 34188 30100 34190
rect 29708 33628 29876 33684
rect 29708 33460 29764 33470
rect 29708 33366 29764 33404
rect 29708 30436 29764 30446
rect 29596 30434 29764 30436
rect 29596 30382 29710 30434
rect 29762 30382 29764 30434
rect 29596 30380 29764 30382
rect 29708 30370 29764 30380
rect 29596 30100 29652 30110
rect 29596 30006 29652 30044
rect 29708 29986 29764 29998
rect 29708 29934 29710 29986
rect 29762 29934 29764 29986
rect 29372 29820 29652 29876
rect 29484 29652 29540 29662
rect 29484 29558 29540 29596
rect 29372 29538 29428 29550
rect 29372 29486 29374 29538
rect 29426 29486 29428 29538
rect 29372 28532 29428 29486
rect 29596 29428 29652 29820
rect 29372 28466 29428 28476
rect 29484 29372 29652 29428
rect 29260 28242 29316 28252
rect 29484 26908 29540 29372
rect 29596 29202 29652 29214
rect 29596 29150 29598 29202
rect 29650 29150 29652 29202
rect 29596 28420 29652 29150
rect 29708 28868 29764 29934
rect 29708 28802 29764 28812
rect 29596 28354 29652 28364
rect 28252 26450 28308 26460
rect 28700 26450 28756 26460
rect 28812 26852 28980 26908
rect 29260 26852 29540 26908
rect 28476 26292 28532 26302
rect 28028 26236 28420 26292
rect 27692 25730 27860 25732
rect 27692 25678 27694 25730
rect 27746 25678 27860 25730
rect 27692 25676 27860 25678
rect 28252 25956 28308 25966
rect 27692 25666 27748 25676
rect 27692 25396 27748 25406
rect 27580 25394 27748 25396
rect 27580 25342 27694 25394
rect 27746 25342 27748 25394
rect 27580 25340 27748 25342
rect 27356 25218 27412 25228
rect 27244 25004 27524 25060
rect 27020 24948 27076 24958
rect 26908 24946 27076 24948
rect 26908 24894 27022 24946
rect 27074 24894 27076 24946
rect 26908 24892 27076 24894
rect 27020 24882 27076 24892
rect 27244 24836 27300 24846
rect 27244 24742 27300 24780
rect 26908 24722 26964 24734
rect 26908 24670 26910 24722
rect 26962 24670 26964 24722
rect 26796 24052 26852 24062
rect 26796 23716 26852 23996
rect 26908 23828 26964 24670
rect 27356 24722 27412 24734
rect 27356 24670 27358 24722
rect 27410 24670 27412 24722
rect 26908 23762 26964 23772
rect 27020 24388 27076 24398
rect 26796 23650 26852 23660
rect 27020 23154 27076 24332
rect 27244 23828 27300 23838
rect 27244 23734 27300 23772
rect 27020 23102 27022 23154
rect 27074 23102 27076 23154
rect 27020 23090 27076 23102
rect 26796 22596 26852 22606
rect 26684 22594 26852 22596
rect 26684 22542 26798 22594
rect 26850 22542 26852 22594
rect 26684 22540 26852 22542
rect 26796 22530 26852 22540
rect 27244 22596 27300 22606
rect 26348 22318 26350 22370
rect 26402 22318 26404 22370
rect 26348 22306 26404 22318
rect 26460 21812 26516 21822
rect 26460 20916 26516 21756
rect 26684 21700 26740 21710
rect 26684 21606 26740 21644
rect 26572 21588 26628 21598
rect 26572 21494 26628 21532
rect 27020 21586 27076 21598
rect 27020 21534 27022 21586
rect 27074 21534 27076 21586
rect 26908 21476 26964 21486
rect 26908 21382 26964 21420
rect 27020 21028 27076 21534
rect 27244 21588 27300 22540
rect 27356 21812 27412 24670
rect 27468 23268 27524 25004
rect 27692 23938 27748 25340
rect 27804 25396 27860 25406
rect 27804 25394 28196 25396
rect 27804 25342 27806 25394
rect 27858 25342 28196 25394
rect 27804 25340 28196 25342
rect 27804 25330 27860 25340
rect 28140 24946 28196 25340
rect 28252 25282 28308 25900
rect 28252 25230 28254 25282
rect 28306 25230 28308 25282
rect 28252 25172 28308 25230
rect 28252 25106 28308 25116
rect 28140 24894 28142 24946
rect 28194 24894 28196 24946
rect 28140 24882 28196 24894
rect 28028 24722 28084 24734
rect 28028 24670 28030 24722
rect 28082 24670 28084 24722
rect 28028 24052 28084 24670
rect 28252 24724 28308 24734
rect 28252 24630 28308 24668
rect 28364 24500 28420 26236
rect 27692 23886 27694 23938
rect 27746 23886 27748 23938
rect 27692 23874 27748 23886
rect 27804 23996 28084 24052
rect 28140 24444 28420 24500
rect 27804 23716 27860 23996
rect 28028 23826 28084 23838
rect 28028 23774 28030 23826
rect 28082 23774 28084 23826
rect 27804 23650 27860 23660
rect 27916 23714 27972 23726
rect 27916 23662 27918 23714
rect 27970 23662 27972 23714
rect 27916 23380 27972 23662
rect 27916 23314 27972 23324
rect 27804 23268 27860 23278
rect 27468 23266 27860 23268
rect 27468 23214 27806 23266
rect 27858 23214 27860 23266
rect 27468 23212 27860 23214
rect 27468 23042 27524 23054
rect 27468 22990 27470 23042
rect 27522 22990 27524 23042
rect 27468 22370 27524 22990
rect 27468 22318 27470 22370
rect 27522 22318 27524 22370
rect 27468 22306 27524 22318
rect 27804 21924 27860 23212
rect 27804 21858 27860 21868
rect 27916 23154 27972 23166
rect 27916 23102 27918 23154
rect 27970 23102 27972 23154
rect 27692 21812 27748 21822
rect 27356 21810 27748 21812
rect 27356 21758 27694 21810
rect 27746 21758 27748 21810
rect 27356 21756 27748 21758
rect 27692 21746 27748 21756
rect 27804 21700 27860 21710
rect 27804 21606 27860 21644
rect 27580 21588 27636 21598
rect 27244 21532 27412 21588
rect 26460 20822 26516 20860
rect 26908 20972 27076 21028
rect 27244 21364 27300 21374
rect 26236 20190 26238 20242
rect 26290 20190 26292 20242
rect 26236 20178 26292 20190
rect 26796 20468 26852 20478
rect 26236 20020 26292 20030
rect 26236 19926 26292 19964
rect 26460 20018 26516 20030
rect 26460 19966 26462 20018
rect 26514 19966 26516 20018
rect 26460 19684 26516 19966
rect 26460 19618 26516 19628
rect 26572 19348 26628 19358
rect 26348 19236 26404 19246
rect 26348 19142 26404 19180
rect 26572 19234 26628 19292
rect 26572 19182 26574 19234
rect 26626 19182 26628 19234
rect 26572 19170 26628 19182
rect 26460 19012 26516 19022
rect 26460 18918 26516 18956
rect 26796 19012 26852 20412
rect 26908 20132 26964 20972
rect 27132 20690 27188 20702
rect 27132 20638 27134 20690
rect 27186 20638 27188 20690
rect 27132 20132 27188 20638
rect 26908 20076 27076 20132
rect 26908 19906 26964 19918
rect 26908 19854 26910 19906
rect 26962 19854 26964 19906
rect 26908 19794 26964 19854
rect 26908 19742 26910 19794
rect 26962 19742 26964 19794
rect 26908 19730 26964 19742
rect 27020 19460 27076 20076
rect 27132 20066 27188 20076
rect 27244 19794 27300 21308
rect 27356 20242 27412 21532
rect 27580 20914 27636 21532
rect 27580 20862 27582 20914
rect 27634 20862 27636 20914
rect 27580 20850 27636 20862
rect 27692 21364 27748 21374
rect 27692 21252 27748 21308
rect 27916 21252 27972 23102
rect 28028 22260 28084 23774
rect 28140 22484 28196 24444
rect 28252 23716 28308 23726
rect 28252 22596 28308 23660
rect 28476 23380 28532 26236
rect 28588 26290 28644 26302
rect 28588 26238 28590 26290
rect 28642 26238 28644 26290
rect 28588 26180 28644 26238
rect 28644 26124 28756 26180
rect 28588 26114 28644 26124
rect 28588 24948 28644 24958
rect 28588 24722 28644 24892
rect 28588 24670 28590 24722
rect 28642 24670 28644 24722
rect 28588 24658 28644 24670
rect 28588 24164 28644 24174
rect 28700 24164 28756 26124
rect 28812 25282 28868 26852
rect 28812 25230 28814 25282
rect 28866 25230 28868 25282
rect 28812 24612 28868 25230
rect 28924 26516 28980 26526
rect 28924 24948 28980 26460
rect 29036 26180 29092 26190
rect 29036 26086 29092 26124
rect 29260 25284 29316 26852
rect 29484 26404 29540 26414
rect 29484 26310 29540 26348
rect 29260 25218 29316 25228
rect 29484 25282 29540 25294
rect 29484 25230 29486 25282
rect 29538 25230 29540 25282
rect 28924 24882 28980 24892
rect 29372 25172 29428 25182
rect 29260 24834 29316 24846
rect 29260 24782 29262 24834
rect 29314 24782 29316 24834
rect 28812 24546 28868 24556
rect 29148 24724 29204 24734
rect 29148 24610 29204 24668
rect 29148 24558 29150 24610
rect 29202 24558 29204 24610
rect 29148 24546 29204 24558
rect 29260 24612 29316 24782
rect 29260 24546 29316 24556
rect 29372 24500 29428 25116
rect 29484 24836 29540 25230
rect 29484 24770 29540 24780
rect 29484 24500 29540 24510
rect 29372 24498 29540 24500
rect 29372 24446 29486 24498
rect 29538 24446 29540 24498
rect 29372 24444 29540 24446
rect 28588 24162 29204 24164
rect 28588 24110 28590 24162
rect 28642 24110 29204 24162
rect 28588 24108 29204 24110
rect 28588 24098 28644 24108
rect 28700 23828 28756 23838
rect 28700 23734 28756 23772
rect 28700 23380 28756 23390
rect 28252 22530 28308 22540
rect 28364 23378 28756 23380
rect 28364 23326 28702 23378
rect 28754 23326 28756 23378
rect 28364 23324 28756 23326
rect 28140 22418 28196 22428
rect 28252 22260 28308 22270
rect 28028 22258 28308 22260
rect 28028 22206 28254 22258
rect 28306 22206 28308 22258
rect 28028 22204 28308 22206
rect 28252 22194 28308 22204
rect 28364 21586 28420 23324
rect 28700 23314 28756 23324
rect 28812 23380 28868 23390
rect 28364 21534 28366 21586
rect 28418 21534 28420 21586
rect 28028 21476 28084 21486
rect 28028 21382 28084 21420
rect 27692 21196 27972 21252
rect 27692 20802 27748 21196
rect 28252 20916 28308 20926
rect 27692 20750 27694 20802
rect 27746 20750 27748 20802
rect 27692 20738 27748 20750
rect 28140 20804 28196 20814
rect 27356 20190 27358 20242
rect 27410 20190 27412 20242
rect 27356 20178 27412 20190
rect 27468 20580 27524 20590
rect 27692 20580 27748 20590
rect 27244 19742 27246 19794
rect 27298 19742 27300 19794
rect 27244 19730 27300 19742
rect 27356 19460 27412 19470
rect 27020 19458 27412 19460
rect 27020 19406 27358 19458
rect 27410 19406 27412 19458
rect 27020 19404 27412 19406
rect 27020 19234 27076 19404
rect 27356 19394 27412 19404
rect 27020 19182 27022 19234
rect 27074 19182 27076 19234
rect 27020 19170 27076 19182
rect 27468 19122 27524 20524
rect 27468 19070 27470 19122
rect 27522 19070 27524 19122
rect 27468 19058 27524 19070
rect 27580 20524 27692 20580
rect 27580 19572 27636 20524
rect 27692 20514 27748 20524
rect 28140 20468 28196 20748
rect 28140 20402 28196 20412
rect 26796 18946 26852 18956
rect 27132 19012 27188 19022
rect 27020 18788 27076 18798
rect 26236 18676 26292 18686
rect 26236 18582 26292 18620
rect 27020 18674 27076 18732
rect 27020 18622 27022 18674
rect 27074 18622 27076 18674
rect 26572 18450 26628 18462
rect 26572 18398 26574 18450
rect 26626 18398 26628 18450
rect 26348 17668 26404 17678
rect 26236 17556 26292 17566
rect 26348 17556 26404 17612
rect 26460 17556 26516 17566
rect 26348 17554 26516 17556
rect 26348 17502 26462 17554
rect 26514 17502 26516 17554
rect 26348 17500 26516 17502
rect 26236 17462 26292 17500
rect 26460 17490 26516 17500
rect 26572 17556 26628 18398
rect 26572 17554 26852 17556
rect 26572 17502 26574 17554
rect 26626 17502 26852 17554
rect 26572 17500 26852 17502
rect 26572 17490 26628 17500
rect 26572 16996 26628 17006
rect 26572 16902 26628 16940
rect 26124 16158 26126 16210
rect 26178 16158 26180 16210
rect 26124 16146 26180 16158
rect 26460 16882 26516 16894
rect 26460 16830 26462 16882
rect 26514 16830 26516 16882
rect 26348 16100 26404 16110
rect 26460 16100 26516 16830
rect 26572 16660 26628 16670
rect 26572 16566 26628 16604
rect 26348 16098 26516 16100
rect 26348 16046 26350 16098
rect 26402 16046 26516 16098
rect 26348 16044 26516 16046
rect 26572 16100 26628 16110
rect 26012 15988 26068 15998
rect 26012 15894 26068 15932
rect 25788 15486 25790 15538
rect 25842 15486 25844 15538
rect 25788 15474 25844 15486
rect 25900 15316 25956 15326
rect 25900 13860 25956 15260
rect 26348 15202 26404 16044
rect 26572 16006 26628 16044
rect 26684 15764 26740 15774
rect 26348 15150 26350 15202
rect 26402 15150 26404 15202
rect 26348 15138 26404 15150
rect 26460 15426 26516 15438
rect 26460 15374 26462 15426
rect 26514 15374 26516 15426
rect 26124 15090 26180 15102
rect 26124 15038 26126 15090
rect 26178 15038 26180 15090
rect 26124 14756 26180 15038
rect 26236 14756 26292 14766
rect 26124 14754 26292 14756
rect 26124 14702 26238 14754
rect 26290 14702 26292 14754
rect 26124 14700 26292 14702
rect 26236 14690 26292 14700
rect 26460 14532 26516 15374
rect 26684 15426 26740 15708
rect 26684 15374 26686 15426
rect 26738 15374 26740 15426
rect 26684 15362 26740 15374
rect 25788 13858 25956 13860
rect 25788 13806 25902 13858
rect 25954 13806 25956 13858
rect 25788 13804 25956 13806
rect 25788 13634 25844 13804
rect 25900 13794 25956 13804
rect 26124 14476 26516 14532
rect 26572 15316 26628 15326
rect 25788 13582 25790 13634
rect 25842 13582 25844 13634
rect 25788 13570 25844 13582
rect 26012 12068 26068 12078
rect 26124 12068 26180 14476
rect 26572 14418 26628 15260
rect 26572 14366 26574 14418
rect 26626 14366 26628 14418
rect 26348 14306 26404 14318
rect 26348 14254 26350 14306
rect 26402 14254 26404 14306
rect 26348 13748 26404 14254
rect 26012 12066 26180 12068
rect 26012 12014 26014 12066
rect 26066 12014 26180 12066
rect 26012 12012 26180 12014
rect 26236 13692 26404 13748
rect 26236 12292 26292 13692
rect 26348 13522 26404 13534
rect 26348 13470 26350 13522
rect 26402 13470 26404 13522
rect 26348 13300 26404 13470
rect 26348 13234 26404 13244
rect 26460 12964 26516 12974
rect 26572 12964 26628 14366
rect 26460 12962 26628 12964
rect 26460 12910 26462 12962
rect 26514 12910 26628 12962
rect 26460 12908 26628 12910
rect 26460 12898 26516 12908
rect 26572 12740 26628 12750
rect 26460 12292 26516 12302
rect 26236 12290 26516 12292
rect 26236 12238 26462 12290
rect 26514 12238 26516 12290
rect 26236 12236 26516 12238
rect 26012 11954 26068 12012
rect 26012 11902 26014 11954
rect 26066 11902 26068 11954
rect 26012 11890 26068 11902
rect 26124 11620 26180 11630
rect 26124 11526 26180 11564
rect 25788 11396 25844 11406
rect 25788 11302 25844 11340
rect 26124 11172 26180 11182
rect 25676 10276 25732 10556
rect 25564 10220 25732 10276
rect 25788 10836 25844 10846
rect 25340 7970 25396 7980
rect 25452 9714 25508 9726
rect 25452 9662 25454 9714
rect 25506 9662 25508 9714
rect 25452 8372 25508 9662
rect 25564 8820 25620 10220
rect 25676 10052 25732 10062
rect 25788 10052 25844 10780
rect 26124 10834 26180 11116
rect 26124 10782 26126 10834
rect 26178 10782 26180 10834
rect 26124 10770 26180 10782
rect 25676 10050 25844 10052
rect 25676 9998 25678 10050
rect 25730 9998 25844 10050
rect 25676 9996 25844 9998
rect 26124 10052 26180 10062
rect 25676 9986 25732 9996
rect 25900 9828 25956 9838
rect 25900 9734 25956 9772
rect 26124 9826 26180 9996
rect 26124 9774 26126 9826
rect 26178 9774 26180 9826
rect 26124 9380 26180 9774
rect 25788 9324 26180 9380
rect 25788 9044 25844 9324
rect 25788 8950 25844 8988
rect 26012 9044 26068 9054
rect 26012 8950 26068 8988
rect 25900 8930 25956 8942
rect 25900 8878 25902 8930
rect 25954 8878 25956 8930
rect 25900 8820 25956 8878
rect 25564 8764 25956 8820
rect 25452 7476 25508 8316
rect 25564 8148 25620 8158
rect 25564 8054 25620 8092
rect 25676 7698 25732 8764
rect 25676 7646 25678 7698
rect 25730 7646 25732 7698
rect 25676 7634 25732 7646
rect 26124 8148 26180 8158
rect 26124 7924 26180 8092
rect 26124 7586 26180 7868
rect 26124 7534 26126 7586
rect 26178 7534 26180 7586
rect 26124 7522 26180 7534
rect 25452 7410 25508 7420
rect 25676 7476 25732 7486
rect 25228 6850 25284 6860
rect 24892 6526 24894 6578
rect 24946 6526 24948 6578
rect 24892 6514 24948 6526
rect 25228 6580 25284 6590
rect 25676 6580 25732 7420
rect 25228 6578 25732 6580
rect 25228 6526 25230 6578
rect 25282 6526 25678 6578
rect 25730 6526 25732 6578
rect 25228 6524 25732 6526
rect 24332 6018 24612 6020
rect 24332 5966 24334 6018
rect 24386 5966 24612 6018
rect 24332 5964 24612 5966
rect 23772 5906 23828 5918
rect 23772 5854 23774 5906
rect 23826 5854 23828 5906
rect 23660 5236 23716 5246
rect 23548 5234 23716 5236
rect 23548 5182 23662 5234
rect 23714 5182 23716 5234
rect 23548 5180 23716 5182
rect 23660 5170 23716 5180
rect 23436 4946 23492 4956
rect 23772 5012 23828 5854
rect 24332 5572 24388 5964
rect 24332 5506 24388 5516
rect 24668 5906 24724 5918
rect 24668 5854 24670 5906
rect 24722 5854 24724 5906
rect 23772 4946 23828 4956
rect 24108 5122 24164 5134
rect 24108 5070 24110 5122
rect 24162 5070 24164 5122
rect 24108 5012 24164 5070
rect 24108 4946 24164 4956
rect 24668 5012 24724 5854
rect 24668 4946 24724 4956
rect 24892 5122 24948 5134
rect 24892 5070 24894 5122
rect 24946 5070 24948 5122
rect 24892 5012 24948 5070
rect 23212 3714 23268 3724
rect 24332 3780 24388 3790
rect 20188 3614 20190 3666
rect 20242 3614 20244 3666
rect 18732 3502 18734 3554
rect 18786 3502 18788 3554
rect 18732 3490 18788 3502
rect 20188 3556 20244 3614
rect 20188 3490 20244 3500
rect 24332 3554 24388 3724
rect 24892 3668 24948 4956
rect 25228 4900 25284 6524
rect 25676 6514 25732 6524
rect 25788 6916 25844 6926
rect 25788 6244 25844 6860
rect 26124 6580 26180 6590
rect 26124 6486 26180 6524
rect 25564 6188 25844 6244
rect 25564 6130 25620 6188
rect 25564 6078 25566 6130
rect 25618 6078 25620 6130
rect 25564 6066 25620 6078
rect 25228 4834 25284 4844
rect 24892 3602 24948 3612
rect 25340 3780 25396 3790
rect 25340 3666 25396 3724
rect 25340 3614 25342 3666
rect 25394 3614 25396 3666
rect 25340 3602 25396 3614
rect 24332 3502 24334 3554
rect 24386 3502 24388 3554
rect 24332 3490 24388 3502
rect 13916 2884 13972 3164
rect 13916 2818 13972 2828
rect 17612 3442 17668 3454
rect 17612 3390 17614 3442
rect 17666 3390 17668 3442
rect 16828 924 17220 980
rect 16828 800 16884 924
rect 0 200 112 800
rect 5376 200 5488 800
rect 11424 200 11536 800
rect 16800 200 16912 800
rect 17164 756 17220 924
rect 17612 756 17668 3390
rect 23212 3442 23268 3454
rect 23212 3390 23214 3442
rect 23266 3390 23268 3442
rect 23212 3388 23268 3390
rect 26236 3388 26292 12236
rect 26460 12226 26516 12236
rect 26572 11844 26628 12684
rect 26684 12738 26740 12750
rect 26684 12686 26686 12738
rect 26738 12686 26740 12738
rect 26684 12628 26740 12686
rect 26684 12068 26740 12572
rect 26684 12002 26740 12012
rect 26460 11788 26628 11844
rect 26348 9828 26404 9838
rect 26460 9828 26516 11788
rect 26572 10052 26628 10062
rect 26796 10052 26852 17500
rect 27020 17332 27076 18622
rect 27020 17266 27076 17276
rect 27020 16996 27076 17006
rect 27020 16210 27076 16940
rect 27020 16158 27022 16210
rect 27074 16158 27076 16210
rect 27020 16146 27076 16158
rect 26908 15988 26964 15998
rect 26908 15148 26964 15932
rect 26908 15092 27076 15148
rect 27020 14306 27076 15092
rect 27020 14254 27022 14306
rect 27074 14254 27076 14306
rect 27020 13300 27076 14254
rect 27020 13234 27076 13244
rect 26572 10050 26852 10052
rect 26572 9998 26574 10050
rect 26626 9998 26852 10050
rect 26572 9996 26852 9998
rect 26908 11396 26964 11406
rect 26908 11170 26964 11340
rect 26908 11118 26910 11170
rect 26962 11118 26964 11170
rect 26572 9986 26628 9996
rect 26460 9772 26628 9828
rect 26348 9042 26404 9772
rect 26348 8990 26350 9042
rect 26402 8990 26404 9042
rect 26348 8978 26404 8990
rect 26460 9044 26516 9054
rect 26460 8146 26516 8988
rect 26460 8094 26462 8146
rect 26514 8094 26516 8146
rect 26460 8082 26516 8094
rect 26572 7924 26628 9772
rect 26908 9604 26964 11118
rect 27020 10948 27076 10958
rect 27020 10834 27076 10892
rect 27020 10782 27022 10834
rect 27074 10782 27076 10834
rect 27020 10770 27076 10782
rect 27132 10276 27188 18956
rect 27580 18674 27636 19516
rect 27692 20132 27748 20142
rect 27692 19124 27748 20076
rect 28140 20020 28196 20030
rect 28140 19926 28196 19964
rect 28252 19908 28308 20860
rect 28364 20244 28420 21534
rect 28364 20178 28420 20188
rect 28476 23156 28532 23166
rect 28476 22258 28532 23100
rect 28700 22596 28756 22606
rect 28588 22372 28644 22382
rect 28588 22278 28644 22316
rect 28476 22206 28478 22258
rect 28530 22206 28532 22258
rect 28476 21812 28532 22206
rect 28252 19842 28308 19852
rect 28476 19348 28532 21756
rect 28700 20690 28756 22540
rect 28700 20638 28702 20690
rect 28754 20638 28756 20690
rect 28700 20626 28756 20638
rect 28364 19292 28532 19348
rect 28588 19906 28644 19918
rect 28588 19854 28590 19906
rect 28642 19854 28644 19906
rect 27692 19030 27748 19068
rect 28028 19234 28084 19246
rect 28028 19182 28030 19234
rect 28082 19182 28084 19234
rect 27580 18622 27582 18674
rect 27634 18622 27636 18674
rect 27580 18610 27636 18622
rect 27916 18450 27972 18462
rect 27916 18398 27918 18450
rect 27970 18398 27972 18450
rect 27244 17892 27300 17902
rect 27244 17798 27300 17836
rect 27356 17668 27412 17678
rect 27244 17442 27300 17454
rect 27244 17390 27246 17442
rect 27298 17390 27300 17442
rect 27244 16548 27300 17390
rect 27356 16770 27412 17612
rect 27916 17444 27972 18398
rect 28028 18340 28084 19182
rect 28364 18676 28420 19292
rect 28364 18610 28420 18620
rect 28476 19122 28532 19134
rect 28476 19070 28478 19122
rect 28530 19070 28532 19122
rect 28028 18274 28084 18284
rect 28364 18452 28420 18462
rect 28364 18116 28420 18396
rect 28364 18050 28420 18060
rect 28476 17892 28532 19070
rect 28588 18788 28644 19854
rect 28812 19122 28868 23324
rect 29036 23156 29092 23166
rect 28924 21588 28980 21598
rect 28924 21494 28980 21532
rect 29036 20580 29092 23100
rect 29148 21588 29204 24108
rect 29484 23716 29540 24444
rect 29820 24164 29876 33628
rect 29932 33572 29988 34188
rect 30044 34178 30100 34188
rect 30156 34132 30212 34142
rect 30156 34038 30212 34076
rect 29932 33346 29988 33516
rect 29932 33294 29934 33346
rect 29986 33294 29988 33346
rect 29932 32452 29988 33294
rect 30268 33124 30324 33134
rect 30268 33030 30324 33068
rect 29932 32386 29988 32396
rect 30380 31106 30436 38612
rect 30716 38162 30772 38174
rect 30716 38110 30718 38162
rect 30770 38110 30772 38162
rect 30716 38052 30772 38110
rect 30716 37986 30772 37996
rect 30828 37826 30884 37838
rect 30828 37774 30830 37826
rect 30882 37774 30884 37826
rect 30828 37716 30884 37774
rect 30828 37268 30884 37660
rect 30828 37202 30884 37212
rect 30716 36260 30772 36270
rect 30492 36036 30548 36046
rect 30492 35922 30548 35980
rect 30492 35870 30494 35922
rect 30546 35870 30548 35922
rect 30492 35858 30548 35870
rect 30716 35698 30772 36204
rect 30940 35924 30996 38612
rect 31052 37940 31108 37950
rect 31052 37156 31108 37884
rect 31052 37062 31108 37100
rect 31164 37380 31220 37390
rect 31164 37154 31220 37324
rect 31164 37102 31166 37154
rect 31218 37102 31220 37154
rect 30940 35868 31108 35924
rect 30716 35646 30718 35698
rect 30770 35646 30772 35698
rect 30492 35588 30548 35598
rect 30492 32676 30548 35532
rect 30604 35586 30660 35598
rect 30604 35534 30606 35586
rect 30658 35534 30660 35586
rect 30604 35364 30660 35534
rect 30604 35298 30660 35308
rect 30716 34356 30772 35646
rect 30604 34300 30772 34356
rect 30940 34580 30996 34590
rect 30940 34354 30996 34524
rect 30940 34302 30942 34354
rect 30994 34302 30996 34354
rect 30604 33572 30660 34300
rect 30940 34290 30996 34302
rect 30604 33506 30660 33516
rect 30716 34130 30772 34142
rect 30716 34078 30718 34130
rect 30770 34078 30772 34130
rect 30716 33460 30772 34078
rect 30828 34132 30884 34142
rect 30828 34038 30884 34076
rect 30716 33394 30772 33404
rect 30828 33124 30884 33134
rect 30828 33030 30884 33068
rect 30492 32620 30660 32676
rect 30380 31054 30382 31106
rect 30434 31054 30436 31106
rect 30380 31042 30436 31054
rect 30492 32452 30548 32462
rect 29932 30994 29988 31006
rect 29932 30942 29934 30994
rect 29986 30942 29988 30994
rect 29932 30212 29988 30942
rect 30156 30882 30212 30894
rect 30492 30884 30548 32396
rect 30156 30830 30158 30882
rect 30210 30830 30212 30882
rect 30156 30436 30212 30830
rect 30156 30370 30212 30380
rect 30380 30828 30548 30884
rect 29932 29540 29988 30156
rect 30268 29540 30324 29550
rect 29932 29538 30324 29540
rect 29932 29486 30270 29538
rect 30322 29486 30324 29538
rect 29932 29484 30324 29486
rect 30268 29204 30324 29484
rect 30268 29138 30324 29148
rect 30268 28532 30324 28542
rect 30268 28438 30324 28476
rect 30156 27076 30212 27086
rect 30156 26982 30212 27020
rect 30268 26964 30324 27002
rect 30268 26898 30324 26908
rect 30380 26908 30436 30828
rect 30492 29986 30548 29998
rect 30492 29934 30494 29986
rect 30546 29934 30548 29986
rect 30492 29652 30548 29934
rect 30492 29586 30548 29596
rect 30604 29428 30660 32620
rect 30716 31554 30772 31566
rect 30716 31502 30718 31554
rect 30770 31502 30772 31554
rect 30716 30212 30772 31502
rect 30716 30146 30772 30156
rect 30940 30212 30996 30222
rect 30940 30118 30996 30156
rect 30828 30100 30884 30110
rect 30828 30006 30884 30044
rect 30716 29988 30772 29998
rect 30716 29894 30772 29932
rect 30492 29372 30660 29428
rect 30716 29764 30772 29774
rect 31052 29764 31108 35868
rect 31164 35588 31220 37102
rect 31276 36260 31332 36270
rect 31276 36166 31332 36204
rect 31164 35532 31332 35588
rect 31164 34356 31220 34366
rect 31164 34262 31220 34300
rect 31276 34132 31332 35532
rect 31164 34076 31332 34132
rect 31164 31332 31220 34076
rect 31388 32788 31444 38612
rect 31500 37828 31556 37838
rect 31500 37734 31556 37772
rect 31500 35698 31556 35710
rect 31500 35646 31502 35698
rect 31554 35646 31556 35698
rect 31500 35588 31556 35646
rect 31500 35522 31556 35532
rect 31612 35476 31668 38612
rect 31724 37826 31780 39678
rect 31948 39284 32004 39294
rect 31836 37940 31892 37950
rect 31836 37846 31892 37884
rect 31724 37774 31726 37826
rect 31778 37774 31780 37826
rect 31724 37716 31780 37774
rect 31724 37650 31780 37660
rect 31836 37268 31892 37278
rect 31836 37174 31892 37212
rect 31948 36036 32004 39228
rect 32060 37156 32116 47628
rect 32172 44994 32228 45006
rect 32172 44942 32174 44994
rect 32226 44942 32228 44994
rect 32172 44212 32228 44942
rect 32172 44118 32228 44156
rect 32284 43650 32340 50372
rect 32508 50372 32564 50382
rect 32508 49700 32564 50316
rect 32396 49698 32564 49700
rect 32396 49646 32510 49698
rect 32562 49646 32564 49698
rect 32396 49644 32564 49646
rect 32396 49028 32452 49644
rect 32508 49634 32564 49644
rect 32396 48934 32452 48972
rect 32508 48020 32564 48030
rect 32508 47926 32564 47964
rect 32620 47348 32676 51886
rect 33628 51380 33684 51996
rect 33740 51380 33796 51390
rect 33628 51378 33796 51380
rect 33628 51326 33742 51378
rect 33794 51326 33796 51378
rect 33628 51324 33796 51326
rect 33740 51314 33796 51324
rect 32732 51154 32788 51166
rect 32732 51102 32734 51154
rect 32786 51102 32788 51154
rect 32732 50820 32788 51102
rect 32732 50754 32788 50764
rect 33068 50370 33124 50382
rect 33068 50318 33070 50370
rect 33122 50318 33124 50370
rect 33068 49700 33124 50318
rect 33516 50372 33572 50382
rect 33516 50278 33572 50316
rect 33068 49634 33124 49644
rect 33740 49924 33796 49934
rect 33628 49588 33684 49598
rect 33292 49586 33684 49588
rect 33292 49534 33630 49586
rect 33682 49534 33684 49586
rect 33292 49532 33684 49534
rect 32732 49252 32788 49262
rect 32732 48466 32788 49196
rect 33292 49250 33348 49532
rect 33628 49522 33684 49532
rect 33292 49198 33294 49250
rect 33346 49198 33348 49250
rect 33292 49186 33348 49198
rect 33740 49138 33796 49868
rect 33964 49588 34020 49598
rect 33740 49086 33742 49138
rect 33794 49086 33796 49138
rect 33516 49028 33572 49038
rect 32732 48414 32734 48466
rect 32786 48414 32788 48466
rect 32732 48402 32788 48414
rect 32844 49026 33572 49028
rect 32844 48974 33518 49026
rect 33570 48974 33572 49026
rect 32844 48972 33572 48974
rect 32844 48130 32900 48972
rect 33516 48962 33572 48972
rect 33628 49028 33684 49038
rect 33628 48692 33684 48972
rect 33740 48916 33796 49086
rect 33740 48850 33796 48860
rect 33852 49586 34020 49588
rect 33852 49534 33966 49586
rect 34018 49534 34020 49586
rect 33852 49532 34020 49534
rect 33628 48636 33796 48692
rect 32844 48078 32846 48130
rect 32898 48078 32900 48130
rect 32844 48066 32900 48078
rect 33628 48132 33684 48142
rect 33292 48020 33348 48030
rect 33292 47458 33348 47964
rect 33292 47406 33294 47458
rect 33346 47406 33348 47458
rect 33292 47394 33348 47406
rect 32620 47282 32676 47292
rect 33628 47348 33684 48076
rect 33740 48020 33796 48636
rect 33852 48244 33908 49532
rect 33964 49522 34020 49532
rect 34076 49588 34132 52332
rect 34188 52164 34244 52174
rect 34188 51380 34244 52108
rect 34188 51286 34244 51324
rect 34076 49028 34132 49532
rect 34188 49698 34244 49710
rect 34188 49646 34190 49698
rect 34242 49646 34244 49698
rect 34188 49252 34244 49646
rect 34188 49186 34244 49196
rect 34188 49028 34244 49038
rect 34076 49026 34244 49028
rect 34076 48974 34190 49026
rect 34242 48974 34244 49026
rect 34076 48972 34244 48974
rect 34188 48962 34244 48972
rect 34300 48916 34356 52668
rect 34412 50148 34468 55022
rect 37548 54628 37604 54638
rect 37660 54628 37716 55244
rect 37772 55234 37828 55244
rect 39676 55298 40068 55300
rect 39676 55246 39790 55298
rect 39842 55246 40068 55298
rect 39676 55244 40068 55246
rect 40236 55300 40292 55310
rect 40572 55300 40628 55412
rect 40236 55298 40628 55300
rect 40236 55246 40238 55298
rect 40290 55246 40628 55298
rect 40236 55244 40628 55246
rect 39340 55188 39396 55198
rect 37548 54626 37716 54628
rect 37548 54574 37550 54626
rect 37602 54574 37716 54626
rect 37548 54572 37716 54574
rect 39228 55186 39396 55188
rect 39228 55134 39342 55186
rect 39394 55134 39396 55186
rect 39228 55132 39396 55134
rect 37548 54562 37604 54572
rect 38220 54516 38276 54526
rect 38220 54422 38276 54460
rect 39116 54516 39172 54526
rect 38444 54404 38500 54414
rect 38444 54310 38500 54348
rect 39004 54404 39060 54414
rect 35196 54124 35460 54134
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35196 54058 35460 54068
rect 39004 53730 39060 54348
rect 39004 53678 39006 53730
rect 39058 53678 39060 53730
rect 35980 53620 36036 53630
rect 35084 53172 35140 53182
rect 34860 53116 35084 53172
rect 34748 52836 34804 52846
rect 34748 52742 34804 52780
rect 34860 52388 34916 53116
rect 35084 53078 35140 53116
rect 35980 53172 36036 53564
rect 35980 53040 36036 53116
rect 38892 53058 38948 53070
rect 38892 53006 38894 53058
rect 38946 53006 38948 53058
rect 34860 52256 34916 52332
rect 34972 52836 35028 52846
rect 34972 52276 35028 52780
rect 35644 52836 35700 52846
rect 35644 52742 35700 52780
rect 36540 52834 36596 52846
rect 38332 52836 38388 52846
rect 36540 52782 36542 52834
rect 36594 52782 36596 52834
rect 35196 52556 35460 52566
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35196 52490 35460 52500
rect 35084 52276 35140 52286
rect 35028 52274 35140 52276
rect 35028 52222 35086 52274
rect 35138 52222 35140 52274
rect 35028 52220 35140 52222
rect 34972 52144 35028 52220
rect 35084 52210 35140 52220
rect 36316 52276 36372 52286
rect 34524 52052 34580 52062
rect 34524 51958 34580 51996
rect 35868 52052 35924 52062
rect 35308 51380 35364 51390
rect 35868 51380 35924 51996
rect 36092 52050 36148 52062
rect 36092 51998 36094 52050
rect 36146 51998 36148 52050
rect 36092 51940 36148 51998
rect 36092 51874 36148 51884
rect 36204 52050 36260 52062
rect 36204 51998 36206 52050
rect 36258 51998 36260 52050
rect 36092 51380 36148 51390
rect 35868 51378 36148 51380
rect 35868 51326 36094 51378
rect 36146 51326 36148 51378
rect 35868 51324 36148 51326
rect 35308 51286 35364 51324
rect 34636 51268 34692 51278
rect 34636 51174 34692 51212
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35196 50922 35460 50932
rect 36092 50596 36148 51324
rect 36092 50502 36148 50540
rect 34748 50484 34804 50494
rect 34748 50390 34804 50428
rect 35196 50484 35252 50494
rect 36204 50428 36260 51998
rect 36316 50818 36372 52220
rect 36428 52162 36484 52174
rect 36428 52110 36430 52162
rect 36482 52110 36484 52162
rect 36428 51604 36484 52110
rect 36540 52052 36596 52782
rect 38108 52834 38388 52836
rect 38108 52782 38334 52834
rect 38386 52782 38388 52834
rect 38108 52780 38388 52782
rect 37884 52724 37940 52734
rect 36652 52276 36708 52286
rect 36652 52182 36708 52220
rect 36540 51986 36596 51996
rect 37436 52162 37492 52174
rect 37436 52110 37438 52162
rect 37490 52110 37492 52162
rect 37436 51940 37492 52110
rect 37436 51874 37492 51884
rect 37884 51938 37940 52668
rect 37884 51886 37886 51938
rect 37938 51886 37940 51938
rect 37548 51604 37604 51614
rect 36428 51548 36596 51604
rect 36316 50766 36318 50818
rect 36370 50766 36372 50818
rect 36316 50754 36372 50766
rect 36428 51380 36484 51390
rect 35196 50390 35252 50428
rect 35644 50372 35700 50382
rect 35532 50370 35700 50372
rect 35532 50318 35646 50370
rect 35698 50318 35700 50370
rect 35532 50316 35700 50318
rect 34412 50092 35028 50148
rect 34524 49028 34580 49038
rect 34300 48860 34468 48916
rect 33964 48804 34020 48814
rect 33964 48710 34020 48748
rect 34076 48802 34132 48814
rect 34076 48750 34078 48802
rect 34130 48750 34132 48802
rect 34076 48244 34132 48750
rect 33852 48188 34020 48244
rect 33852 48020 33908 48030
rect 33740 48018 33908 48020
rect 33740 47966 33854 48018
rect 33906 47966 33908 48018
rect 33740 47964 33908 47966
rect 33852 47908 33908 47964
rect 33964 48020 34020 48188
rect 34076 48178 34132 48188
rect 34076 48020 34132 48030
rect 34020 48018 34132 48020
rect 34020 47966 34078 48018
rect 34130 47966 34132 48018
rect 34020 47964 34132 47966
rect 33964 47888 34020 47964
rect 34076 47954 34132 47964
rect 33740 47796 33796 47806
rect 33740 47570 33796 47740
rect 33740 47518 33742 47570
rect 33794 47518 33796 47570
rect 33740 47506 33796 47518
rect 33628 47254 33684 47292
rect 33852 47346 33908 47852
rect 33852 47294 33854 47346
rect 33906 47294 33908 47346
rect 33852 47282 33908 47294
rect 34300 47348 34356 47358
rect 34300 47254 34356 47292
rect 34412 47236 34468 48860
rect 34524 48466 34580 48972
rect 34860 48916 34916 48926
rect 34524 48414 34526 48466
rect 34578 48414 34580 48466
rect 34524 48402 34580 48414
rect 34636 48914 34916 48916
rect 34636 48862 34862 48914
rect 34914 48862 34916 48914
rect 34636 48860 34916 48862
rect 34636 48244 34692 48860
rect 34860 48850 34916 48860
rect 34524 48188 34692 48244
rect 34748 48692 34804 48702
rect 34972 48692 35028 50092
rect 35532 49812 35588 50316
rect 35644 50306 35700 50316
rect 36092 50372 36260 50428
rect 36316 50372 36372 50382
rect 36092 49922 36148 50372
rect 36092 49870 36094 49922
rect 36146 49870 36148 49922
rect 36092 49858 36148 49870
rect 35532 49756 36036 49812
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35084 49028 35140 49038
rect 35084 48934 35140 48972
rect 35532 49026 35588 49756
rect 35980 49700 36036 49756
rect 36204 49810 36260 49822
rect 36204 49758 36206 49810
rect 36258 49758 36260 49810
rect 36204 49700 36260 49758
rect 35980 49644 36260 49700
rect 35644 49588 35700 49598
rect 35644 49494 35700 49532
rect 35532 48974 35534 49026
rect 35586 48974 35588 49026
rect 35532 48962 35588 48974
rect 35868 48916 35924 48926
rect 35196 48804 35252 48814
rect 35196 48710 35252 48748
rect 35308 48802 35364 48814
rect 35308 48750 35310 48802
rect 35362 48750 35364 48802
rect 34524 47796 34580 48188
rect 34748 48132 34804 48636
rect 34860 48636 35028 48692
rect 34860 48468 34916 48636
rect 35084 48580 35140 48590
rect 34860 48412 35028 48468
rect 34524 47730 34580 47740
rect 34636 48076 34804 48132
rect 34860 48130 34916 48142
rect 34860 48078 34862 48130
rect 34914 48078 34916 48130
rect 34636 47348 34692 48076
rect 34748 47908 34804 47918
rect 34748 47682 34804 47852
rect 34748 47630 34750 47682
rect 34802 47630 34804 47682
rect 34748 47570 34804 47630
rect 34748 47518 34750 47570
rect 34802 47518 34804 47570
rect 34748 47506 34804 47518
rect 34860 47572 34916 48078
rect 34860 47506 34916 47516
rect 34636 47292 34916 47348
rect 34412 47180 34804 47236
rect 33964 46900 34020 46910
rect 33740 46788 33796 46798
rect 33796 46732 33908 46788
rect 33740 46694 33796 46732
rect 32396 46676 32452 46686
rect 32396 43764 32452 46620
rect 32508 46564 32564 46574
rect 32508 46470 32564 46508
rect 33628 46564 33684 46574
rect 33628 46470 33684 46508
rect 33068 45666 33124 45678
rect 33068 45614 33070 45666
rect 33122 45614 33124 45666
rect 32620 45106 32676 45118
rect 33068 45108 33124 45614
rect 32620 45054 32622 45106
rect 32674 45054 32676 45106
rect 32620 43988 32676 45054
rect 32620 43922 32676 43932
rect 32732 45052 33124 45108
rect 33628 45666 33684 45678
rect 33628 45614 33630 45666
rect 33682 45614 33684 45666
rect 32732 44212 32788 45052
rect 32732 44098 32788 44156
rect 33628 44324 33684 45614
rect 33740 45444 33796 45454
rect 33740 45106 33796 45388
rect 33740 45054 33742 45106
rect 33794 45054 33796 45106
rect 33740 45042 33796 45054
rect 32732 44046 32734 44098
rect 32786 44046 32788 44098
rect 32396 43708 32676 43764
rect 32284 43598 32286 43650
rect 32338 43598 32340 43650
rect 32284 43540 32340 43598
rect 32284 43474 32340 43484
rect 32620 42980 32676 43708
rect 32732 43316 32788 44046
rect 32844 44100 32900 44110
rect 32844 44006 32900 44044
rect 32956 44098 33012 44110
rect 32956 44046 32958 44098
rect 33010 44046 33012 44098
rect 32956 43988 33012 44046
rect 33180 44100 33236 44110
rect 33180 44006 33236 44044
rect 32956 43922 33012 43932
rect 33628 43764 33684 44268
rect 33516 43708 33684 43764
rect 33516 43540 33572 43708
rect 33068 43484 33572 43540
rect 32844 43428 32900 43438
rect 32844 43426 33012 43428
rect 32844 43374 32846 43426
rect 32898 43374 33012 43426
rect 32844 43372 33012 43374
rect 32844 43362 32900 43372
rect 32732 43250 32788 43260
rect 32396 42924 32676 42980
rect 32396 42868 32452 42924
rect 32284 42812 32452 42868
rect 32284 41860 32340 42812
rect 32508 42756 32564 42766
rect 32396 42084 32452 42094
rect 32508 42084 32564 42700
rect 32732 42756 32788 42766
rect 32732 42662 32788 42700
rect 32620 42644 32676 42654
rect 32620 42550 32676 42588
rect 32956 42532 33012 43372
rect 32956 42438 33012 42476
rect 32396 42082 32564 42084
rect 32396 42030 32398 42082
rect 32450 42030 32564 42082
rect 32396 42028 32564 42030
rect 32396 42018 32452 42028
rect 32284 41804 32452 41860
rect 32284 39618 32340 39630
rect 32284 39566 32286 39618
rect 32338 39566 32340 39618
rect 32284 39060 32340 39566
rect 32284 38994 32340 39004
rect 32396 38668 32452 41804
rect 32956 39620 33012 39630
rect 32844 39508 32900 39518
rect 32844 39414 32900 39452
rect 32956 38668 33012 39564
rect 32060 37090 32116 37100
rect 32172 38612 32452 38668
rect 32844 38612 33012 38668
rect 32172 36932 32228 38612
rect 32396 37826 32452 37838
rect 32732 37828 32788 37838
rect 32396 37774 32398 37826
rect 32450 37774 32452 37826
rect 32396 37380 32452 37774
rect 32396 37314 32452 37324
rect 32620 37826 32788 37828
rect 32620 37774 32734 37826
rect 32786 37774 32788 37826
rect 32620 37772 32788 37774
rect 32620 37380 32676 37772
rect 32732 37762 32788 37772
rect 32620 37286 32676 37324
rect 32732 37378 32788 37390
rect 32732 37326 32734 37378
rect 32786 37326 32788 37378
rect 32732 37268 32788 37326
rect 32732 37202 32788 37212
rect 31948 35970 32004 35980
rect 32060 36876 32228 36932
rect 31836 35924 31892 35934
rect 31836 35830 31892 35868
rect 31612 35410 31668 35420
rect 31836 34692 31892 34702
rect 31836 34598 31892 34636
rect 31724 34580 31780 34590
rect 31724 34356 31780 34524
rect 31724 34354 31892 34356
rect 31724 34302 31726 34354
rect 31778 34302 31892 34354
rect 31724 34300 31892 34302
rect 31724 34290 31780 34300
rect 31388 32732 31668 32788
rect 31500 32564 31556 32574
rect 31388 32562 31556 32564
rect 31388 32510 31502 32562
rect 31554 32510 31556 32562
rect 31388 32508 31556 32510
rect 31388 31892 31444 32508
rect 31500 32498 31556 32508
rect 31164 31266 31220 31276
rect 31276 31666 31332 31678
rect 31276 31614 31278 31666
rect 31330 31614 31332 31666
rect 30716 29426 30772 29708
rect 30716 29374 30718 29426
rect 30770 29374 30772 29426
rect 30492 28420 30548 29372
rect 30716 29362 30772 29374
rect 30940 29708 31108 29764
rect 31164 31108 31220 31118
rect 31276 31108 31332 31614
rect 31164 31106 31332 31108
rect 31164 31054 31166 31106
rect 31218 31054 31332 31106
rect 31164 31052 31332 31054
rect 31388 31554 31444 31836
rect 31388 31502 31390 31554
rect 31442 31502 31444 31554
rect 31388 31108 31444 31502
rect 31164 30098 31220 31052
rect 31388 31042 31444 31052
rect 31500 31220 31556 31230
rect 31500 31106 31556 31164
rect 31500 31054 31502 31106
rect 31554 31054 31556 31106
rect 31500 31042 31556 31054
rect 31164 30046 31166 30098
rect 31218 30046 31220 30098
rect 30828 29314 30884 29326
rect 30828 29262 30830 29314
rect 30882 29262 30884 29314
rect 30604 28644 30660 28654
rect 30604 28550 30660 28588
rect 30492 28364 30772 28420
rect 30604 27858 30660 27870
rect 30604 27806 30606 27858
rect 30658 27806 30660 27858
rect 30492 27076 30548 27086
rect 30604 27076 30660 27806
rect 30492 27074 30660 27076
rect 30492 27022 30494 27074
rect 30546 27022 30660 27074
rect 30492 27020 30660 27022
rect 30492 27010 30548 27020
rect 30380 26852 30660 26908
rect 30044 26178 30100 26190
rect 30044 26126 30046 26178
rect 30098 26126 30100 26178
rect 30044 26068 30100 26126
rect 30044 26002 30100 26012
rect 29932 25282 29988 25294
rect 29932 25230 29934 25282
rect 29986 25230 29988 25282
rect 29932 24948 29988 25230
rect 29932 24612 29988 24892
rect 29932 24610 30100 24612
rect 29932 24558 29934 24610
rect 29986 24558 30100 24610
rect 29932 24556 30100 24558
rect 29932 24546 29988 24556
rect 29820 24098 29876 24108
rect 29484 23622 29540 23660
rect 29708 23828 29764 23838
rect 29484 23380 29540 23390
rect 29484 23286 29540 23324
rect 29372 22596 29428 22606
rect 29148 21532 29316 21588
rect 29036 20514 29092 20524
rect 29148 21362 29204 21374
rect 29148 21310 29150 21362
rect 29202 21310 29204 21362
rect 29036 20132 29092 20142
rect 29036 20038 29092 20076
rect 28812 19070 28814 19122
rect 28866 19070 28868 19122
rect 28812 19058 28868 19070
rect 29148 18788 29204 21310
rect 28588 18732 29204 18788
rect 28924 18564 28980 18574
rect 28476 17826 28532 17836
rect 28700 18452 28756 18462
rect 28252 17780 28308 17790
rect 28252 17666 28308 17724
rect 28252 17614 28254 17666
rect 28306 17614 28308 17666
rect 28252 17602 28308 17614
rect 28588 17780 28644 17790
rect 27972 17388 28196 17444
rect 27916 17350 27972 17388
rect 28140 17106 28196 17388
rect 28140 17054 28142 17106
rect 28194 17054 28196 17106
rect 28140 17042 28196 17054
rect 28252 17332 28308 17342
rect 28028 16996 28084 17006
rect 27356 16718 27358 16770
rect 27410 16718 27412 16770
rect 27356 16706 27412 16718
rect 27692 16882 27748 16894
rect 27692 16830 27694 16882
rect 27746 16830 27748 16882
rect 27692 16548 27748 16830
rect 27244 16492 27748 16548
rect 27244 15316 27300 15326
rect 27244 15222 27300 15260
rect 27468 15204 27524 15214
rect 27356 13746 27412 13758
rect 27356 13694 27358 13746
rect 27410 13694 27412 13746
rect 27356 13636 27412 13694
rect 27356 13570 27412 13580
rect 27356 13186 27412 13198
rect 27356 13134 27358 13186
rect 27410 13134 27412 13186
rect 27356 13074 27412 13134
rect 27356 13022 27358 13074
rect 27410 13022 27412 13074
rect 27356 13010 27412 13022
rect 27468 12740 27524 15148
rect 27580 14308 27636 14318
rect 27692 14308 27748 16492
rect 27916 16436 27972 16446
rect 27916 16098 27972 16380
rect 27916 16046 27918 16098
rect 27970 16046 27972 16098
rect 27916 16034 27972 16046
rect 28028 15538 28084 16940
rect 28252 16210 28308 17276
rect 28252 16158 28254 16210
rect 28306 16158 28308 16210
rect 28252 15652 28308 16158
rect 28252 15586 28308 15596
rect 28588 17106 28644 17724
rect 28588 17054 28590 17106
rect 28642 17054 28644 17106
rect 28028 15486 28030 15538
rect 28082 15486 28084 15538
rect 27804 15316 27860 15326
rect 27804 15222 27860 15260
rect 28028 15148 28084 15486
rect 28588 15316 28644 17054
rect 28028 15092 28196 15148
rect 27580 14306 27748 14308
rect 27580 14254 27582 14306
rect 27634 14254 27748 14306
rect 27580 14252 27748 14254
rect 27580 14242 27636 14252
rect 27468 12684 27636 12740
rect 27580 12402 27636 12684
rect 27580 12350 27582 12402
rect 27634 12350 27636 12402
rect 27580 12338 27636 12350
rect 27468 12292 27524 12302
rect 27468 12198 27524 12236
rect 27692 12180 27748 14252
rect 27916 14308 27972 14318
rect 27916 14214 27972 14252
rect 28140 13748 28196 15092
rect 28476 14308 28532 14318
rect 28252 13748 28308 13758
rect 28140 13746 28308 13748
rect 28140 13694 28254 13746
rect 28306 13694 28308 13746
rect 28140 13692 28308 13694
rect 27804 13636 27860 13646
rect 27804 12740 27860 13580
rect 28140 13186 28196 13692
rect 28252 13682 28308 13692
rect 28476 13746 28532 14252
rect 28476 13694 28478 13746
rect 28530 13694 28532 13746
rect 28252 13524 28308 13534
rect 28252 13430 28308 13468
rect 28140 13134 28142 13186
rect 28194 13134 28196 13186
rect 27804 12738 27972 12740
rect 27804 12686 27806 12738
rect 27858 12686 27972 12738
rect 27804 12684 27972 12686
rect 27804 12674 27860 12684
rect 27580 12124 27748 12180
rect 27244 11394 27300 11406
rect 27244 11342 27246 11394
rect 27298 11342 27300 11394
rect 27244 11284 27300 11342
rect 27244 10836 27300 11228
rect 27244 10612 27300 10780
rect 27468 11394 27524 11406
rect 27468 11342 27470 11394
rect 27522 11342 27524 11394
rect 27468 10724 27524 11342
rect 27580 10948 27636 12124
rect 27692 11956 27748 11966
rect 27916 11956 27972 12684
rect 27692 11954 27972 11956
rect 27692 11902 27694 11954
rect 27746 11902 27972 11954
rect 27692 11900 27972 11902
rect 27692 11890 27748 11900
rect 27580 10892 27860 10948
rect 27580 10724 27636 10734
rect 27468 10722 27636 10724
rect 27468 10670 27582 10722
rect 27634 10670 27636 10722
rect 27468 10668 27636 10670
rect 27356 10612 27412 10622
rect 27244 10610 27412 10612
rect 27244 10558 27358 10610
rect 27410 10558 27412 10610
rect 27244 10556 27412 10558
rect 27356 10546 27412 10556
rect 27132 10220 27300 10276
rect 27132 10052 27188 10062
rect 27020 9828 27076 9838
rect 27020 9734 27076 9772
rect 26908 9548 27076 9604
rect 26908 9044 26964 9054
rect 26908 8950 26964 8988
rect 22876 3332 23268 3388
rect 26012 3332 26292 3388
rect 26348 7868 26628 7924
rect 26684 8258 26740 8270
rect 26684 8206 26686 8258
rect 26738 8206 26740 8258
rect 26684 8036 26740 8206
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 22876 800 22932 3332
rect 26012 2548 26068 3332
rect 26348 2660 26404 7868
rect 26460 7588 26516 7598
rect 26684 7588 26740 7980
rect 26908 7924 26964 7934
rect 26908 7698 26964 7868
rect 26908 7646 26910 7698
rect 26962 7646 26964 7698
rect 26908 7634 26964 7646
rect 26460 7586 26740 7588
rect 26460 7534 26462 7586
rect 26514 7534 26740 7586
rect 26460 7532 26740 7534
rect 26460 7476 26516 7532
rect 26460 7410 26516 7420
rect 26908 7140 26964 7150
rect 26572 6468 26628 6478
rect 26572 6374 26628 6412
rect 26348 2594 26404 2604
rect 26012 2482 26068 2492
rect 26908 2324 26964 7084
rect 27020 3332 27076 9548
rect 27132 9042 27188 9996
rect 27132 8990 27134 9042
rect 27186 8990 27188 9042
rect 27132 8978 27188 8990
rect 27244 8820 27300 10220
rect 27356 9940 27412 9950
rect 27356 9714 27412 9884
rect 27356 9662 27358 9714
rect 27410 9662 27412 9714
rect 27356 9650 27412 9662
rect 27468 9044 27524 10668
rect 27580 10658 27636 10668
rect 27804 10276 27860 10892
rect 27468 8978 27524 8988
rect 27580 10220 27860 10276
rect 27468 8820 27524 8830
rect 27244 8818 27524 8820
rect 27244 8766 27470 8818
rect 27522 8766 27524 8818
rect 27244 8764 27524 8766
rect 27244 8036 27300 8046
rect 27244 7942 27300 7980
rect 27356 5124 27412 8764
rect 27468 8754 27524 8764
rect 27356 5058 27412 5068
rect 27020 3266 27076 3276
rect 26908 2258 26964 2268
rect 27580 1428 27636 10220
rect 27916 10164 27972 11900
rect 28028 11508 28084 11518
rect 28028 11414 28084 11452
rect 28140 11284 28196 13134
rect 28364 13188 28420 13198
rect 28476 13188 28532 13694
rect 28364 13186 28532 13188
rect 28364 13134 28366 13186
rect 28418 13134 28532 13186
rect 28364 13132 28532 13134
rect 28364 13122 28420 13132
rect 28476 12852 28532 12862
rect 28364 12796 28476 12852
rect 28364 11394 28420 12796
rect 28476 12758 28532 12796
rect 28588 12402 28644 15260
rect 28700 14420 28756 18396
rect 28924 18450 28980 18508
rect 28924 18398 28926 18450
rect 28978 18398 28980 18450
rect 28924 18386 28980 18398
rect 28812 17442 28868 17454
rect 28812 17390 28814 17442
rect 28866 17390 28868 17442
rect 28812 16884 28868 17390
rect 28812 16818 28868 16828
rect 28924 17444 28980 17454
rect 28924 16548 28980 17388
rect 28924 16482 28980 16492
rect 28812 16436 28868 16446
rect 28812 16210 28868 16380
rect 28812 16158 28814 16210
rect 28866 16158 28868 16210
rect 28812 16146 28868 16158
rect 28812 15316 28868 15326
rect 28812 15222 28868 15260
rect 28812 14420 28868 14430
rect 28700 14418 28868 14420
rect 28700 14366 28814 14418
rect 28866 14366 28868 14418
rect 28700 14364 28868 14366
rect 28812 14354 28868 14364
rect 28588 12350 28590 12402
rect 28642 12350 28644 12402
rect 28364 11342 28366 11394
rect 28418 11342 28420 11394
rect 28364 11330 28420 11342
rect 28476 12292 28532 12302
rect 28028 11228 28196 11284
rect 28028 10388 28084 11228
rect 28252 11172 28308 11182
rect 28140 10612 28196 10622
rect 28140 10518 28196 10556
rect 28028 10332 28196 10388
rect 27804 10108 27972 10164
rect 27804 9604 27860 10108
rect 27804 9602 28084 9604
rect 27804 9550 27806 9602
rect 27858 9550 28084 9602
rect 27804 9548 28084 9550
rect 27804 9538 27860 9548
rect 27916 8930 27972 8942
rect 27916 8878 27918 8930
rect 27970 8878 27972 8930
rect 27916 8818 27972 8878
rect 27916 8766 27918 8818
rect 27970 8766 27972 8818
rect 27916 8754 27972 8766
rect 27692 8034 27748 8046
rect 27692 7982 27694 8034
rect 27746 7982 27748 8034
rect 27692 7924 27748 7982
rect 27692 7858 27748 7868
rect 28028 6804 28084 9548
rect 28028 6738 28084 6748
rect 28028 4898 28084 4910
rect 28028 4846 28030 4898
rect 28082 4846 28084 4898
rect 28028 4004 28084 4846
rect 28140 4564 28196 10332
rect 28252 9938 28308 11116
rect 28476 10948 28532 12236
rect 28252 9886 28254 9938
rect 28306 9886 28308 9938
rect 28252 8818 28308 9886
rect 28364 10892 28532 10948
rect 28588 11506 28644 12350
rect 28924 12180 28980 12190
rect 28924 12086 28980 12124
rect 28588 11454 28590 11506
rect 28642 11454 28644 11506
rect 28364 9940 28420 10892
rect 28588 10836 28644 11454
rect 29036 11396 29092 18732
rect 29260 17668 29316 21532
rect 29372 20916 29428 22540
rect 29596 22482 29652 22494
rect 29596 22430 29598 22482
rect 29650 22430 29652 22482
rect 29596 22372 29652 22430
rect 29596 22306 29652 22316
rect 29484 21364 29540 21374
rect 29484 21270 29540 21308
rect 29708 21140 29764 23772
rect 29932 23828 29988 23838
rect 29932 23734 29988 23772
rect 29596 21084 29764 21140
rect 29820 23716 29876 23726
rect 29484 20916 29540 20926
rect 29372 20914 29540 20916
rect 29372 20862 29486 20914
rect 29538 20862 29540 20914
rect 29372 20860 29540 20862
rect 29484 20850 29540 20860
rect 29596 20132 29652 21084
rect 29484 20076 29652 20132
rect 29820 20132 29876 23660
rect 29932 23156 29988 23166
rect 29932 23062 29988 23100
rect 29932 22596 29988 22606
rect 29932 22502 29988 22540
rect 30044 22484 30100 24556
rect 30380 24610 30436 24622
rect 30380 24558 30382 24610
rect 30434 24558 30436 24610
rect 30380 24388 30436 24558
rect 30436 24332 30548 24388
rect 30380 24322 30436 24332
rect 30044 22428 30324 22484
rect 30156 22260 30212 22270
rect 30156 22166 30212 22204
rect 30268 21812 30324 22428
rect 30268 21756 30436 21812
rect 30044 21700 30100 21710
rect 30044 21606 30100 21644
rect 30268 21586 30324 21598
rect 30268 21534 30270 21586
rect 30322 21534 30324 21586
rect 30268 20802 30324 21534
rect 30268 20750 30270 20802
rect 30322 20750 30324 20802
rect 29932 20692 29988 20702
rect 29932 20242 29988 20636
rect 30044 20580 30100 20590
rect 30044 20486 30100 20524
rect 29932 20190 29934 20242
rect 29986 20190 29988 20242
rect 29932 20178 29988 20190
rect 29260 17602 29316 17612
rect 29372 18450 29428 18462
rect 29372 18398 29374 18450
rect 29426 18398 29428 18450
rect 29148 16996 29204 17006
rect 29372 16996 29428 18398
rect 29484 17780 29540 20076
rect 29820 20066 29876 20076
rect 29708 20020 29764 20030
rect 29708 19926 29764 19964
rect 30156 20018 30212 20030
rect 30156 19966 30158 20018
rect 30210 19966 30212 20018
rect 30156 19908 30212 19966
rect 30156 19842 30212 19852
rect 29596 19122 29652 19134
rect 29596 19070 29598 19122
rect 29650 19070 29652 19122
rect 29596 18452 29652 19070
rect 29932 19124 29988 19134
rect 29932 19030 29988 19068
rect 30268 19124 30324 20750
rect 30380 20580 30436 21756
rect 30380 20514 30436 20524
rect 30492 20132 30548 24332
rect 30604 23604 30660 26852
rect 30604 23538 30660 23548
rect 30716 22484 30772 28364
rect 30828 27076 30884 29262
rect 30940 27300 30996 29708
rect 31052 29428 31108 29438
rect 31164 29428 31220 30046
rect 31052 29426 31220 29428
rect 31052 29374 31054 29426
rect 31106 29374 31220 29426
rect 31052 29372 31220 29374
rect 31276 30884 31332 30894
rect 31052 28644 31108 29372
rect 31276 29316 31332 30828
rect 31500 30436 31556 30446
rect 31500 30342 31556 30380
rect 31500 30210 31556 30222
rect 31500 30158 31502 30210
rect 31554 30158 31556 30210
rect 31388 30100 31444 30110
rect 31500 30100 31556 30158
rect 31388 30098 31556 30100
rect 31388 30046 31390 30098
rect 31442 30046 31556 30098
rect 31388 30044 31556 30046
rect 31388 30034 31444 30044
rect 31052 28578 31108 28588
rect 31164 29260 31332 29316
rect 31052 28084 31108 28094
rect 31052 27990 31108 28028
rect 31164 28082 31220 29260
rect 31276 28868 31332 28878
rect 31276 28774 31332 28812
rect 31276 28532 31332 28542
rect 31276 28308 31332 28476
rect 31388 28532 31444 28542
rect 31388 28530 31556 28532
rect 31388 28478 31390 28530
rect 31442 28478 31556 28530
rect 31388 28476 31556 28478
rect 31388 28466 31444 28476
rect 31500 28420 31556 28476
rect 31276 28252 31444 28308
rect 31164 28030 31166 28082
rect 31218 28030 31220 28082
rect 31164 28018 31220 28030
rect 30940 27234 30996 27244
rect 31276 27858 31332 27870
rect 31276 27806 31278 27858
rect 31330 27806 31332 27858
rect 30940 27076 30996 27086
rect 30828 27074 30996 27076
rect 30828 27022 30942 27074
rect 30994 27022 30996 27074
rect 30828 27020 30996 27022
rect 30828 26964 30884 27020
rect 30940 27010 30996 27020
rect 31164 27074 31220 27086
rect 31164 27022 31166 27074
rect 31218 27022 31220 27074
rect 31164 26908 31220 27022
rect 30828 24836 30884 26908
rect 31052 26852 31220 26908
rect 31276 27076 31332 27806
rect 31276 26908 31332 27020
rect 31388 27074 31444 28252
rect 31500 27412 31556 28364
rect 31500 27346 31556 27356
rect 31500 27188 31556 27198
rect 31612 27188 31668 32732
rect 31836 32674 31892 34300
rect 31836 32622 31838 32674
rect 31890 32622 31892 32674
rect 31836 30324 31892 32622
rect 31948 33346 32004 33358
rect 31948 33294 31950 33346
rect 32002 33294 32004 33346
rect 31948 31892 32004 33294
rect 31948 31826 32004 31836
rect 31948 31220 32004 31230
rect 31948 31126 32004 31164
rect 31724 30268 31892 30324
rect 31724 29540 31780 30268
rect 31836 30098 31892 30110
rect 31836 30046 31838 30098
rect 31890 30046 31892 30098
rect 31836 29988 31892 30046
rect 31836 29922 31892 29932
rect 31724 29484 31892 29540
rect 31724 29314 31780 29326
rect 31724 29262 31726 29314
rect 31778 29262 31780 29314
rect 31724 29204 31780 29262
rect 31724 29138 31780 29148
rect 31836 28644 31892 29484
rect 31724 28588 31892 28644
rect 31724 28084 31780 28588
rect 32060 28308 32116 36876
rect 32172 36484 32228 36494
rect 32172 28756 32228 36428
rect 32284 36482 32340 36494
rect 32284 36430 32286 36482
rect 32338 36430 32340 36482
rect 32284 35140 32340 36430
rect 32732 36484 32788 36494
rect 32732 36390 32788 36428
rect 32396 36036 32452 36046
rect 32396 35922 32452 35980
rect 32396 35870 32398 35922
rect 32450 35870 32452 35922
rect 32396 35858 32452 35870
rect 32732 35588 32788 35598
rect 32844 35588 32900 38612
rect 32956 37492 33012 37502
rect 32956 37398 33012 37436
rect 32732 35586 32900 35588
rect 32732 35534 32734 35586
rect 32786 35534 32900 35586
rect 32732 35532 32900 35534
rect 33068 35924 33124 43484
rect 33404 43316 33460 43326
rect 33180 36596 33236 36606
rect 33180 36502 33236 36540
rect 32732 35476 32788 35532
rect 32732 35410 32788 35420
rect 32396 35140 32452 35150
rect 32284 35138 32452 35140
rect 32284 35086 32398 35138
rect 32450 35086 32452 35138
rect 32284 35084 32452 35086
rect 32284 34356 32340 35084
rect 32396 35074 32452 35084
rect 32956 35028 33012 35038
rect 33068 35028 33124 35868
rect 32508 35026 33124 35028
rect 32508 34974 32958 35026
rect 33010 34974 33124 35026
rect 32508 34972 33124 34974
rect 33180 36372 33236 36382
rect 32508 34914 32564 34972
rect 32956 34962 33012 34972
rect 32508 34862 32510 34914
rect 32562 34862 32564 34914
rect 32508 34850 32564 34862
rect 32396 34692 32452 34702
rect 32396 34598 32452 34636
rect 32284 34290 32340 34300
rect 32508 33348 32564 33358
rect 32508 33254 32564 33292
rect 32396 33124 32452 33134
rect 32396 33030 32452 33068
rect 32620 33124 32676 33134
rect 32620 33122 32788 33124
rect 32620 33070 32622 33122
rect 32674 33070 32788 33122
rect 32620 33068 32788 33070
rect 32620 33058 32676 33068
rect 32732 32452 32788 33068
rect 32844 32452 32900 32462
rect 32732 32396 32844 32452
rect 32844 32358 32900 32396
rect 32956 32004 33012 32014
rect 32732 31220 32788 31230
rect 32284 30212 32340 30222
rect 32284 30118 32340 30156
rect 32508 29538 32564 29550
rect 32508 29486 32510 29538
rect 32562 29486 32564 29538
rect 32508 28980 32564 29486
rect 32172 28690 32228 28700
rect 32284 28868 32340 28878
rect 32284 28754 32340 28812
rect 32284 28702 32286 28754
rect 32338 28702 32340 28754
rect 32284 28690 32340 28702
rect 32172 28532 32228 28542
rect 32172 28438 32228 28476
rect 32396 28530 32452 28542
rect 32396 28478 32398 28530
rect 32450 28478 32452 28530
rect 32396 28308 32452 28478
rect 32060 28252 32452 28308
rect 31724 27636 31780 28028
rect 32396 28084 32452 28252
rect 32396 28018 32452 28028
rect 31724 27580 31892 27636
rect 31500 27186 31668 27188
rect 31500 27134 31502 27186
rect 31554 27134 31668 27186
rect 31500 27132 31668 27134
rect 31724 27412 31780 27422
rect 31500 27122 31556 27132
rect 31388 27022 31390 27074
rect 31442 27022 31444 27074
rect 31388 27010 31444 27022
rect 31276 26852 31444 26908
rect 31052 25620 31108 26852
rect 31276 26290 31332 26302
rect 31276 26238 31278 26290
rect 31330 26238 31332 26290
rect 31276 25956 31332 26238
rect 31276 25890 31332 25900
rect 31388 25732 31444 26852
rect 31612 26850 31668 26862
rect 31612 26798 31614 26850
rect 31666 26798 31668 26850
rect 30940 25396 30996 25406
rect 31052 25396 31108 25564
rect 31276 25676 31444 25732
rect 31500 26292 31556 26302
rect 31276 25506 31332 25676
rect 31276 25454 31278 25506
rect 31330 25454 31332 25506
rect 31276 25442 31332 25454
rect 30940 25394 31108 25396
rect 30940 25342 30942 25394
rect 30994 25342 31108 25394
rect 30940 25340 31108 25342
rect 31388 25396 31444 25406
rect 31500 25396 31556 26236
rect 31612 25956 31668 26798
rect 31724 26402 31780 27356
rect 31724 26350 31726 26402
rect 31778 26350 31780 26402
rect 31724 26338 31780 26350
rect 31724 26180 31780 26190
rect 31724 26086 31780 26124
rect 31612 25890 31668 25900
rect 31836 25508 31892 27580
rect 32284 27188 32340 27198
rect 31388 25394 31556 25396
rect 31388 25342 31390 25394
rect 31442 25342 31556 25394
rect 31388 25340 31556 25342
rect 31612 25452 31892 25508
rect 31948 27186 32340 27188
rect 31948 27134 32286 27186
rect 32338 27134 32340 27186
rect 31948 27132 32340 27134
rect 31948 26180 32004 27132
rect 32284 27122 32340 27132
rect 32172 26964 32228 26974
rect 32172 26628 32228 26908
rect 32396 26962 32452 26974
rect 32396 26910 32398 26962
rect 32450 26910 32452 26962
rect 32396 26852 32452 26910
rect 32396 26786 32452 26796
rect 32172 26572 32452 26628
rect 32172 26404 32228 26414
rect 32172 26310 32228 26348
rect 32060 26292 32116 26302
rect 32060 26198 32116 26236
rect 31948 25506 32004 26124
rect 32284 25956 32340 25966
rect 32060 25620 32116 25630
rect 32060 25526 32116 25564
rect 31948 25454 31950 25506
rect 32002 25454 32004 25506
rect 30940 25330 30996 25340
rect 31388 25330 31444 25340
rect 31164 25282 31220 25294
rect 31164 25230 31166 25282
rect 31218 25230 31220 25282
rect 30828 24780 30996 24836
rect 30828 24610 30884 24622
rect 30828 24558 30830 24610
rect 30882 24558 30884 24610
rect 30828 24276 30884 24558
rect 30828 24210 30884 24220
rect 30940 23938 30996 24780
rect 31164 24612 31220 25230
rect 31164 24546 31220 24556
rect 31276 25172 31332 25182
rect 31612 25172 31668 25452
rect 31948 25442 32004 25454
rect 32284 25396 32340 25900
rect 32284 25302 32340 25340
rect 31164 24164 31220 24174
rect 31164 24070 31220 24108
rect 30940 23886 30942 23938
rect 30994 23886 30996 23938
rect 30940 23156 30996 23886
rect 31164 23156 31220 23166
rect 30940 23154 31220 23156
rect 30940 23102 31166 23154
rect 31218 23102 31220 23154
rect 30940 23100 31220 23102
rect 31164 23090 31220 23100
rect 30716 22418 30772 22428
rect 30604 22260 30660 22270
rect 30604 22166 30660 22204
rect 30828 21812 30884 21822
rect 30828 21718 30884 21756
rect 31276 21812 31332 25116
rect 31388 25116 31668 25172
rect 31724 25284 31780 25294
rect 31388 23716 31444 25116
rect 31612 24612 31668 24622
rect 31612 24518 31668 24556
rect 31724 24388 31780 25228
rect 32172 24612 32228 24622
rect 31612 24332 31780 24388
rect 32060 24500 32116 24510
rect 31500 23940 31556 23950
rect 31500 23846 31556 23884
rect 31388 23660 31556 23716
rect 31388 22484 31444 22494
rect 31388 22390 31444 22428
rect 31276 21746 31332 21756
rect 31276 21588 31332 21598
rect 31276 21494 31332 21532
rect 30716 21364 30772 21374
rect 30716 20132 30772 21308
rect 30828 20804 30884 20814
rect 30828 20710 30884 20748
rect 31500 20692 31556 23660
rect 31500 20626 31556 20636
rect 30492 20076 30660 20132
rect 30380 20020 30436 20030
rect 30380 20018 30548 20020
rect 30380 19966 30382 20018
rect 30434 19966 30548 20018
rect 30380 19964 30548 19966
rect 30380 19954 30436 19964
rect 30492 19794 30548 19964
rect 30492 19742 30494 19794
rect 30546 19742 30548 19794
rect 30492 19730 30548 19742
rect 30268 19058 30324 19068
rect 30604 19122 30660 20076
rect 30716 20076 31220 20132
rect 30716 19234 30772 20076
rect 30716 19182 30718 19234
rect 30770 19182 30772 19234
rect 30716 19170 30772 19182
rect 30828 19906 30884 19918
rect 30828 19854 30830 19906
rect 30882 19854 30884 19906
rect 30828 19794 30884 19854
rect 30828 19742 30830 19794
rect 30882 19742 30884 19794
rect 30604 19070 30606 19122
rect 30658 19070 30660 19122
rect 30380 19010 30436 19022
rect 30380 18958 30382 19010
rect 30434 18958 30436 19010
rect 30268 18900 30324 18910
rect 29708 18788 29764 18798
rect 29708 18674 29764 18732
rect 29708 18622 29710 18674
rect 29762 18622 29764 18674
rect 29708 18610 29764 18622
rect 30156 18788 30212 18798
rect 30156 18674 30212 18732
rect 30156 18622 30158 18674
rect 30210 18622 30212 18674
rect 30156 18610 30212 18622
rect 29596 18386 29652 18396
rect 29484 17714 29540 17724
rect 29820 17668 29876 17678
rect 29876 17612 29988 17668
rect 29820 17574 29876 17612
rect 29484 17444 29540 17454
rect 29484 17350 29540 17388
rect 29708 17442 29764 17454
rect 29708 17390 29710 17442
rect 29762 17390 29764 17442
rect 29148 16994 29428 16996
rect 29148 16942 29150 16994
rect 29202 16942 29428 16994
rect 29148 16940 29428 16942
rect 29148 16884 29204 16940
rect 29148 16818 29204 16828
rect 29484 16884 29540 16894
rect 29708 16884 29764 17390
rect 29932 17106 29988 17612
rect 29932 17054 29934 17106
rect 29986 17054 29988 17106
rect 29932 17042 29988 17054
rect 29484 16882 29764 16884
rect 29484 16830 29486 16882
rect 29538 16830 29764 16882
rect 29484 16828 29764 16830
rect 29484 15988 29540 16828
rect 29932 16100 29988 16110
rect 29932 16006 29988 16044
rect 29596 15988 29652 15998
rect 29484 15986 29652 15988
rect 29484 15934 29598 15986
rect 29650 15934 29652 15986
rect 29484 15932 29652 15934
rect 29484 15764 29540 15932
rect 29596 15922 29652 15932
rect 29484 15698 29540 15708
rect 29596 15652 29652 15662
rect 29260 15540 29316 15550
rect 29260 15148 29316 15484
rect 29036 11330 29092 11340
rect 29148 15092 29316 15148
rect 29372 15092 29428 15102
rect 28588 10770 28644 10780
rect 28364 9874 28420 9884
rect 28476 10722 28532 10734
rect 28476 10670 28478 10722
rect 28530 10670 28532 10722
rect 28476 10500 28532 10670
rect 28364 9268 28420 9278
rect 28364 9174 28420 9212
rect 28252 8766 28254 8818
rect 28306 8766 28308 8818
rect 28252 8754 28308 8766
rect 28476 6020 28532 10444
rect 28700 10612 28756 10622
rect 28700 9602 28756 10556
rect 28700 9550 28702 9602
rect 28754 9550 28756 9602
rect 28700 9492 28756 9550
rect 28700 9426 28756 9436
rect 28476 5954 28532 5964
rect 28812 5236 28868 5246
rect 28812 5142 28868 5180
rect 28364 5012 28420 5022
rect 28364 4918 28420 4956
rect 28140 4498 28196 4508
rect 28028 3938 28084 3948
rect 27580 1362 27636 1372
rect 28252 3444 28308 3454
rect 28252 800 28308 3388
rect 29148 1316 29204 15092
rect 29260 10500 29316 10510
rect 29260 10406 29316 10444
rect 29372 8260 29428 15036
rect 29596 14642 29652 15596
rect 29932 15652 29988 15662
rect 29932 15538 29988 15596
rect 29932 15486 29934 15538
rect 29986 15486 29988 15538
rect 29932 15474 29988 15486
rect 30156 15314 30212 15326
rect 30156 15262 30158 15314
rect 30210 15262 30212 15314
rect 30044 15202 30100 15214
rect 30044 15150 30046 15202
rect 30098 15150 30100 15202
rect 30044 15092 30100 15150
rect 30044 15026 30100 15036
rect 30156 15204 30212 15262
rect 29596 14590 29598 14642
rect 29650 14590 29652 14642
rect 29596 14578 29652 14590
rect 29708 14644 29764 14654
rect 29484 14532 29540 14542
rect 29484 13746 29540 14476
rect 29708 14420 29764 14588
rect 30044 14532 30100 14542
rect 30044 14438 30100 14476
rect 29484 13694 29486 13746
rect 29538 13694 29540 13746
rect 29484 13682 29540 13694
rect 29596 14364 29764 14420
rect 29596 13074 29652 14364
rect 30156 13970 30212 15148
rect 30268 15148 30324 18844
rect 30380 17220 30436 18958
rect 30604 18788 30660 19070
rect 30604 18722 30660 18732
rect 30828 18228 30884 19742
rect 31164 19348 31220 20076
rect 30492 18226 30884 18228
rect 30492 18174 30830 18226
rect 30882 18174 30884 18226
rect 30492 18172 30884 18174
rect 30492 17444 30548 18172
rect 30828 18162 30884 18172
rect 31052 19346 31220 19348
rect 31052 19294 31166 19346
rect 31218 19294 31220 19346
rect 31052 19292 31220 19294
rect 31052 17556 31108 19292
rect 31164 19282 31220 19292
rect 31276 19908 31332 19918
rect 31276 18900 31332 19852
rect 31276 18834 31332 18844
rect 31276 18676 31332 18686
rect 31276 18582 31332 18620
rect 31500 18676 31556 18686
rect 31500 18582 31556 18620
rect 31164 18564 31220 18574
rect 31164 18450 31220 18508
rect 31164 18398 31166 18450
rect 31218 18398 31220 18450
rect 31164 17890 31220 18398
rect 31164 17838 31166 17890
rect 31218 17838 31220 17890
rect 31164 17826 31220 17838
rect 31388 18338 31444 18350
rect 31388 18286 31390 18338
rect 31442 18286 31444 18338
rect 31164 17556 31220 17566
rect 30492 17350 30548 17388
rect 30716 17554 31220 17556
rect 30716 17502 31166 17554
rect 31218 17502 31220 17554
rect 30716 17500 31220 17502
rect 30380 17154 30436 17164
rect 30716 17108 30772 17500
rect 31164 17490 31220 17500
rect 31276 17554 31332 17566
rect 31276 17502 31278 17554
rect 31330 17502 31332 17554
rect 30604 17106 30772 17108
rect 30604 17054 30718 17106
rect 30770 17054 30772 17106
rect 30604 17052 30772 17054
rect 30380 16100 30436 16110
rect 30380 16006 30436 16044
rect 30604 15540 30660 17052
rect 30716 17042 30772 17052
rect 31052 17332 31108 17342
rect 30828 16324 30884 16334
rect 30828 16210 30884 16268
rect 30828 16158 30830 16210
rect 30882 16158 30884 16210
rect 30828 16146 30884 16158
rect 30380 15316 30436 15354
rect 30380 15250 30436 15260
rect 30604 15314 30660 15484
rect 30604 15262 30606 15314
rect 30658 15262 30660 15314
rect 30604 15250 30660 15262
rect 30828 15876 30884 15886
rect 30828 15316 30884 15820
rect 30716 15204 30772 15214
rect 30268 15092 30548 15148
rect 30268 14644 30324 14654
rect 30268 14550 30324 14588
rect 30492 14306 30548 15092
rect 30492 14254 30494 14306
rect 30546 14254 30548 14306
rect 30492 14084 30548 14254
rect 30604 14308 30660 14318
rect 30604 14214 30660 14252
rect 30716 14306 30772 15148
rect 30828 15090 30884 15260
rect 30828 15038 30830 15090
rect 30882 15038 30884 15090
rect 30828 14532 30884 15038
rect 30828 14466 30884 14476
rect 30716 14254 30718 14306
rect 30770 14254 30772 14306
rect 30492 14018 30548 14028
rect 30156 13918 30158 13970
rect 30210 13918 30212 13970
rect 30156 13906 30212 13918
rect 30716 13972 30772 14254
rect 30940 13972 30996 13982
rect 30716 13916 30940 13972
rect 30940 13878 30996 13916
rect 30380 13748 30436 13758
rect 29932 13636 29988 13646
rect 29932 13542 29988 13580
rect 30268 13634 30324 13646
rect 30268 13582 30270 13634
rect 30322 13582 30324 13634
rect 29596 13022 29598 13074
rect 29650 13022 29652 13074
rect 29596 13010 29652 13022
rect 29708 13522 29764 13534
rect 29708 13470 29710 13522
rect 29762 13470 29764 13522
rect 29708 12628 29764 13470
rect 29708 12562 29764 12572
rect 29820 13076 29876 13086
rect 29820 12852 29876 13020
rect 29820 12402 29876 12796
rect 29932 12738 29988 12750
rect 29932 12686 29934 12738
rect 29986 12686 29988 12738
rect 29932 12628 29988 12686
rect 29932 12562 29988 12572
rect 29820 12350 29822 12402
rect 29874 12350 29876 12402
rect 29820 12338 29876 12350
rect 30268 12292 30324 13582
rect 30380 13074 30436 13692
rect 30380 13022 30382 13074
rect 30434 13022 30436 13074
rect 30380 13010 30436 13022
rect 30492 13076 30548 13086
rect 30268 12236 30436 12292
rect 29596 12178 29652 12190
rect 29596 12126 29598 12178
rect 29650 12126 29652 12178
rect 29596 11844 29652 12126
rect 29596 11778 29652 11788
rect 30268 12066 30324 12078
rect 30268 12014 30270 12066
rect 30322 12014 30324 12066
rect 30268 11844 30324 12014
rect 30268 11778 30324 11788
rect 29596 11284 29652 11294
rect 29596 11190 29652 11228
rect 29932 11282 29988 11294
rect 29932 11230 29934 11282
rect 29986 11230 29988 11282
rect 29820 10836 29876 10846
rect 29820 10742 29876 10780
rect 29932 10500 29988 11230
rect 30156 10724 30212 10734
rect 30156 10630 30212 10668
rect 29932 10434 29988 10444
rect 29484 9940 29540 9950
rect 29484 9846 29540 9884
rect 29372 8194 29428 8204
rect 30380 6132 30436 12236
rect 30492 11506 30548 13020
rect 30828 13076 30884 13086
rect 30828 12982 30884 13020
rect 30492 11454 30494 11506
rect 30546 11454 30548 11506
rect 30492 11442 30548 11454
rect 30716 12180 30772 12190
rect 30716 12066 30772 12124
rect 30716 12014 30718 12066
rect 30770 12014 30772 12066
rect 30716 10388 30772 12014
rect 30828 11170 30884 11182
rect 30828 11118 30830 11170
rect 30882 11118 30884 11170
rect 30828 11060 30884 11118
rect 30828 10994 30884 11004
rect 30716 10322 30772 10332
rect 30380 6066 30436 6076
rect 31052 5236 31108 17276
rect 31276 17108 31332 17502
rect 31276 17042 31332 17052
rect 31276 15876 31332 15886
rect 31164 15874 31332 15876
rect 31164 15822 31278 15874
rect 31330 15822 31332 15874
rect 31164 15820 31332 15822
rect 31164 14868 31220 15820
rect 31276 15810 31332 15820
rect 31164 14802 31220 14812
rect 31276 15204 31332 15280
rect 31276 14642 31332 15148
rect 31388 15148 31444 18286
rect 31612 17332 31668 24332
rect 31836 24052 31892 24062
rect 31836 23266 31892 23996
rect 31836 23214 31838 23266
rect 31890 23214 31892 23266
rect 31836 23202 31892 23214
rect 31724 23154 31780 23166
rect 31724 23102 31726 23154
rect 31778 23102 31780 23154
rect 31724 22596 31780 23102
rect 32060 22932 32116 24444
rect 32060 22866 32116 22876
rect 31724 22540 32004 22596
rect 31948 22482 32004 22540
rect 31948 22430 31950 22482
rect 32002 22430 32004 22482
rect 31948 22418 32004 22430
rect 31836 22372 31892 22382
rect 31836 22278 31892 22316
rect 32060 22146 32116 22158
rect 32060 22094 32062 22146
rect 32114 22094 32116 22146
rect 32060 22036 32116 22094
rect 32060 21970 32116 21980
rect 31948 21476 32004 21486
rect 32172 21476 32228 24556
rect 32284 23940 32340 23950
rect 32284 23378 32340 23884
rect 32396 23492 32452 26572
rect 32508 26404 32564 28924
rect 32620 28084 32676 28094
rect 32620 27990 32676 28028
rect 32508 25284 32564 26348
rect 32620 26962 32676 26974
rect 32620 26910 32622 26962
rect 32674 26910 32676 26962
rect 32620 26180 32676 26910
rect 32732 26964 32788 31164
rect 32844 30436 32900 30446
rect 32844 29650 32900 30380
rect 32844 29598 32846 29650
rect 32898 29598 32900 29650
rect 32844 29586 32900 29598
rect 32956 26908 33012 31948
rect 33180 31220 33236 36316
rect 33292 33348 33348 33358
rect 33292 33254 33348 33292
rect 33180 31154 33236 31164
rect 33180 29988 33236 29998
rect 33180 29894 33236 29932
rect 33180 29092 33236 29102
rect 33068 28868 33124 28878
rect 33068 28754 33124 28812
rect 33068 28702 33070 28754
rect 33122 28702 33124 28754
rect 33068 28690 33124 28702
rect 33180 28532 33236 29036
rect 32732 26898 32788 26908
rect 32620 26114 32676 26124
rect 32844 26852 33012 26908
rect 33068 28476 33236 28532
rect 32732 25284 32788 25294
rect 32508 25282 32788 25284
rect 32508 25230 32734 25282
rect 32786 25230 32788 25282
rect 32508 25228 32788 25230
rect 32508 25060 32564 25070
rect 32508 24946 32564 25004
rect 32508 24894 32510 24946
rect 32562 24894 32564 24946
rect 32508 24882 32564 24894
rect 32732 23828 32788 25228
rect 32508 23716 32564 23726
rect 32732 23716 32788 23772
rect 32508 23714 32788 23716
rect 32508 23662 32510 23714
rect 32562 23662 32788 23714
rect 32508 23660 32788 23662
rect 32508 23650 32564 23660
rect 32396 23436 32564 23492
rect 32284 23326 32286 23378
rect 32338 23326 32340 23378
rect 32284 23314 32340 23326
rect 32396 23268 32452 23278
rect 32396 23174 32452 23212
rect 32284 23044 32340 23054
rect 32284 22370 32340 22988
rect 32508 22484 32564 23436
rect 32620 23380 32676 23390
rect 32620 23286 32676 23324
rect 32284 22318 32286 22370
rect 32338 22318 32340 22370
rect 32284 22306 32340 22318
rect 32396 22428 32564 22484
rect 31948 21474 32228 21476
rect 31948 21422 31950 21474
rect 32002 21422 32228 21474
rect 31948 21420 32228 21422
rect 31948 21026 32004 21420
rect 31948 20974 31950 21026
rect 32002 20974 32004 21026
rect 31948 20962 32004 20974
rect 32284 20916 32340 20926
rect 32284 20822 32340 20860
rect 31836 20578 31892 20590
rect 31836 20526 31838 20578
rect 31890 20526 31892 20578
rect 31836 20244 31892 20526
rect 31836 20178 31892 20188
rect 31948 20580 32004 20590
rect 31724 19906 31780 19918
rect 31724 19854 31726 19906
rect 31778 19854 31780 19906
rect 31724 19684 31780 19854
rect 31724 19618 31780 19628
rect 31836 19012 31892 19022
rect 31948 19012 32004 20524
rect 31836 19010 32004 19012
rect 31836 18958 31838 19010
rect 31890 18958 32004 19010
rect 31836 18956 32004 18958
rect 31836 18788 31892 18956
rect 31836 18722 31892 18732
rect 32172 18564 32228 18574
rect 32172 18470 32228 18508
rect 32284 18340 32340 18350
rect 32172 18338 32340 18340
rect 32172 18286 32286 18338
rect 32338 18286 32340 18338
rect 32172 18284 32340 18286
rect 32060 17556 32116 17566
rect 32060 17462 32116 17500
rect 31612 17266 31668 17276
rect 32172 17332 32228 18284
rect 32284 18274 32340 18284
rect 32172 17266 32228 17276
rect 32284 17554 32340 17566
rect 32284 17502 32286 17554
rect 32338 17502 32340 17554
rect 31724 17220 31780 17230
rect 31724 17106 31780 17164
rect 32284 17220 32340 17502
rect 32284 17154 32340 17164
rect 31724 17054 31726 17106
rect 31778 17054 31780 17106
rect 31724 17042 31780 17054
rect 32172 17108 32228 17118
rect 32172 17014 32228 17052
rect 31948 16996 32004 17006
rect 31948 15986 32004 16940
rect 32060 16884 32116 16894
rect 32060 16098 32116 16828
rect 32060 16046 32062 16098
rect 32114 16046 32116 16098
rect 32060 16034 32116 16046
rect 31948 15934 31950 15986
rect 32002 15934 32004 15986
rect 31948 15922 32004 15934
rect 31724 15876 31780 15886
rect 31724 15782 31780 15820
rect 31724 15540 31780 15550
rect 32396 15540 32452 22428
rect 32508 22258 32564 22270
rect 32508 22206 32510 22258
rect 32562 22206 32564 22258
rect 32508 21700 32564 22206
rect 32732 22036 32788 23660
rect 32844 23268 32900 26852
rect 32956 24948 33012 24958
rect 32956 24854 33012 24892
rect 33068 24276 33124 28476
rect 33404 26908 33460 43260
rect 33852 42868 33908 46732
rect 33964 46786 34020 46844
rect 33964 46734 33966 46786
rect 34018 46734 34020 46786
rect 33964 46722 34020 46734
rect 34412 46676 34468 46686
rect 34412 46582 34468 46620
rect 34524 45444 34580 45454
rect 34188 45106 34244 45118
rect 34188 45054 34190 45106
rect 34242 45054 34244 45106
rect 34188 44548 34244 45054
rect 34188 44482 34244 44492
rect 34524 43762 34580 45388
rect 34524 43710 34526 43762
rect 34578 43710 34580 43762
rect 34524 43652 34580 43710
rect 34524 43586 34580 43596
rect 34748 43204 34804 47180
rect 34860 46898 34916 47292
rect 34860 46846 34862 46898
rect 34914 46846 34916 46898
rect 34860 46788 34916 46846
rect 34860 46722 34916 46732
rect 34972 45220 35028 48412
rect 35084 47682 35140 48524
rect 35308 48020 35364 48750
rect 35868 48354 35924 48860
rect 35868 48302 35870 48354
rect 35922 48302 35924 48354
rect 35868 48290 35924 48302
rect 35980 48802 36036 48814
rect 35980 48750 35982 48802
rect 36034 48750 36036 48802
rect 35756 48244 35812 48254
rect 35756 48150 35812 48188
rect 35532 48020 35588 48030
rect 35308 47964 35532 48020
rect 35532 47926 35588 47964
rect 35980 48020 36036 48750
rect 35980 47954 36036 47964
rect 36092 48018 36148 48030
rect 36316 48020 36372 50316
rect 36428 49810 36484 51324
rect 36540 50596 36596 51548
rect 37436 51380 37492 51390
rect 37436 51286 37492 51324
rect 37548 51266 37604 51548
rect 37548 51214 37550 51266
rect 37602 51214 37604 51266
rect 37548 51202 37604 51214
rect 37436 50820 37492 50830
rect 36652 50818 37492 50820
rect 36652 50766 37438 50818
rect 37490 50766 37492 50818
rect 36652 50764 37492 50766
rect 36652 50596 36708 50764
rect 37436 50706 37492 50764
rect 37884 50818 37940 51886
rect 37884 50766 37886 50818
rect 37938 50766 37940 50818
rect 37884 50754 37940 50766
rect 37996 52276 38052 52286
rect 37436 50654 37438 50706
rect 37490 50654 37492 50706
rect 37436 50642 37492 50654
rect 36540 50594 36708 50596
rect 36540 50542 36542 50594
rect 36594 50542 36708 50594
rect 36540 50540 36708 50542
rect 36540 50530 36596 50540
rect 36428 49758 36430 49810
rect 36482 49758 36484 49810
rect 36428 49746 36484 49758
rect 36092 47966 36094 48018
rect 36146 47966 36148 48018
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 36092 47796 36148 47966
rect 36092 47730 36148 47740
rect 36204 48018 36372 48020
rect 36204 47966 36318 48018
rect 36370 47966 36372 48018
rect 36204 47964 36372 47966
rect 35084 47630 35086 47682
rect 35138 47630 35140 47682
rect 35084 47572 35140 47630
rect 35196 47572 35252 47582
rect 35084 47570 35252 47572
rect 35084 47518 35198 47570
rect 35250 47518 35252 47570
rect 35084 47516 35252 47518
rect 35196 47506 35252 47516
rect 34636 43148 34804 43204
rect 34860 45164 35028 45220
rect 35084 47348 35140 47358
rect 33964 42868 34020 42878
rect 33852 42866 34020 42868
rect 33852 42814 33966 42866
rect 34018 42814 34020 42866
rect 33852 42812 34020 42814
rect 33852 42756 33908 42812
rect 33964 42802 34020 42812
rect 33852 42690 33908 42700
rect 33516 42532 33572 42542
rect 33516 42438 33572 42476
rect 34076 42084 34132 42094
rect 34076 41990 34132 42028
rect 33628 41972 33684 41982
rect 33628 41878 33684 41916
rect 34300 41748 34356 41758
rect 34188 41188 34244 41198
rect 33964 41186 34244 41188
rect 33964 41134 34190 41186
rect 34242 41134 34244 41186
rect 33964 41132 34244 41134
rect 33852 41076 33908 41086
rect 33852 40982 33908 41020
rect 33740 40514 33796 40526
rect 33740 40462 33742 40514
rect 33794 40462 33796 40514
rect 33516 40402 33572 40414
rect 33516 40350 33518 40402
rect 33570 40350 33572 40402
rect 33516 39730 33572 40350
rect 33516 39678 33518 39730
rect 33570 39678 33572 39730
rect 33516 39666 33572 39678
rect 33628 40404 33684 40414
rect 33628 39618 33684 40348
rect 33628 39566 33630 39618
rect 33682 39566 33684 39618
rect 33628 39554 33684 39566
rect 33628 39060 33684 39070
rect 33628 38966 33684 39004
rect 33740 38724 33796 40462
rect 33852 40516 33908 40526
rect 33852 40422 33908 40460
rect 33964 39844 34020 41132
rect 34188 41122 34244 41132
rect 34300 41186 34356 41692
rect 34300 41134 34302 41186
rect 34354 41134 34356 41186
rect 34300 41122 34356 41134
rect 34076 40964 34132 40974
rect 34076 40870 34132 40908
rect 33740 38658 33796 38668
rect 33852 39788 34020 39844
rect 34076 40516 34132 40526
rect 33740 38164 33796 38174
rect 33516 38050 33572 38062
rect 33516 37998 33518 38050
rect 33570 37998 33572 38050
rect 33516 37492 33572 37998
rect 33516 37426 33572 37436
rect 33628 37268 33684 37278
rect 33628 37174 33684 37212
rect 33740 37266 33796 38108
rect 33740 37214 33742 37266
rect 33794 37214 33796 37266
rect 33740 37202 33796 37214
rect 33852 37826 33908 39788
rect 34076 38946 34132 40460
rect 34076 38894 34078 38946
rect 34130 38894 34132 38946
rect 34076 38882 34132 38894
rect 34300 40404 34356 40414
rect 34300 38946 34356 40348
rect 34300 38894 34302 38946
rect 34354 38894 34356 38946
rect 34300 38882 34356 38894
rect 34188 38834 34244 38846
rect 34188 38782 34190 38834
rect 34242 38782 34244 38834
rect 34188 38724 34244 38782
rect 34188 38658 34244 38668
rect 33964 38612 34020 38622
rect 33964 38162 34020 38556
rect 33964 38110 33966 38162
rect 34018 38110 34020 38162
rect 33964 38098 34020 38110
rect 34076 38164 34132 38174
rect 34076 38050 34132 38108
rect 34076 37998 34078 38050
rect 34130 37998 34132 38050
rect 34076 37986 34132 37998
rect 34300 38052 34356 38062
rect 33852 37774 33854 37826
rect 33906 37774 33908 37826
rect 33852 37268 33908 37774
rect 34076 37268 34132 37278
rect 33852 37266 34132 37268
rect 33852 37214 34078 37266
rect 34130 37214 34132 37266
rect 33852 37212 34132 37214
rect 34076 37202 34132 37212
rect 33628 36484 33684 36494
rect 33628 36390 33684 36428
rect 34188 36036 34244 36046
rect 33628 34802 33684 34814
rect 33628 34750 33630 34802
rect 33682 34750 33684 34802
rect 33516 33348 33572 33358
rect 33516 33254 33572 33292
rect 33628 33124 33684 34750
rect 33740 34692 33796 34702
rect 33740 34598 33796 34636
rect 33964 34690 34020 34702
rect 33964 34638 33966 34690
rect 34018 34638 34020 34690
rect 33964 34130 34020 34638
rect 33964 34078 33966 34130
rect 34018 34078 34020 34130
rect 33964 34066 34020 34078
rect 33628 33058 33684 33068
rect 33740 34018 33796 34030
rect 33740 33966 33742 34018
rect 33794 33966 33796 34018
rect 33740 33572 33796 33966
rect 33740 32452 33796 33516
rect 34188 33458 34244 35980
rect 34188 33406 34190 33458
rect 34242 33406 34244 33458
rect 34188 33394 34244 33406
rect 33740 32386 33796 32396
rect 33852 33124 33908 33134
rect 33740 31780 33796 31790
rect 33628 31108 33684 31118
rect 33628 31014 33684 31052
rect 33516 30436 33572 30446
rect 33516 29650 33572 30380
rect 33740 29876 33796 31724
rect 33852 30994 33908 33068
rect 34188 32452 34244 32462
rect 33964 31890 34020 31902
rect 33964 31838 33966 31890
rect 34018 31838 34020 31890
rect 33964 31106 34020 31838
rect 33964 31054 33966 31106
rect 34018 31054 34020 31106
rect 33964 31042 34020 31054
rect 33852 30942 33854 30994
rect 33906 30942 33908 30994
rect 33852 30100 33908 30942
rect 34188 30884 34244 32396
rect 34300 31890 34356 37996
rect 34412 37268 34468 37278
rect 34412 34916 34468 37212
rect 34412 34860 34580 34916
rect 34412 34692 34468 34702
rect 34412 34598 34468 34636
rect 34524 32004 34580 34860
rect 34636 34242 34692 43148
rect 34748 42530 34804 42542
rect 34748 42478 34750 42530
rect 34802 42478 34804 42530
rect 34748 42308 34804 42478
rect 34748 41970 34804 42252
rect 34748 41918 34750 41970
rect 34802 41918 34804 41970
rect 34748 41906 34804 41918
rect 34748 40964 34804 40974
rect 34748 40626 34804 40908
rect 34748 40574 34750 40626
rect 34802 40574 34804 40626
rect 34748 40562 34804 40574
rect 34860 38668 34916 45164
rect 35084 44436 35140 47292
rect 35644 47236 35700 47246
rect 36204 47236 36260 47964
rect 36316 47954 36372 47964
rect 36652 48802 36708 50540
rect 36652 48750 36654 48802
rect 36706 48750 36708 48802
rect 36652 47796 36708 48750
rect 36652 47730 36708 47740
rect 36764 50596 36820 50606
rect 36764 48468 36820 50540
rect 37884 50596 37940 50606
rect 37996 50596 38052 52220
rect 37884 50594 38052 50596
rect 37884 50542 37886 50594
rect 37938 50542 38052 50594
rect 37884 50540 38052 50542
rect 38108 52164 38164 52780
rect 38332 52770 38388 52780
rect 38332 52276 38388 52286
rect 38388 52220 38500 52276
rect 38332 52182 38388 52220
rect 37884 50530 37940 50540
rect 36988 49700 37044 49710
rect 36988 49698 37156 49700
rect 36988 49646 36990 49698
rect 37042 49646 37156 49698
rect 36988 49644 37156 49646
rect 36988 49634 37044 49644
rect 36764 47570 36820 48412
rect 36988 48244 37044 48254
rect 36988 47796 37044 48188
rect 37100 48020 37156 49644
rect 37436 49698 37492 49710
rect 37436 49646 37438 49698
rect 37490 49646 37492 49698
rect 37436 48804 37492 49646
rect 37660 49700 37716 49710
rect 37548 48804 37604 48814
rect 37436 48802 37604 48804
rect 37436 48750 37550 48802
rect 37602 48750 37604 48802
rect 37436 48748 37604 48750
rect 37324 48468 37380 48478
rect 37324 48374 37380 48412
rect 37548 48244 37604 48748
rect 37548 48178 37604 48188
rect 37100 47954 37156 47964
rect 36988 47740 37380 47796
rect 36764 47518 36766 47570
rect 36818 47518 36820 47570
rect 36764 47506 36820 47518
rect 35644 47234 36260 47236
rect 35644 47182 35646 47234
rect 35698 47182 36260 47234
rect 35644 47180 36260 47182
rect 36316 47234 36372 47246
rect 36316 47182 36318 47234
rect 36370 47182 36372 47234
rect 35644 47124 35700 47180
rect 35644 47058 35700 47068
rect 36316 46676 36372 47182
rect 36988 46900 37044 46910
rect 36876 46788 36932 46798
rect 36988 46788 37044 46844
rect 36876 46786 37044 46788
rect 36876 46734 36878 46786
rect 36930 46734 37044 46786
rect 36876 46732 37044 46734
rect 36876 46722 36932 46732
rect 36316 46610 36372 46620
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35308 46004 35364 46014
rect 35196 46002 35364 46004
rect 35196 45950 35310 46002
rect 35362 45950 35364 46002
rect 35196 45948 35364 45950
rect 35196 45444 35252 45948
rect 35308 45938 35364 45948
rect 37212 45892 37268 45902
rect 36652 45780 36708 45790
rect 36652 45686 36708 45724
rect 35196 45378 35252 45388
rect 36540 45668 36596 45678
rect 35532 45220 35588 45230
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35084 44370 35140 44380
rect 35420 44324 35476 44334
rect 35532 44324 35588 45164
rect 36428 45220 36484 45230
rect 35476 44268 35588 44324
rect 36204 44884 36260 44894
rect 35420 44230 35476 44268
rect 35084 44212 35140 44222
rect 35084 44118 35140 44156
rect 36204 44212 36260 44828
rect 36428 44660 36484 45164
rect 36428 44594 36484 44604
rect 36316 44548 36372 44558
rect 36316 44454 36372 44492
rect 36428 44324 36484 44334
rect 36540 44324 36596 45612
rect 36428 44322 36596 44324
rect 36428 44270 36430 44322
rect 36482 44270 36596 44322
rect 36428 44268 36596 44270
rect 36652 45556 36708 45566
rect 36428 44258 36484 44268
rect 36316 44212 36372 44222
rect 36652 44212 36708 45500
rect 37212 45330 37268 45836
rect 37212 45278 37214 45330
rect 37266 45278 37268 45330
rect 37212 45266 37268 45278
rect 36260 44210 36372 44212
rect 36260 44158 36318 44210
rect 36370 44158 36372 44210
rect 36260 44156 36372 44158
rect 36204 44080 36260 44156
rect 35868 43652 35924 43662
rect 35868 43538 35924 43596
rect 35868 43486 35870 43538
rect 35922 43486 35924 43538
rect 35868 43474 35924 43486
rect 36316 43540 36372 44156
rect 36540 44156 36708 44212
rect 36428 43540 36484 43550
rect 36316 43538 36484 43540
rect 36316 43486 36430 43538
rect 36482 43486 36484 43538
rect 36316 43484 36484 43486
rect 36428 43474 36484 43484
rect 35084 43428 35140 43438
rect 35084 42756 35140 43372
rect 35420 43426 35476 43438
rect 35420 43374 35422 43426
rect 35474 43374 35476 43426
rect 35420 43316 35476 43374
rect 35420 43260 35700 43316
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35084 42700 35476 42756
rect 35420 42532 35476 42700
rect 35644 42644 35700 43260
rect 36092 42868 36148 42878
rect 35644 42642 35812 42644
rect 35644 42590 35646 42642
rect 35698 42590 35812 42642
rect 35644 42588 35812 42590
rect 35644 42578 35700 42588
rect 35420 42438 35476 42476
rect 35532 42530 35588 42542
rect 35532 42478 35534 42530
rect 35586 42478 35588 42530
rect 34972 41860 35028 41870
rect 34972 41766 35028 41804
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35420 41188 35476 41198
rect 35420 41094 35476 41132
rect 35532 41076 35588 42478
rect 35756 42084 35812 42588
rect 35868 42532 35924 42542
rect 35868 42194 35924 42476
rect 35868 42142 35870 42194
rect 35922 42142 35924 42194
rect 35868 42130 35924 42142
rect 36092 42308 36148 42812
rect 36092 42194 36148 42252
rect 36092 42142 36094 42194
rect 36146 42142 36148 42194
rect 35756 42018 35812 42028
rect 35980 42084 36036 42094
rect 35644 41972 35700 41982
rect 35644 41878 35700 41916
rect 35756 41858 35812 41870
rect 35756 41806 35758 41858
rect 35810 41806 35812 41858
rect 35756 41748 35812 41806
rect 35756 41682 35812 41692
rect 35980 41524 36036 42028
rect 35644 41468 36036 41524
rect 35644 41298 35700 41468
rect 35644 41246 35646 41298
rect 35698 41246 35700 41298
rect 35644 41234 35700 41246
rect 35532 41010 35588 41020
rect 35644 41074 35700 41086
rect 35644 41022 35646 41074
rect 35698 41022 35700 41074
rect 35308 40628 35364 40638
rect 35308 40402 35364 40572
rect 35308 40350 35310 40402
rect 35362 40350 35364 40402
rect 35308 40338 35364 40350
rect 35644 40404 35700 41022
rect 36092 41074 36148 42142
rect 36092 41022 36094 41074
rect 36146 41022 36148 41074
rect 36092 41010 36148 41022
rect 36316 41186 36372 41198
rect 36316 41134 36318 41186
rect 36370 41134 36372 41186
rect 36204 40628 36260 40638
rect 36204 40534 36260 40572
rect 36316 40626 36372 41134
rect 36316 40574 36318 40626
rect 36370 40574 36372 40626
rect 36316 40562 36372 40574
rect 36428 40740 36484 40750
rect 36428 40626 36484 40684
rect 36428 40574 36430 40626
rect 36482 40574 36484 40626
rect 35644 40338 35700 40348
rect 35756 40402 35812 40414
rect 35756 40350 35758 40402
rect 35810 40350 35812 40402
rect 35532 40292 35588 40302
rect 35084 40180 35140 40190
rect 35084 40086 35140 40124
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39396 35140 39406
rect 35084 38668 35140 39340
rect 35532 38836 35588 40236
rect 35644 39844 35700 39854
rect 35756 39844 35812 40350
rect 35644 39842 35812 39844
rect 35644 39790 35646 39842
rect 35698 39790 35812 39842
rect 35644 39788 35812 39790
rect 35644 39778 35700 39788
rect 36204 39732 36260 39742
rect 36428 39732 36484 40574
rect 36540 40292 36596 44156
rect 37324 44100 37380 47740
rect 37548 47458 37604 47470
rect 37548 47406 37550 47458
rect 37602 47406 37604 47458
rect 37548 46900 37604 47406
rect 37660 47348 37716 49644
rect 37884 49028 37940 49038
rect 37884 48934 37940 48972
rect 37772 48468 37828 48478
rect 37772 47458 37828 48412
rect 38108 47684 38164 52108
rect 38332 51604 38388 51614
rect 38332 51510 38388 51548
rect 38220 51492 38276 51502
rect 38220 50708 38276 51436
rect 38332 51380 38388 51390
rect 38444 51380 38500 52220
rect 38332 51378 38500 51380
rect 38332 51326 38334 51378
rect 38386 51326 38500 51378
rect 38332 51324 38500 51326
rect 38892 51940 38948 53006
rect 39004 52386 39060 53678
rect 39116 54402 39172 54460
rect 39116 54350 39118 54402
rect 39170 54350 39172 54402
rect 39116 53506 39172 54350
rect 39228 53844 39284 55132
rect 39340 55122 39396 55132
rect 39676 54738 39732 55244
rect 39788 55234 39844 55244
rect 40236 55234 40292 55244
rect 39676 54686 39678 54738
rect 39730 54686 39732 54738
rect 39676 54674 39732 54686
rect 40572 54738 40628 55244
rect 41132 55300 41188 55918
rect 41132 55234 41188 55244
rect 41244 55636 41300 55646
rect 40572 54686 40574 54738
rect 40626 54686 40628 54738
rect 40572 54674 40628 54686
rect 40796 54516 40852 54526
rect 40796 54422 40852 54460
rect 39340 54404 39396 54414
rect 39340 54310 39396 54348
rect 40460 54404 40516 54414
rect 39228 53778 39284 53788
rect 40460 53842 40516 54348
rect 40460 53790 40462 53842
rect 40514 53790 40516 53842
rect 40460 53778 40516 53790
rect 39340 53732 39396 53742
rect 39340 53638 39396 53676
rect 40348 53732 40404 53742
rect 40348 53638 40404 53676
rect 40460 53620 40516 53630
rect 40460 53526 40516 53564
rect 39116 53454 39118 53506
rect 39170 53454 39172 53506
rect 39116 52500 39172 53454
rect 40908 53172 40964 53182
rect 40908 53078 40964 53116
rect 40684 53060 40740 53070
rect 40684 53058 40852 53060
rect 40684 53006 40686 53058
rect 40738 53006 40852 53058
rect 40684 53004 40852 53006
rect 40684 52994 40740 53004
rect 39228 52948 39284 52958
rect 40572 52948 40628 52958
rect 39228 52946 39396 52948
rect 39228 52894 39230 52946
rect 39282 52894 39396 52946
rect 39228 52892 39396 52894
rect 39228 52882 39284 52892
rect 39116 52444 39284 52500
rect 39004 52334 39006 52386
rect 39058 52334 39060 52386
rect 39004 52322 39060 52334
rect 39116 52164 39172 52174
rect 38332 51314 38388 51324
rect 38780 51268 38836 51278
rect 38444 51154 38500 51166
rect 38444 51102 38446 51154
rect 38498 51102 38500 51154
rect 38444 50818 38500 51102
rect 38444 50766 38446 50818
rect 38498 50766 38500 50818
rect 38444 50754 38500 50766
rect 38668 51154 38724 51166
rect 38668 51102 38670 51154
rect 38722 51102 38724 51154
rect 38332 50708 38388 50718
rect 38220 50706 38388 50708
rect 38220 50654 38334 50706
rect 38386 50654 38388 50706
rect 38220 50652 38388 50654
rect 38220 50596 38276 50652
rect 38332 50642 38388 50652
rect 38220 50530 38276 50540
rect 38668 50484 38724 51102
rect 38668 50418 38724 50428
rect 38332 48802 38388 48814
rect 38332 48750 38334 48802
rect 38386 48750 38388 48802
rect 38332 48244 38388 48750
rect 38332 48178 38388 48188
rect 38108 47618 38164 47628
rect 38220 48130 38276 48142
rect 38220 48078 38222 48130
rect 38274 48078 38276 48130
rect 37772 47406 37774 47458
rect 37826 47406 37828 47458
rect 37772 47394 37828 47406
rect 37996 47458 38052 47470
rect 37996 47406 37998 47458
rect 38050 47406 38052 47458
rect 37660 47282 37716 47292
rect 37548 46834 37604 46844
rect 37772 47236 37828 47246
rect 37548 46674 37604 46686
rect 37548 46622 37550 46674
rect 37602 46622 37604 46674
rect 37548 46452 37604 46622
rect 37772 46674 37828 47180
rect 37772 46622 37774 46674
rect 37826 46622 37828 46674
rect 37772 46610 37828 46622
rect 37996 46676 38052 47406
rect 37996 46610 38052 46620
rect 38220 46452 38276 48078
rect 38668 48130 38724 48142
rect 38668 48078 38670 48130
rect 38722 48078 38724 48130
rect 38668 47460 38724 48078
rect 38668 47394 38724 47404
rect 37548 46396 38276 46452
rect 38332 46562 38388 46574
rect 38332 46510 38334 46562
rect 38386 46510 38388 46562
rect 37436 45668 37492 45678
rect 37436 45574 37492 45612
rect 37548 45220 37604 46396
rect 37660 46116 37716 46126
rect 37660 45666 37716 46060
rect 38332 46116 38388 46510
rect 38332 46050 38388 46060
rect 37772 45892 37828 45902
rect 37772 45798 37828 45836
rect 38780 45892 38836 51212
rect 38892 49924 38948 51884
rect 39004 52108 39116 52164
rect 39004 51604 39060 52108
rect 39116 52070 39172 52108
rect 39228 51940 39284 52444
rect 39004 51538 39060 51548
rect 39116 51884 39284 51940
rect 39004 50594 39060 50606
rect 39004 50542 39006 50594
rect 39058 50542 39060 50594
rect 39004 50372 39060 50542
rect 39004 50306 39060 50316
rect 38892 49868 39060 49924
rect 38892 49700 38948 49710
rect 38892 49606 38948 49644
rect 39004 49586 39060 49868
rect 39004 49534 39006 49586
rect 39058 49534 39060 49586
rect 39004 49522 39060 49534
rect 39116 47682 39172 51884
rect 39340 51492 39396 52892
rect 40348 52946 40628 52948
rect 40348 52894 40574 52946
rect 40626 52894 40628 52946
rect 40348 52892 40628 52894
rect 39788 52834 39844 52846
rect 39788 52782 39790 52834
rect 39842 52782 39844 52834
rect 39788 52724 39844 52782
rect 39788 52658 39844 52668
rect 39228 51436 39396 51492
rect 39788 52162 39844 52174
rect 39788 52110 39790 52162
rect 39842 52110 39844 52162
rect 39228 50484 39284 51436
rect 39340 51268 39396 51278
rect 39340 51174 39396 51212
rect 39676 51266 39732 51278
rect 39676 51214 39678 51266
rect 39730 51214 39732 51266
rect 39676 50428 39732 51214
rect 39788 50932 39844 52110
rect 40348 52052 40404 52892
rect 40572 52882 40628 52892
rect 40796 52386 40852 53004
rect 40796 52334 40798 52386
rect 40850 52334 40852 52386
rect 40460 52276 40516 52286
rect 40460 52182 40516 52220
rect 40236 51996 40348 52052
rect 40124 51380 40180 51390
rect 40124 51286 40180 51324
rect 39788 50866 39844 50876
rect 40012 51268 40068 51278
rect 40012 50820 40068 51212
rect 40124 50820 40180 50830
rect 40012 50818 40180 50820
rect 40012 50766 40126 50818
rect 40178 50766 40180 50818
rect 40012 50764 40180 50766
rect 40124 50754 40180 50764
rect 39228 50390 39284 50428
rect 39452 50372 39732 50428
rect 39340 49700 39396 49710
rect 39340 49606 39396 49644
rect 39228 49028 39284 49038
rect 39228 48934 39284 48972
rect 39340 48804 39396 48814
rect 39116 47630 39118 47682
rect 39170 47630 39172 47682
rect 39116 47618 39172 47630
rect 39228 48802 39396 48804
rect 39228 48750 39342 48802
rect 39394 48750 39396 48802
rect 39228 48748 39396 48750
rect 38780 45826 38836 45836
rect 39116 45892 39172 45902
rect 39116 45798 39172 45836
rect 39228 45892 39284 48748
rect 39340 48738 39396 48748
rect 39452 48804 39508 50372
rect 39676 50260 39732 50372
rect 39676 50194 39732 50204
rect 39788 50706 39844 50718
rect 39788 50654 39790 50706
rect 39842 50654 39844 50706
rect 39788 50372 39844 50654
rect 39788 49698 39844 50316
rect 39900 50482 39956 50494
rect 39900 50430 39902 50482
rect 39954 50430 39956 50482
rect 39900 50260 39956 50430
rect 40236 50428 40292 51996
rect 40348 51920 40404 51996
rect 40796 51716 40852 52334
rect 40908 52612 40964 52622
rect 40908 52274 40964 52556
rect 40908 52222 40910 52274
rect 40962 52222 40964 52274
rect 40908 52210 40964 52222
rect 40460 51660 40964 51716
rect 40348 51490 40404 51502
rect 40348 51438 40350 51490
rect 40402 51438 40404 51490
rect 40348 50596 40404 51438
rect 40460 51378 40516 51660
rect 40460 51326 40462 51378
rect 40514 51326 40516 51378
rect 40460 51314 40516 51326
rect 40348 50540 40852 50596
rect 39900 50194 39956 50204
rect 40124 50372 40292 50428
rect 39788 49646 39790 49698
rect 39842 49646 39844 49698
rect 39564 49586 39620 49598
rect 39564 49534 39566 49586
rect 39618 49534 39620 49586
rect 39564 48804 39620 49534
rect 39788 49028 39844 49646
rect 39900 49700 39956 49710
rect 39900 49250 39956 49644
rect 40012 49586 40068 49598
rect 40012 49534 40014 49586
rect 40066 49534 40068 49586
rect 40012 49364 40068 49534
rect 40012 49298 40068 49308
rect 39900 49198 39902 49250
rect 39954 49198 39956 49250
rect 39900 49186 39956 49198
rect 40124 49138 40180 50372
rect 40684 50370 40740 50382
rect 40684 50318 40686 50370
rect 40738 50318 40740 50370
rect 40684 49924 40740 50318
rect 40684 49858 40740 49868
rect 40460 49700 40516 49710
rect 40460 49606 40516 49644
rect 40124 49086 40126 49138
rect 40178 49086 40180 49138
rect 40124 49074 40180 49086
rect 40236 49586 40292 49598
rect 40236 49534 40238 49586
rect 40290 49534 40292 49586
rect 39788 48962 39844 48972
rect 40012 49026 40068 49038
rect 40012 48974 40014 49026
rect 40066 48974 40068 49026
rect 40012 48916 40068 48974
rect 40012 48804 40068 48860
rect 39564 48748 40068 48804
rect 40236 49028 40292 49534
rect 39452 48468 39508 48748
rect 39564 48468 39620 48478
rect 39452 48466 39620 48468
rect 39452 48414 39566 48466
rect 39618 48414 39620 48466
rect 39452 48412 39620 48414
rect 39564 48402 39620 48412
rect 39340 48242 39396 48254
rect 39340 48190 39342 48242
rect 39394 48190 39396 48242
rect 39340 46676 39396 48190
rect 40124 48242 40180 48254
rect 40124 48190 40126 48242
rect 40178 48190 40180 48242
rect 40124 48132 40180 48190
rect 40124 48066 40180 48076
rect 39452 47908 39508 47918
rect 39452 47458 39508 47852
rect 40236 47682 40292 48972
rect 40460 49364 40516 49374
rect 40460 49026 40516 49308
rect 40460 48974 40462 49026
rect 40514 48974 40516 49026
rect 40348 48244 40404 48254
rect 40348 48150 40404 48188
rect 40460 48020 40516 48974
rect 40684 49028 40740 49038
rect 40684 48934 40740 48972
rect 40796 48466 40852 50540
rect 40908 50034 40964 51660
rect 41020 51380 41076 51390
rect 41020 50594 41076 51324
rect 41020 50542 41022 50594
rect 41074 50542 41076 50594
rect 41020 50484 41076 50542
rect 41020 50418 41076 50428
rect 41132 50596 41188 50606
rect 41244 50596 41300 55580
rect 41580 54516 41636 56030
rect 42924 56082 42980 56094
rect 42924 56030 42926 56082
rect 42978 56030 42980 56082
rect 42476 55972 42532 55982
rect 42476 55878 42532 55916
rect 42924 55972 42980 56030
rect 43596 55972 43652 57036
rect 46956 56084 47012 56094
rect 43708 55972 43764 55982
rect 43596 55970 43764 55972
rect 43596 55918 43710 55970
rect 43762 55918 43764 55970
rect 43596 55916 43764 55918
rect 42924 55906 42980 55916
rect 43708 55906 43764 55916
rect 42588 55298 42644 55310
rect 42588 55246 42590 55298
rect 42642 55246 42644 55298
rect 42252 55188 42308 55198
rect 41580 54450 41636 54460
rect 42028 55186 42308 55188
rect 42028 55134 42254 55186
rect 42306 55134 42308 55186
rect 42028 55132 42308 55134
rect 41580 53844 41636 53854
rect 41580 53730 41636 53788
rect 41580 53678 41582 53730
rect 41634 53678 41636 53730
rect 41580 53666 41636 53678
rect 41692 53618 41748 53630
rect 41692 53566 41694 53618
rect 41746 53566 41748 53618
rect 41468 52946 41524 52958
rect 41468 52894 41470 52946
rect 41522 52894 41524 52946
rect 41356 52162 41412 52174
rect 41356 52110 41358 52162
rect 41410 52110 41412 52162
rect 41356 51940 41412 52110
rect 41468 52052 41524 52894
rect 41692 52834 41748 53566
rect 42028 53172 42084 55132
rect 42252 55122 42308 55132
rect 42140 54628 42196 54638
rect 42140 54534 42196 54572
rect 42476 54514 42532 54526
rect 42476 54462 42478 54514
rect 42530 54462 42532 54514
rect 42252 54404 42308 54414
rect 42252 54310 42308 54348
rect 42476 54404 42532 54462
rect 42476 54338 42532 54348
rect 42476 53506 42532 53518
rect 42476 53454 42478 53506
rect 42530 53454 42532 53506
rect 42476 53396 42532 53454
rect 42476 53330 42532 53340
rect 42588 53172 42644 55246
rect 43708 55300 43764 55310
rect 43708 55206 43764 55244
rect 44156 55188 44212 55198
rect 44156 55094 44212 55132
rect 46620 55188 46676 55198
rect 46620 55094 46676 55132
rect 46956 55186 47012 56028
rect 48412 55972 48468 59200
rect 50556 56476 50820 56486
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50556 56410 50820 56420
rect 54236 56196 54292 56206
rect 54236 56102 54292 56140
rect 48860 56084 48916 56094
rect 48860 55990 48916 56028
rect 48412 55906 48468 55916
rect 49532 55972 49588 55982
rect 49532 55878 49588 55916
rect 54460 55972 54516 59200
rect 54684 56196 54740 56206
rect 54684 56082 54740 56140
rect 57820 56196 57876 56206
rect 57820 56102 57876 56140
rect 59836 56196 59892 59200
rect 59836 56130 59892 56140
rect 54684 56030 54686 56082
rect 54738 56030 54740 56082
rect 54684 56018 54740 56030
rect 56700 56082 56756 56094
rect 56700 56030 56702 56082
rect 56754 56030 56756 56082
rect 54460 55906 54516 55916
rect 55468 55972 55524 55982
rect 55468 55878 55524 55916
rect 46956 55134 46958 55186
rect 47010 55134 47012 55186
rect 46956 55122 47012 55134
rect 49308 55636 49364 55646
rect 43708 54628 43764 54638
rect 42700 54516 42756 54526
rect 43260 54516 43316 54526
rect 42700 54514 42980 54516
rect 42700 54462 42702 54514
rect 42754 54462 42980 54514
rect 42700 54460 42980 54462
rect 42700 54450 42756 54460
rect 42028 53170 42532 53172
rect 42028 53118 42030 53170
rect 42082 53118 42532 53170
rect 42028 53116 42532 53118
rect 42028 53106 42084 53116
rect 41692 52782 41694 52834
rect 41746 52782 41748 52834
rect 41692 52770 41748 52782
rect 41804 52946 41860 52958
rect 41804 52894 41806 52946
rect 41858 52894 41860 52946
rect 41804 52386 41860 52894
rect 41804 52334 41806 52386
rect 41858 52334 41860 52386
rect 41804 52322 41860 52334
rect 42028 52612 42084 52622
rect 42028 52388 42084 52556
rect 42028 52256 42084 52332
rect 42140 52276 42196 52286
rect 41468 51986 41524 51996
rect 41356 51874 41412 51884
rect 41468 51492 41524 51502
rect 41468 51398 41524 51436
rect 42028 51268 42084 51278
rect 42028 51174 42084 51212
rect 41244 50540 41412 50596
rect 40908 49982 40910 50034
rect 40962 49982 40964 50034
rect 40908 49970 40964 49982
rect 40796 48414 40798 48466
rect 40850 48414 40852 48466
rect 40796 48402 40852 48414
rect 40236 47630 40238 47682
rect 40290 47630 40292 47682
rect 40236 47618 40292 47630
rect 40348 47964 40516 48020
rect 40572 48242 40628 48254
rect 40572 48190 40574 48242
rect 40626 48190 40628 48242
rect 39452 47406 39454 47458
rect 39506 47406 39508 47458
rect 39452 47394 39508 47406
rect 39676 47460 39732 47470
rect 39676 47366 39732 47404
rect 40236 47124 40292 47134
rect 39564 46786 39620 46798
rect 39564 46734 39566 46786
rect 39618 46734 39620 46786
rect 39564 46676 39620 46734
rect 39340 46674 39508 46676
rect 39340 46622 39342 46674
rect 39394 46622 39508 46674
rect 39340 46620 39508 46622
rect 39340 46610 39396 46620
rect 39340 45892 39396 45902
rect 39228 45836 39340 45892
rect 37660 45614 37662 45666
rect 37714 45614 37716 45666
rect 37660 45556 37716 45614
rect 37660 45490 37716 45500
rect 38220 45666 38276 45678
rect 38220 45614 38222 45666
rect 38274 45614 38276 45666
rect 38220 45444 38276 45614
rect 38780 45668 38836 45678
rect 39228 45668 39284 45836
rect 39340 45826 39396 45836
rect 38780 45574 38836 45612
rect 38892 45612 39284 45668
rect 38220 45378 38276 45388
rect 38892 45220 38948 45612
rect 37548 45164 37828 45220
rect 37660 44994 37716 45006
rect 37660 44942 37662 44994
rect 37714 44942 37716 44994
rect 37436 44100 37492 44110
rect 37324 44098 37492 44100
rect 37324 44046 37438 44098
rect 37490 44046 37492 44098
rect 37324 44044 37492 44046
rect 36652 43876 36708 43886
rect 36652 42868 36708 43820
rect 37436 43428 37492 44044
rect 37436 43362 37492 43372
rect 36652 42736 36708 42812
rect 36764 42756 36820 42766
rect 36540 40226 36596 40236
rect 36652 42532 36708 42542
rect 36652 42308 36708 42476
rect 36652 40068 36708 42252
rect 35756 39730 36484 39732
rect 35756 39678 36206 39730
rect 36258 39678 36484 39730
rect 35756 39676 36484 39678
rect 36540 39732 36596 39742
rect 35756 39618 35812 39676
rect 35756 39566 35758 39618
rect 35810 39566 35812 39618
rect 35756 39554 35812 39566
rect 35644 39508 35700 39518
rect 35644 39394 35700 39452
rect 35644 39342 35646 39394
rect 35698 39342 35700 39394
rect 35644 39284 35700 39342
rect 35644 39218 35700 39228
rect 35532 38834 35700 38836
rect 35532 38782 35534 38834
rect 35586 38782 35700 38834
rect 35532 38780 35700 38782
rect 35532 38770 35588 38780
rect 34748 38612 34916 38668
rect 34972 38612 35140 38668
rect 34748 37492 34804 38612
rect 34860 38164 34916 38202
rect 34860 38098 34916 38108
rect 34860 37940 34916 37978
rect 34860 37874 34916 37884
rect 34972 37604 35028 38612
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35308 37938 35364 37950
rect 35308 37886 35310 37938
rect 35362 37886 35364 37938
rect 35084 37828 35140 37838
rect 35084 37734 35140 37772
rect 34972 37548 35140 37604
rect 34748 37436 34916 37492
rect 34748 35588 34804 35598
rect 34748 35494 34804 35532
rect 34636 34190 34638 34242
rect 34690 34190 34692 34242
rect 34636 34178 34692 34190
rect 34524 31938 34580 31948
rect 34636 33348 34692 33358
rect 34636 33124 34692 33292
rect 34748 33124 34804 33134
rect 34636 33122 34804 33124
rect 34636 33070 34750 33122
rect 34802 33070 34804 33122
rect 34636 33068 34804 33070
rect 34300 31838 34302 31890
rect 34354 31838 34356 31890
rect 34300 31826 34356 31838
rect 34188 30790 34244 30828
rect 34300 30996 34356 31006
rect 33852 30034 33908 30044
rect 34188 30100 34244 30110
rect 33740 29810 33796 29820
rect 33516 29598 33518 29650
rect 33570 29598 33572 29650
rect 33516 29586 33572 29598
rect 33964 28756 34020 28766
rect 33964 28662 34020 28700
rect 33516 28644 33572 28654
rect 33516 28550 33572 28588
rect 33180 26852 33236 26862
rect 33180 24612 33236 26796
rect 33180 24546 33236 24556
rect 33292 26852 33460 26908
rect 33628 28196 33684 28206
rect 33068 24220 33236 24276
rect 33068 24050 33124 24062
rect 33068 23998 33070 24050
rect 33122 23998 33124 24050
rect 33068 23380 33124 23998
rect 33180 23604 33236 24220
rect 33292 24052 33348 26852
rect 33516 26180 33572 26190
rect 33404 26068 33460 26078
rect 33404 25284 33460 26012
rect 33516 25508 33572 26124
rect 33516 25442 33572 25452
rect 33404 25190 33460 25228
rect 33292 23986 33348 23996
rect 33404 24948 33460 24958
rect 33292 23828 33348 23838
rect 33292 23734 33348 23772
rect 33404 23604 33460 24892
rect 33516 24610 33572 24622
rect 33516 24558 33518 24610
rect 33570 24558 33572 24610
rect 33516 24500 33572 24558
rect 33516 24434 33572 24444
rect 33628 23940 33684 28140
rect 33852 28084 33908 28094
rect 33852 27298 33908 28028
rect 33852 27246 33854 27298
rect 33906 27246 33908 27298
rect 33852 27234 33908 27246
rect 34076 28084 34132 28094
rect 33964 26180 34020 26190
rect 33740 25394 33796 25406
rect 33740 25342 33742 25394
rect 33794 25342 33796 25394
rect 33740 24836 33796 25342
rect 33964 24946 34020 26124
rect 33964 24894 33966 24946
rect 34018 24894 34020 24946
rect 33964 24882 34020 24894
rect 33740 24770 33796 24780
rect 33852 24500 33908 24510
rect 33628 23884 33796 23940
rect 33516 23828 33572 23838
rect 33516 23734 33572 23772
rect 33628 23714 33684 23726
rect 33628 23662 33630 23714
rect 33682 23662 33684 23714
rect 33628 23604 33684 23662
rect 33180 23548 33348 23604
rect 33404 23548 33628 23604
rect 33068 23314 33124 23324
rect 32844 23202 32900 23212
rect 32956 23156 33012 23166
rect 32956 23154 33124 23156
rect 32956 23102 32958 23154
rect 33010 23102 33124 23154
rect 32956 23100 33124 23102
rect 32956 23090 33012 23100
rect 32956 22932 33012 22942
rect 32732 21970 32788 21980
rect 32844 22148 32900 22158
rect 32508 21698 32676 21700
rect 32508 21646 32510 21698
rect 32562 21646 32676 21698
rect 32508 21644 32676 21646
rect 32508 21634 32564 21644
rect 32620 21026 32676 21644
rect 32620 20974 32622 21026
rect 32674 20974 32676 21026
rect 32620 20692 32676 20974
rect 32844 21698 32900 22092
rect 32844 21646 32846 21698
rect 32898 21646 32900 21698
rect 32732 20916 32788 20926
rect 32844 20916 32900 21646
rect 32732 20914 32900 20916
rect 32732 20862 32734 20914
rect 32786 20862 32900 20914
rect 32732 20860 32900 20862
rect 32732 20850 32788 20860
rect 32956 20804 33012 22876
rect 33068 20914 33124 23100
rect 33180 22148 33236 22158
rect 33180 22054 33236 22092
rect 33068 20862 33070 20914
rect 33122 20862 33124 20914
rect 33068 20850 33124 20862
rect 32844 20748 33012 20804
rect 32620 20636 32788 20692
rect 32508 20580 32564 20590
rect 32508 20130 32564 20524
rect 32508 20078 32510 20130
rect 32562 20078 32564 20130
rect 32508 20066 32564 20078
rect 32508 19012 32564 19050
rect 32508 18946 32564 18956
rect 32508 18788 32564 18798
rect 32508 18562 32564 18732
rect 32508 18510 32510 18562
rect 32562 18510 32564 18562
rect 32508 18498 32564 18510
rect 32620 18676 32676 18686
rect 32620 18450 32676 18620
rect 32620 18398 32622 18450
rect 32674 18398 32676 18450
rect 32508 17780 32564 17790
rect 32620 17780 32676 18398
rect 32732 18228 32788 20636
rect 32732 18162 32788 18172
rect 32508 17778 32676 17780
rect 32508 17726 32510 17778
rect 32562 17726 32676 17778
rect 32508 17724 32676 17726
rect 32508 17714 32564 17724
rect 32732 17666 32788 17678
rect 32732 17614 32734 17666
rect 32786 17614 32788 17666
rect 32732 17444 32788 17614
rect 32732 17378 32788 17388
rect 32732 16996 32788 17006
rect 32508 16884 32564 16894
rect 32508 16790 32564 16828
rect 32732 16882 32788 16940
rect 32732 16830 32734 16882
rect 32786 16830 32788 16882
rect 32620 15988 32676 15998
rect 32732 15988 32788 16830
rect 32620 15986 32788 15988
rect 32620 15934 32622 15986
rect 32674 15934 32788 15986
rect 32620 15932 32788 15934
rect 32620 15922 32676 15932
rect 31724 15446 31780 15484
rect 31948 15484 32452 15540
rect 32508 15540 32564 15550
rect 31388 15092 31556 15148
rect 31276 14590 31278 14642
rect 31330 14590 31332 14642
rect 31276 14578 31332 14590
rect 31388 13636 31444 13646
rect 31388 13542 31444 13580
rect 31276 12964 31332 12974
rect 31276 12870 31332 12908
rect 31164 12292 31220 12302
rect 31164 12198 31220 12236
rect 31500 10612 31556 15092
rect 31724 14306 31780 14318
rect 31724 14254 31726 14306
rect 31778 14254 31780 14306
rect 31724 14084 31780 14254
rect 31724 14018 31780 14028
rect 31948 13524 32004 15484
rect 32508 15446 32564 15484
rect 32284 15316 32340 15326
rect 32284 15222 32340 15260
rect 31948 13458 32004 13468
rect 32396 15202 32452 15214
rect 32396 15150 32398 15202
rect 32450 15150 32452 15202
rect 31500 10546 31556 10556
rect 31052 5170 31108 5180
rect 32396 5236 32452 15150
rect 32844 13074 32900 20748
rect 33180 20690 33236 20702
rect 33180 20638 33182 20690
rect 33234 20638 33236 20690
rect 33180 20468 33236 20638
rect 33180 20402 33236 20412
rect 33292 20244 33348 23548
rect 33628 23472 33684 23548
rect 33628 23380 33684 23390
rect 33516 23268 33572 23278
rect 33516 23174 33572 23212
rect 33516 22260 33572 22270
rect 33516 22166 33572 22204
rect 33628 21812 33684 23324
rect 33740 21924 33796 23884
rect 33852 23938 33908 24444
rect 33852 23886 33854 23938
rect 33906 23886 33908 23938
rect 33852 23874 33908 23886
rect 33964 23604 34020 23614
rect 33964 23378 34020 23548
rect 33964 23326 33966 23378
rect 34018 23326 34020 23378
rect 33964 23314 34020 23326
rect 34076 21924 34132 28028
rect 34188 27970 34244 30044
rect 34188 27918 34190 27970
rect 34242 27918 34244 27970
rect 34188 27906 34244 27918
rect 34300 29314 34356 30940
rect 34412 30772 34468 30782
rect 34636 30772 34692 33068
rect 34748 33058 34804 33068
rect 34860 32788 34916 37436
rect 34972 33906 35028 33918
rect 34972 33854 34974 33906
rect 35026 33854 35028 33906
rect 34972 33572 35028 33854
rect 34972 33506 35028 33516
rect 34748 32732 34916 32788
rect 34748 31556 34804 32732
rect 34972 32450 35028 32462
rect 34972 32398 34974 32450
rect 35026 32398 35028 32450
rect 34860 31780 34916 31790
rect 34860 31686 34916 31724
rect 34972 31556 35028 32398
rect 34748 31500 34916 31556
rect 34412 30770 34692 30772
rect 34412 30718 34414 30770
rect 34466 30718 34692 30770
rect 34412 30716 34692 30718
rect 34748 30884 34804 30894
rect 34412 30100 34468 30716
rect 34748 30324 34804 30828
rect 34748 30210 34804 30268
rect 34748 30158 34750 30210
rect 34802 30158 34804 30210
rect 34748 30146 34804 30158
rect 34412 30034 34468 30044
rect 34524 29988 34580 29998
rect 34524 29876 34580 29932
rect 34300 29262 34302 29314
rect 34354 29262 34356 29314
rect 34188 27746 34244 27758
rect 34188 27694 34190 27746
rect 34242 27694 34244 27746
rect 34188 27300 34244 27694
rect 34188 27168 34244 27244
rect 33740 21868 33908 21924
rect 33628 21756 33796 21812
rect 33404 21700 33460 21710
rect 33404 20916 33460 21644
rect 33404 20802 33460 20860
rect 33404 20750 33406 20802
rect 33458 20750 33460 20802
rect 33404 20738 33460 20750
rect 33628 20580 33684 20618
rect 33628 20514 33684 20524
rect 33068 20188 33348 20244
rect 33628 20356 33684 20366
rect 33628 20242 33684 20300
rect 33628 20190 33630 20242
rect 33682 20190 33684 20242
rect 32956 19906 33012 19918
rect 32956 19854 32958 19906
rect 33010 19854 33012 19906
rect 32956 19796 33012 19854
rect 32956 19730 33012 19740
rect 32956 19236 33012 19246
rect 32956 19142 33012 19180
rect 33068 17780 33124 20188
rect 33628 20020 33684 20190
rect 33404 19964 33684 20020
rect 33404 19346 33460 19964
rect 33404 19294 33406 19346
rect 33458 19294 33460 19346
rect 33404 19282 33460 19294
rect 33516 19794 33572 19806
rect 33516 19742 33518 19794
rect 33570 19742 33572 19794
rect 33068 17714 33124 17724
rect 33404 17780 33460 17790
rect 33180 17444 33236 17454
rect 33068 17332 33124 17342
rect 32956 15988 33012 15998
rect 32956 15894 33012 15932
rect 32956 15316 33012 15326
rect 32956 15222 33012 15260
rect 32844 13022 32846 13074
rect 32898 13022 32900 13074
rect 32844 12964 32900 13022
rect 32844 12898 32900 12908
rect 32396 5170 32452 5180
rect 32844 12292 32900 12302
rect 32844 12066 32900 12236
rect 32844 12014 32846 12066
rect 32898 12014 32900 12066
rect 31052 4116 31108 4126
rect 31052 3666 31108 4060
rect 31052 3614 31054 3666
rect 31106 3614 31108 3666
rect 30492 3556 30548 3566
rect 29372 3444 29428 3482
rect 30492 3462 30548 3500
rect 31052 3556 31108 3614
rect 31052 3490 31108 3500
rect 29372 3378 29428 3388
rect 32844 2772 32900 12014
rect 33068 11396 33124 17276
rect 33180 12964 33236 17388
rect 33292 12964 33348 12974
rect 33180 12962 33348 12964
rect 33180 12910 33294 12962
rect 33346 12910 33348 12962
rect 33180 12908 33348 12910
rect 33292 12852 33348 12908
rect 33292 12786 33348 12796
rect 33068 11330 33124 11340
rect 33404 8148 33460 17724
rect 33516 17666 33572 19742
rect 33740 19124 33796 21756
rect 33852 20804 33908 21868
rect 34076 21858 34132 21868
rect 34188 25396 34244 25406
rect 34076 21700 34132 21710
rect 34076 21606 34132 21644
rect 33964 21588 34020 21598
rect 33964 21494 34020 21532
rect 34188 21474 34244 25340
rect 34300 24948 34356 29262
rect 34412 29820 34580 29876
rect 34412 28308 34468 29820
rect 34636 29426 34692 29438
rect 34636 29374 34638 29426
rect 34690 29374 34692 29426
rect 34524 28532 34580 28542
rect 34524 28438 34580 28476
rect 34412 28252 34580 28308
rect 34412 27858 34468 27870
rect 34412 27806 34414 27858
rect 34466 27806 34468 27858
rect 34412 26964 34468 27806
rect 34524 27748 34580 28252
rect 34636 27972 34692 29374
rect 34748 28980 34804 28990
rect 34748 28644 34804 28924
rect 34748 28530 34804 28588
rect 34748 28478 34750 28530
rect 34802 28478 34804 28530
rect 34748 28466 34804 28478
rect 34636 27906 34692 27916
rect 34524 27692 34804 27748
rect 34412 26898 34468 26908
rect 34524 27300 34580 27310
rect 34412 26402 34468 26414
rect 34412 26350 34414 26402
rect 34466 26350 34468 26402
rect 34412 26180 34468 26350
rect 34412 26114 34468 26124
rect 34524 25618 34580 27244
rect 34748 26514 34804 27692
rect 34860 26908 34916 31500
rect 34972 31490 35028 31500
rect 34972 30884 35028 30894
rect 34972 30790 35028 30828
rect 35084 30660 35140 37548
rect 35308 37490 35364 37886
rect 35644 37940 35700 38780
rect 35644 37874 35700 37884
rect 35308 37438 35310 37490
rect 35362 37438 35364 37490
rect 35308 37426 35364 37438
rect 35756 37044 35812 37054
rect 35756 36950 35812 36988
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35868 36148 35924 39676
rect 36204 39666 36260 39676
rect 36092 38834 36148 38846
rect 36092 38782 36094 38834
rect 36146 38782 36148 38834
rect 35980 38052 36036 38062
rect 36092 38052 36148 38782
rect 36316 38834 36372 38846
rect 36316 38782 36318 38834
rect 36370 38782 36372 38834
rect 36204 38722 36260 38734
rect 36204 38670 36206 38722
rect 36258 38670 36260 38722
rect 36204 38276 36260 38670
rect 36204 38210 36260 38220
rect 35980 38050 36148 38052
rect 35980 37998 35982 38050
rect 36034 37998 36148 38050
rect 35980 37996 36148 37998
rect 35980 37986 36036 37996
rect 35532 36092 35924 36148
rect 35980 37716 36036 37726
rect 35980 37042 36036 37660
rect 35980 36990 35982 37042
rect 36034 36990 36036 37042
rect 35308 35700 35364 35710
rect 35308 35606 35364 35644
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 34018 35252 34030
rect 35196 33966 35198 34018
rect 35250 33966 35252 34018
rect 35196 33906 35252 33966
rect 35196 33854 35198 33906
rect 35250 33854 35252 33906
rect 35196 33842 35252 33854
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35308 33572 35364 33582
rect 35308 32786 35364 33516
rect 35308 32734 35310 32786
rect 35362 32734 35364 32786
rect 35308 32722 35364 32734
rect 35420 33122 35476 33134
rect 35420 33070 35422 33122
rect 35474 33070 35476 33122
rect 35420 32340 35476 33070
rect 35532 32788 35588 36092
rect 35644 35924 35700 35934
rect 35980 35924 36036 36990
rect 35644 35922 36036 35924
rect 35644 35870 35646 35922
rect 35698 35870 36036 35922
rect 35644 35868 36036 35870
rect 35644 35858 35700 35868
rect 36092 35138 36148 37996
rect 36204 38052 36260 38062
rect 36316 38052 36372 38782
rect 36540 38162 36596 39676
rect 36652 39508 36708 40012
rect 36652 39414 36708 39452
rect 36764 42082 36820 42700
rect 37660 42756 37716 44942
rect 37660 42662 37716 42700
rect 37212 42644 37268 42654
rect 36988 42196 37044 42206
rect 36988 42102 37044 42140
rect 36764 42030 36766 42082
rect 36818 42030 36820 42082
rect 36764 39172 36820 42030
rect 37100 41972 37156 41982
rect 37100 41878 37156 41916
rect 36876 41300 36932 41310
rect 36876 40628 36932 41244
rect 36876 40496 36932 40572
rect 36540 38110 36542 38162
rect 36594 38110 36596 38162
rect 36540 38098 36596 38110
rect 36652 39116 36820 39172
rect 36204 38050 36372 38052
rect 36204 37998 36206 38050
rect 36258 37998 36372 38050
rect 36204 37996 36372 37998
rect 36204 37716 36260 37996
rect 36204 37650 36260 37660
rect 36540 37940 36596 37950
rect 36204 37268 36260 37278
rect 36540 37268 36596 37884
rect 36204 37266 36596 37268
rect 36204 37214 36206 37266
rect 36258 37214 36596 37266
rect 36204 37212 36596 37214
rect 36204 37202 36260 37212
rect 36092 35086 36094 35138
rect 36146 35086 36148 35138
rect 36092 35074 36148 35086
rect 36204 37044 36260 37054
rect 36204 36260 36260 36988
rect 36428 36260 36484 36270
rect 36204 36258 36484 36260
rect 36204 36206 36430 36258
rect 36482 36206 36484 36258
rect 36204 36204 36484 36206
rect 36092 34916 36148 34926
rect 35644 34914 36148 34916
rect 35644 34862 36094 34914
rect 36146 34862 36148 34914
rect 35644 34860 36148 34862
rect 35644 34690 35700 34860
rect 36092 34850 36148 34860
rect 35644 34638 35646 34690
rect 35698 34638 35700 34690
rect 35644 33124 35700 34638
rect 36092 34580 36148 34590
rect 35868 34018 35924 34030
rect 35868 33966 35870 34018
rect 35922 33966 35924 34018
rect 35868 33684 35924 33966
rect 35868 33618 35924 33628
rect 35980 33124 36036 33134
rect 35644 33122 36036 33124
rect 35644 33070 35982 33122
rect 36034 33070 36036 33122
rect 35644 33068 36036 33070
rect 35532 32732 35700 32788
rect 35532 32564 35588 32574
rect 35532 32470 35588 32508
rect 35420 32284 35588 32340
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35532 32004 35588 32284
rect 35308 31948 35588 32004
rect 35308 30996 35364 31948
rect 35308 30930 35364 30940
rect 35420 31666 35476 31678
rect 35420 31614 35422 31666
rect 35474 31614 35476 31666
rect 35420 31556 35476 31614
rect 35420 30772 35476 31500
rect 35532 31554 35588 31566
rect 35532 31502 35534 31554
rect 35586 31502 35588 31554
rect 35532 31444 35588 31502
rect 35532 31378 35588 31388
rect 35644 31220 35700 32732
rect 35868 32004 35924 32014
rect 35756 31780 35812 31790
rect 35756 31686 35812 31724
rect 35420 30706 35476 30716
rect 35532 31164 35700 31220
rect 35756 31220 35812 31230
rect 35868 31220 35924 31948
rect 35756 31218 35924 31220
rect 35756 31166 35758 31218
rect 35810 31166 35924 31218
rect 35756 31164 35924 31166
rect 34972 30604 35140 30660
rect 35196 30604 35460 30614
rect 34972 28754 35028 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 30210 35140 30222
rect 35084 30158 35086 30210
rect 35138 30158 35140 30210
rect 35084 30100 35140 30158
rect 35084 29652 35140 30044
rect 35196 29652 35252 29662
rect 35084 29650 35252 29652
rect 35084 29598 35198 29650
rect 35250 29598 35252 29650
rect 35084 29596 35252 29598
rect 35084 28868 35140 29596
rect 35196 29586 35252 29596
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35532 28868 35588 31164
rect 35644 30996 35700 31006
rect 35644 30902 35700 30940
rect 35756 30212 35812 31164
rect 35756 30146 35812 30156
rect 35644 30100 35700 30110
rect 35644 29876 35700 30044
rect 35644 29810 35700 29820
rect 35084 28802 35140 28812
rect 35420 28812 35588 28868
rect 34972 28702 34974 28754
rect 35026 28702 35028 28754
rect 34972 28690 35028 28702
rect 35196 28756 35252 28766
rect 35084 28532 35140 28542
rect 34972 28418 35028 28430
rect 34972 28366 34974 28418
rect 35026 28366 35028 28418
rect 34972 27972 35028 28366
rect 34972 27906 35028 27916
rect 35084 27188 35140 28476
rect 35196 27858 35252 28700
rect 35196 27806 35198 27858
rect 35250 27806 35252 27858
rect 35196 27794 35252 27806
rect 35420 27636 35476 28812
rect 35644 28756 35700 28766
rect 35532 28700 35644 28756
rect 35532 28642 35588 28700
rect 35644 28690 35700 28700
rect 35532 28590 35534 28642
rect 35586 28590 35588 28642
rect 35532 28578 35588 28590
rect 35868 28644 35924 28654
rect 35868 28550 35924 28588
rect 35868 28420 35924 28430
rect 35532 27972 35588 27982
rect 35532 27878 35588 27916
rect 35756 27972 35812 27982
rect 35420 27580 35588 27636
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35532 27300 35588 27580
rect 35420 27244 35588 27300
rect 35196 27188 35252 27198
rect 35084 27186 35252 27188
rect 35084 27134 35198 27186
rect 35250 27134 35252 27186
rect 35084 27132 35252 27134
rect 35196 27076 35252 27132
rect 35196 27010 35252 27020
rect 34860 26852 35140 26908
rect 34748 26462 34750 26514
rect 34802 26462 34804 26514
rect 34748 26450 34804 26462
rect 34636 26292 34692 26302
rect 34860 26292 34916 26302
rect 34636 26290 34804 26292
rect 34636 26238 34638 26290
rect 34690 26238 34804 26290
rect 34636 26236 34804 26238
rect 34636 26226 34692 26236
rect 34524 25566 34526 25618
rect 34578 25566 34580 25618
rect 34524 25554 34580 25566
rect 34412 25508 34468 25518
rect 34412 25414 34468 25452
rect 34300 24882 34356 24892
rect 34636 25282 34692 25294
rect 34636 25230 34638 25282
rect 34690 25230 34692 25282
rect 34412 24836 34468 24846
rect 34412 24742 34468 24780
rect 34636 24836 34692 25230
rect 34636 24770 34692 24780
rect 34748 24612 34804 26236
rect 34860 26290 35028 26292
rect 34860 26238 34862 26290
rect 34914 26238 35028 26290
rect 34860 26236 35028 26238
rect 34860 26226 34916 26236
rect 34860 25506 34916 25518
rect 34860 25454 34862 25506
rect 34914 25454 34916 25506
rect 34860 25396 34916 25454
rect 34860 25330 34916 25340
rect 34972 24836 35028 26236
rect 35084 25732 35140 26852
rect 35420 26852 35476 27244
rect 35420 26786 35476 26796
rect 35756 26850 35812 27916
rect 35756 26798 35758 26850
rect 35810 26798 35812 26850
rect 35756 26786 35812 26798
rect 35644 26740 35700 26750
rect 35420 26628 35476 26638
rect 35644 26628 35700 26684
rect 35644 26572 35812 26628
rect 35420 26402 35476 26572
rect 35420 26350 35422 26402
rect 35474 26350 35476 26402
rect 35420 26338 35476 26350
rect 35532 26404 35588 26414
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35532 25732 35588 26348
rect 35084 25676 35252 25732
rect 35084 25506 35140 25518
rect 35084 25454 35086 25506
rect 35138 25454 35140 25506
rect 35084 25284 35140 25454
rect 35084 25218 35140 25228
rect 35084 24836 35140 24846
rect 34748 24546 34804 24556
rect 34860 24834 35140 24836
rect 34860 24782 35086 24834
rect 35138 24782 35140 24834
rect 34860 24780 35140 24782
rect 34300 23828 34356 23838
rect 34300 23734 34356 23772
rect 34636 23828 34692 23838
rect 34636 23734 34692 23772
rect 34524 23714 34580 23726
rect 34524 23662 34526 23714
rect 34578 23662 34580 23714
rect 34188 21422 34190 21474
rect 34242 21422 34244 21474
rect 34188 21410 34244 21422
rect 34300 23604 34356 23614
rect 34300 22258 34356 23548
rect 34524 23604 34580 23662
rect 34524 23538 34580 23548
rect 34524 23154 34580 23166
rect 34524 23102 34526 23154
rect 34578 23102 34580 23154
rect 34524 22932 34580 23102
rect 34748 23154 34804 23166
rect 34748 23102 34750 23154
rect 34802 23102 34804 23154
rect 34636 23044 34692 23054
rect 34636 22950 34692 22988
rect 34524 22866 34580 22876
rect 34524 22596 34580 22606
rect 34748 22596 34804 23102
rect 34524 22594 34748 22596
rect 34524 22542 34526 22594
rect 34578 22542 34748 22594
rect 34524 22540 34748 22542
rect 34524 22530 34580 22540
rect 34748 22464 34804 22540
rect 34860 22372 34916 24780
rect 35084 24770 35140 24780
rect 35196 24612 35252 25676
rect 35532 25666 35588 25676
rect 35644 26292 35700 26302
rect 35532 25396 35588 25406
rect 35644 25396 35700 26236
rect 35756 26068 35812 26572
rect 35868 26514 35924 28364
rect 35980 26628 36036 33068
rect 36092 32564 36148 34524
rect 36204 33124 36260 36204
rect 36428 36194 36484 36204
rect 36316 35924 36372 35934
rect 36316 35810 36372 35868
rect 36316 35758 36318 35810
rect 36370 35758 36372 35810
rect 36316 35140 36372 35758
rect 36428 35812 36484 35822
rect 36428 35718 36484 35756
rect 36428 35476 36484 35486
rect 36428 35474 36596 35476
rect 36428 35422 36430 35474
rect 36482 35422 36596 35474
rect 36428 35420 36596 35422
rect 36428 35410 36484 35420
rect 36428 35140 36484 35150
rect 36316 35138 36484 35140
rect 36316 35086 36430 35138
rect 36482 35086 36484 35138
rect 36316 35084 36484 35086
rect 36428 35074 36484 35084
rect 36316 34130 36372 34142
rect 36316 34078 36318 34130
rect 36370 34078 36372 34130
rect 36316 33908 36372 34078
rect 36316 33842 36372 33852
rect 36316 33684 36372 33694
rect 36316 33346 36372 33628
rect 36316 33294 36318 33346
rect 36370 33294 36372 33346
rect 36316 33282 36372 33294
rect 36204 33068 36372 33124
rect 36092 32498 36148 32508
rect 36204 32116 36260 32126
rect 36092 29204 36148 29214
rect 36092 29110 36148 29148
rect 36092 28756 36148 28766
rect 36092 27186 36148 28700
rect 36204 27636 36260 32060
rect 36316 31780 36372 33068
rect 36428 32564 36484 32574
rect 36428 32004 36484 32508
rect 36428 31938 36484 31948
rect 36540 31892 36596 35420
rect 36540 31826 36596 31836
rect 36652 31890 36708 39116
rect 37100 39060 37156 39070
rect 37212 39060 37268 42588
rect 37548 42532 37604 42542
rect 37324 42530 37604 42532
rect 37324 42478 37550 42530
rect 37602 42478 37604 42530
rect 37324 42476 37604 42478
rect 37324 42082 37380 42476
rect 37548 42466 37604 42476
rect 37772 42308 37828 45164
rect 38780 45164 38948 45220
rect 38556 45108 38612 45118
rect 38332 44996 38388 45006
rect 38332 44994 38500 44996
rect 38332 44942 38334 44994
rect 38386 44942 38500 44994
rect 38332 44940 38500 44942
rect 38332 44930 38388 44940
rect 37996 44100 38052 44110
rect 37996 44098 38164 44100
rect 37996 44046 37998 44098
rect 38050 44046 38164 44098
rect 37996 44044 38164 44046
rect 37996 44034 38052 44044
rect 37996 43764 38052 43774
rect 37884 42754 37940 42766
rect 37884 42702 37886 42754
rect 37938 42702 37940 42754
rect 37884 42532 37940 42702
rect 37884 42466 37940 42476
rect 37772 42252 37940 42308
rect 37324 42030 37326 42082
rect 37378 42030 37380 42082
rect 37324 42018 37380 42030
rect 37772 41972 37828 41982
rect 37660 41916 37772 41972
rect 37548 40962 37604 40974
rect 37548 40910 37550 40962
rect 37602 40910 37604 40962
rect 37324 40290 37380 40302
rect 37324 40238 37326 40290
rect 37378 40238 37380 40290
rect 37324 40180 37380 40238
rect 37324 40114 37380 40124
rect 37548 39396 37604 40910
rect 37548 39330 37604 39340
rect 37100 39058 37268 39060
rect 37100 39006 37102 39058
rect 37154 39006 37268 39058
rect 37100 39004 37268 39006
rect 37100 38994 37156 39004
rect 36764 38836 36820 38846
rect 36764 38742 36820 38780
rect 36764 38276 36820 38286
rect 36764 38182 36820 38220
rect 37212 37940 37268 39004
rect 37660 38836 37716 41916
rect 37772 41878 37828 41916
rect 37884 41748 37940 42252
rect 37996 42194 38052 43708
rect 38108 42308 38164 44044
rect 38332 44098 38388 44110
rect 38332 44046 38334 44098
rect 38386 44046 38388 44098
rect 38332 42756 38388 44046
rect 38444 43764 38500 44940
rect 38444 43698 38500 43708
rect 38444 42980 38500 42990
rect 38556 42980 38612 45052
rect 38780 44772 38836 45164
rect 38892 44996 38948 45006
rect 38892 44994 39060 44996
rect 38892 44942 38894 44994
rect 38946 44942 39060 44994
rect 38892 44940 39060 44942
rect 38892 44930 38948 44940
rect 38780 44716 38948 44772
rect 38668 44660 38724 44670
rect 38668 43764 38724 44604
rect 38892 44210 38948 44716
rect 38892 44158 38894 44210
rect 38946 44158 38948 44210
rect 38892 44146 38948 44158
rect 38780 44098 38836 44110
rect 38780 44046 38782 44098
rect 38834 44046 38836 44098
rect 38780 43988 38836 44046
rect 38780 43922 38836 43932
rect 38780 43764 38836 43774
rect 38668 43762 38836 43764
rect 38668 43710 38782 43762
rect 38834 43710 38836 43762
rect 38668 43708 38836 43710
rect 38780 43698 38836 43708
rect 38892 43316 38948 43326
rect 38444 42978 38724 42980
rect 38444 42926 38446 42978
rect 38498 42926 38724 42978
rect 38444 42924 38724 42926
rect 38444 42914 38500 42924
rect 38332 42690 38388 42700
rect 38556 42756 38612 42766
rect 38220 42644 38276 42654
rect 38220 42550 38276 42588
rect 38108 42242 38164 42252
rect 37996 42142 37998 42194
rect 38050 42142 38052 42194
rect 37996 42130 38052 42142
rect 38108 42084 38164 42094
rect 38556 42084 38612 42700
rect 38108 42082 38612 42084
rect 38108 42030 38110 42082
rect 38162 42030 38612 42082
rect 38108 42028 38612 42030
rect 38108 42018 38164 42028
rect 37772 41692 37940 41748
rect 38556 41748 38612 42028
rect 38668 41970 38724 42924
rect 38892 42532 38948 43260
rect 39004 42644 39060 44940
rect 39340 44210 39396 44222
rect 39340 44158 39342 44210
rect 39394 44158 39396 44210
rect 39116 44100 39172 44110
rect 39172 44044 39284 44100
rect 39116 43968 39172 44044
rect 39004 42578 39060 42588
rect 38892 42466 38948 42476
rect 38892 42196 38948 42206
rect 38892 42102 38948 42140
rect 38668 41918 38670 41970
rect 38722 41918 38724 41970
rect 38668 41906 38724 41918
rect 38892 41972 38948 41982
rect 38556 41692 38724 41748
rect 37772 39844 37828 41692
rect 37884 41300 37940 41310
rect 37884 41206 37940 41244
rect 38108 41188 38164 41198
rect 37772 39778 37828 39788
rect 37996 40402 38052 40414
rect 37996 40350 37998 40402
rect 38050 40350 38052 40402
rect 37772 39508 37828 39518
rect 37772 39414 37828 39452
rect 37884 39396 37940 39406
rect 37884 39302 37940 39340
rect 37436 38724 37492 38734
rect 37436 38050 37492 38668
rect 37436 37998 37438 38050
rect 37490 37998 37492 38050
rect 37436 37986 37492 37998
rect 37660 37940 37716 38780
rect 37996 38834 38052 40350
rect 38108 39618 38164 41132
rect 38668 41186 38724 41692
rect 38668 41134 38670 41186
rect 38722 41134 38724 41186
rect 38668 41122 38724 41134
rect 38892 41188 38948 41916
rect 39116 41970 39172 41982
rect 39116 41918 39118 41970
rect 39170 41918 39172 41970
rect 39116 41298 39172 41918
rect 39228 41746 39284 44044
rect 39340 43428 39396 44158
rect 39452 43764 39508 46620
rect 39564 46610 39620 46620
rect 40012 46676 40068 46686
rect 40012 45778 40068 46620
rect 40236 46674 40292 47068
rect 40348 46900 40404 47964
rect 40460 46900 40516 46910
rect 40348 46898 40516 46900
rect 40348 46846 40462 46898
rect 40514 46846 40516 46898
rect 40348 46844 40516 46846
rect 40572 46900 40628 48190
rect 40796 48242 40852 48254
rect 40796 48190 40798 48242
rect 40850 48190 40852 48242
rect 40684 48132 40740 48142
rect 40684 47458 40740 48076
rect 40684 47406 40686 47458
rect 40738 47406 40740 47458
rect 40684 47124 40740 47406
rect 40684 47058 40740 47068
rect 40684 46900 40740 46910
rect 40572 46844 40684 46900
rect 40460 46834 40516 46844
rect 40684 46806 40740 46844
rect 40796 46788 40852 48190
rect 40236 46622 40238 46674
rect 40290 46622 40292 46674
rect 40236 46610 40292 46622
rect 40348 46674 40404 46686
rect 40348 46622 40350 46674
rect 40402 46622 40404 46674
rect 40348 46564 40404 46622
rect 40572 46676 40628 46686
rect 40572 46582 40628 46620
rect 40348 46498 40404 46508
rect 40012 45726 40014 45778
rect 40066 45726 40068 45778
rect 39564 45108 39620 45118
rect 39564 45014 39620 45052
rect 39676 44548 39732 44558
rect 39564 43764 39620 43774
rect 39452 43762 39620 43764
rect 39452 43710 39566 43762
rect 39618 43710 39620 43762
rect 39452 43708 39620 43710
rect 39564 43698 39620 43708
rect 39676 43764 39732 44492
rect 39900 44100 39956 44110
rect 39340 43362 39396 43372
rect 39452 43316 39508 43326
rect 39452 42978 39508 43260
rect 39676 42980 39732 43708
rect 39452 42926 39454 42978
rect 39506 42926 39508 42978
rect 39452 42914 39508 42926
rect 39564 42924 39732 42980
rect 39788 44098 39956 44100
rect 39788 44046 39902 44098
rect 39954 44046 39956 44098
rect 39788 44044 39956 44046
rect 39452 42756 39508 42766
rect 39340 42644 39396 42654
rect 39340 42082 39396 42588
rect 39340 42030 39342 42082
rect 39394 42030 39396 42082
rect 39340 42018 39396 42030
rect 39228 41694 39230 41746
rect 39282 41694 39284 41746
rect 39228 41682 39284 41694
rect 39116 41246 39118 41298
rect 39170 41246 39172 41298
rect 39116 41234 39172 41246
rect 38892 41056 38948 41132
rect 39116 41076 39172 41086
rect 39116 40982 39172 41020
rect 38332 40964 38388 40974
rect 38220 40516 38276 40526
rect 38220 40422 38276 40460
rect 38332 40402 38388 40908
rect 39116 40628 39172 40638
rect 39116 40534 39172 40572
rect 38332 40350 38334 40402
rect 38386 40350 38388 40402
rect 38332 40068 38388 40350
rect 38668 40404 38724 40414
rect 38668 40402 38836 40404
rect 38668 40350 38670 40402
rect 38722 40350 38836 40402
rect 38668 40348 38836 40350
rect 38668 40338 38724 40348
rect 38108 39566 38110 39618
rect 38162 39566 38164 39618
rect 38108 39554 38164 39566
rect 38220 40012 38388 40068
rect 37996 38782 37998 38834
rect 38050 38782 38052 38834
rect 37996 38668 38052 38782
rect 38220 38834 38276 40012
rect 38332 39844 38388 39854
rect 38332 39060 38388 39788
rect 38668 39732 38724 39742
rect 38780 39732 38836 40348
rect 39340 39956 39396 39966
rect 39004 39732 39060 39742
rect 38780 39676 39004 39732
rect 38668 39638 38724 39676
rect 39004 39618 39060 39676
rect 39340 39730 39396 39900
rect 39340 39678 39342 39730
rect 39394 39678 39396 39730
rect 39340 39666 39396 39678
rect 39004 39566 39006 39618
rect 39058 39566 39060 39618
rect 39004 39554 39060 39566
rect 38556 39508 38612 39518
rect 38332 38994 38388 39004
rect 38444 39396 38500 39406
rect 38444 38946 38500 39340
rect 38444 38894 38446 38946
rect 38498 38894 38500 38946
rect 38444 38882 38500 38894
rect 38220 38782 38222 38834
rect 38274 38782 38276 38834
rect 38220 38770 38276 38782
rect 37884 38612 38052 38668
rect 38332 38722 38388 38734
rect 38556 38724 38612 39452
rect 39004 39284 39060 39294
rect 39004 38834 39060 39228
rect 39452 39060 39508 42700
rect 39564 40964 39620 42924
rect 39788 42868 39844 44044
rect 39900 44034 39956 44044
rect 40012 43876 40068 45726
rect 40348 46116 40404 46126
rect 40348 45778 40404 46060
rect 40796 46116 40852 46732
rect 40908 48244 40964 48254
rect 40908 47684 40964 48188
rect 41132 47684 41188 50540
rect 41244 48802 41300 48814
rect 41244 48750 41246 48802
rect 41298 48750 41300 48802
rect 41244 48244 41300 48750
rect 41244 48178 41300 48188
rect 41132 47628 41300 47684
rect 40908 47458 40964 47628
rect 40908 47406 40910 47458
rect 40962 47406 40964 47458
rect 40908 46564 40964 47406
rect 41132 47458 41188 47470
rect 41132 47406 41134 47458
rect 41186 47406 41188 47458
rect 41020 47346 41076 47358
rect 41020 47294 41022 47346
rect 41074 47294 41076 47346
rect 41020 47012 41076 47294
rect 41020 46946 41076 46956
rect 41132 46676 41188 47406
rect 41132 46610 41188 46620
rect 40908 46498 40964 46508
rect 40796 46050 40852 46060
rect 40348 45726 40350 45778
rect 40402 45726 40404 45778
rect 40348 45714 40404 45726
rect 40460 45892 40516 45902
rect 41244 45892 41300 47628
rect 40460 45106 40516 45836
rect 40460 45054 40462 45106
rect 40514 45054 40516 45106
rect 40460 45042 40516 45054
rect 40572 45836 41300 45892
rect 40236 44548 40292 44558
rect 40236 44434 40292 44492
rect 40236 44382 40238 44434
rect 40290 44382 40292 44434
rect 40236 44370 40292 44382
rect 39900 43820 40068 43876
rect 39900 42980 39956 43820
rect 40236 43652 40292 43662
rect 40124 43650 40292 43652
rect 40124 43598 40238 43650
rect 40290 43598 40292 43650
rect 40124 43596 40292 43598
rect 39900 42914 39956 42924
rect 40012 43538 40068 43550
rect 40012 43486 40014 43538
rect 40066 43486 40068 43538
rect 39788 42802 39844 42812
rect 40012 42866 40068 43486
rect 40012 42814 40014 42866
rect 40066 42814 40068 42866
rect 40012 42802 40068 42814
rect 39676 42756 39732 42766
rect 39676 42662 39732 42700
rect 40012 42642 40068 42654
rect 40012 42590 40014 42642
rect 40066 42590 40068 42642
rect 40012 42308 40068 42590
rect 39900 41972 39956 41982
rect 39900 41878 39956 41916
rect 40012 41300 40068 42252
rect 40124 42196 40180 43596
rect 40236 43586 40292 43596
rect 40348 43650 40404 43662
rect 40348 43598 40350 43650
rect 40402 43598 40404 43650
rect 40236 43428 40292 43438
rect 40236 43334 40292 43372
rect 40236 42980 40292 42990
rect 40236 42886 40292 42924
rect 40236 42196 40292 42206
rect 40124 42194 40292 42196
rect 40124 42142 40238 42194
rect 40290 42142 40292 42194
rect 40124 42140 40292 42142
rect 40236 42130 40292 42140
rect 39900 41244 40068 41300
rect 40124 41970 40180 41982
rect 40124 41918 40126 41970
rect 40178 41918 40180 41970
rect 39676 41076 39732 41086
rect 39676 40982 39732 41020
rect 39564 40898 39620 40908
rect 39900 40740 39956 41244
rect 40012 41074 40068 41086
rect 40012 41022 40014 41074
rect 40066 41022 40068 41074
rect 40012 40964 40068 41022
rect 40124 41076 40180 41918
rect 40348 41972 40404 43598
rect 40460 42868 40516 42878
rect 40460 42082 40516 42812
rect 40460 42030 40462 42082
rect 40514 42030 40516 42082
rect 40460 42018 40516 42030
rect 40348 41906 40404 41916
rect 40572 41860 40628 45836
rect 40796 45668 40852 45678
rect 40684 45666 40852 45668
rect 40684 45614 40798 45666
rect 40850 45614 40852 45666
rect 40684 45612 40852 45614
rect 40684 45218 40740 45612
rect 40796 45602 40852 45612
rect 41244 45666 41300 45678
rect 41244 45614 41246 45666
rect 41298 45614 41300 45666
rect 40684 45166 40686 45218
rect 40738 45166 40740 45218
rect 40684 44884 40740 45166
rect 41132 45108 41188 45118
rect 40684 44818 40740 44828
rect 40908 44996 40964 45006
rect 40684 44100 40740 44110
rect 40684 43316 40740 44044
rect 40796 43540 40852 43550
rect 40796 43446 40852 43484
rect 40684 43250 40740 43260
rect 40684 42756 40740 42766
rect 40684 42662 40740 42700
rect 40460 41804 40628 41860
rect 40684 42084 40740 42094
rect 40124 41010 40180 41020
rect 40236 41524 40292 41534
rect 40012 40898 40068 40908
rect 39564 40684 39956 40740
rect 39564 40626 39620 40684
rect 39564 40574 39566 40626
rect 39618 40574 39620 40626
rect 39564 40562 39620 40574
rect 39564 39060 39620 39070
rect 39452 39058 39620 39060
rect 39452 39006 39566 39058
rect 39618 39006 39620 39058
rect 39452 39004 39620 39006
rect 39564 38994 39620 39004
rect 39004 38782 39006 38834
rect 39058 38782 39060 38834
rect 39004 38770 39060 38782
rect 38332 38670 38334 38722
rect 38386 38670 38388 38722
rect 37772 38052 37828 38062
rect 37772 37958 37828 37996
rect 37212 37874 37268 37884
rect 37548 37938 37716 37940
rect 37548 37886 37662 37938
rect 37714 37886 37716 37938
rect 37548 37884 37716 37886
rect 36876 37828 36932 37838
rect 36876 37490 36932 37772
rect 36876 37438 36878 37490
rect 36930 37438 36932 37490
rect 36876 37426 36932 37438
rect 36988 37716 37044 37726
rect 36988 37490 37044 37660
rect 36988 37438 36990 37490
rect 37042 37438 37044 37490
rect 36988 37426 37044 37438
rect 36764 37266 36820 37278
rect 36764 37214 36766 37266
rect 36818 37214 36820 37266
rect 36764 37044 36820 37214
rect 37436 37268 37492 37278
rect 37548 37268 37604 37884
rect 37660 37874 37716 37884
rect 37436 37266 37604 37268
rect 37436 37214 37438 37266
rect 37490 37214 37604 37266
rect 37436 37212 37604 37214
rect 37436 37202 37492 37212
rect 36764 36978 36820 36988
rect 37660 37042 37716 37054
rect 37660 36990 37662 37042
rect 37714 36990 37716 37042
rect 36988 36820 37044 36830
rect 36988 35924 37044 36764
rect 37436 36820 37492 36830
rect 37436 36594 37492 36764
rect 37436 36542 37438 36594
rect 37490 36542 37492 36594
rect 37436 36530 37492 36542
rect 36988 35792 37044 35868
rect 37436 35812 37492 35822
rect 37436 35718 37492 35756
rect 37100 35700 37156 35710
rect 36988 34692 37044 34702
rect 36764 33908 36820 33918
rect 36764 33458 36820 33852
rect 36764 33406 36766 33458
rect 36818 33406 36820 33458
rect 36764 33394 36820 33406
rect 36876 33124 36932 33134
rect 36876 32674 36932 33068
rect 36876 32622 36878 32674
rect 36930 32622 36932 32674
rect 36876 32610 36932 32622
rect 36988 32116 37044 34636
rect 36988 32050 37044 32060
rect 36652 31838 36654 31890
rect 36706 31838 36708 31890
rect 36652 31826 36708 31838
rect 36988 31892 37044 31902
rect 36316 31724 36484 31780
rect 36316 31556 36372 31566
rect 36316 31462 36372 31500
rect 36428 29652 36484 31724
rect 36540 31554 36596 31566
rect 36540 31502 36542 31554
rect 36594 31502 36596 31554
rect 36540 31444 36596 31502
rect 36540 31378 36596 31388
rect 36764 31554 36820 31566
rect 36764 31502 36766 31554
rect 36818 31502 36820 31554
rect 36540 31106 36596 31118
rect 36540 31054 36542 31106
rect 36594 31054 36596 31106
rect 36540 29876 36596 31054
rect 36540 29810 36596 29820
rect 36764 29652 36820 31502
rect 36428 29596 36596 29652
rect 36316 29426 36372 29438
rect 36316 29374 36318 29426
rect 36370 29374 36372 29426
rect 36316 28644 36372 29374
rect 36428 28644 36484 28654
rect 36316 28642 36484 28644
rect 36316 28590 36430 28642
rect 36482 28590 36484 28642
rect 36316 28588 36484 28590
rect 36428 28578 36484 28588
rect 36540 28644 36596 29596
rect 36764 29586 36820 29596
rect 36876 29426 36932 29438
rect 36876 29374 36878 29426
rect 36930 29374 36932 29426
rect 36540 28578 36596 28588
rect 36764 28756 36820 28766
rect 36764 28530 36820 28700
rect 36764 28478 36766 28530
rect 36818 28478 36820 28530
rect 36764 28466 36820 28478
rect 36652 28420 36708 28430
rect 36204 27570 36260 27580
rect 36540 28418 36708 28420
rect 36540 28366 36654 28418
rect 36706 28366 36708 28418
rect 36540 28364 36708 28366
rect 36092 27134 36094 27186
rect 36146 27134 36148 27186
rect 36092 27122 36148 27134
rect 36540 27188 36596 28364
rect 36652 28354 36708 28364
rect 36652 27970 36708 27982
rect 36652 27918 36654 27970
rect 36706 27918 36708 27970
rect 36652 27300 36708 27918
rect 36764 27860 36820 27870
rect 36764 27766 36820 27804
rect 36876 27746 36932 29374
rect 36988 29314 37044 31836
rect 36988 29262 36990 29314
rect 37042 29262 37044 29314
rect 36988 29250 37044 29262
rect 36876 27694 36878 27746
rect 36930 27694 36932 27746
rect 36876 27682 36932 27694
rect 36988 29092 37044 29102
rect 36652 27234 36708 27244
rect 36764 27636 36820 27646
rect 36540 27122 36596 27132
rect 36540 26964 36596 26974
rect 36540 26852 36596 26908
rect 36540 26850 36708 26852
rect 36540 26798 36542 26850
rect 36594 26798 36708 26850
rect 36540 26796 36708 26798
rect 36540 26786 36596 26796
rect 35980 26562 36036 26572
rect 36540 26628 36596 26638
rect 35868 26462 35870 26514
rect 35922 26462 35924 26514
rect 35868 26450 35924 26462
rect 36092 26292 36148 26302
rect 36428 26292 36484 26302
rect 36092 26290 36372 26292
rect 36092 26238 36094 26290
rect 36146 26238 36372 26290
rect 36092 26236 36372 26238
rect 36092 26226 36148 26236
rect 35756 26012 36148 26068
rect 35868 25732 35924 25742
rect 35868 25506 35924 25676
rect 35868 25454 35870 25506
rect 35922 25454 35924 25506
rect 35868 25442 35924 25454
rect 35532 25394 35700 25396
rect 35532 25342 35534 25394
rect 35586 25342 35700 25394
rect 35532 25340 35700 25342
rect 35532 25330 35588 25340
rect 35756 25282 35812 25294
rect 35756 25230 35758 25282
rect 35810 25230 35812 25282
rect 35644 24724 35700 24734
rect 34300 22206 34302 22258
rect 34354 22206 34356 22258
rect 34188 21252 34244 21262
rect 33852 20802 34132 20804
rect 33852 20750 33854 20802
rect 33906 20750 34132 20802
rect 33852 20748 34132 20750
rect 33852 20738 33908 20748
rect 34076 20130 34132 20748
rect 34188 20580 34244 21196
rect 34300 21026 34356 22206
rect 34748 22316 34916 22372
rect 34972 24556 35252 24612
rect 35532 24612 35588 24622
rect 34972 22372 35028 24556
rect 35532 24518 35588 24556
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35644 23826 35700 24668
rect 35644 23774 35646 23826
rect 35698 23774 35700 23826
rect 35644 23762 35700 23774
rect 35308 23714 35364 23726
rect 35308 23662 35310 23714
rect 35362 23662 35364 23714
rect 35084 23154 35140 23166
rect 35084 23102 35086 23154
rect 35138 23102 35140 23154
rect 35084 22596 35140 23102
rect 35308 23156 35364 23662
rect 35756 23380 35812 25230
rect 35980 24836 36036 24846
rect 35980 24742 36036 24780
rect 35756 23314 35812 23324
rect 35980 24498 36036 24510
rect 35980 24446 35982 24498
rect 36034 24446 36036 24498
rect 35868 23156 35924 23166
rect 35308 23154 35924 23156
rect 35308 23102 35870 23154
rect 35922 23102 35924 23154
rect 35308 23100 35924 23102
rect 35532 22932 35588 22942
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22540 35476 22596
rect 34972 22316 35140 22372
rect 34300 20974 34302 21026
rect 34354 20974 34356 21026
rect 34300 20962 34356 20974
rect 34412 22146 34468 22158
rect 34412 22094 34414 22146
rect 34466 22094 34468 22146
rect 34412 21588 34468 22094
rect 34412 20916 34468 21532
rect 34412 20850 34468 20860
rect 34524 21924 34580 21934
rect 34524 21586 34580 21868
rect 34524 21534 34526 21586
rect 34578 21534 34580 21586
rect 34300 20580 34356 20590
rect 34188 20578 34468 20580
rect 34188 20526 34302 20578
rect 34354 20526 34468 20578
rect 34188 20524 34468 20526
rect 34300 20514 34356 20524
rect 34076 20078 34078 20130
rect 34130 20078 34132 20130
rect 33852 20018 33908 20030
rect 33852 19966 33854 20018
rect 33906 19966 33908 20018
rect 33852 19796 33908 19966
rect 33852 19730 33908 19740
rect 33852 19348 33908 19358
rect 34076 19348 34132 20078
rect 34300 19348 34356 19358
rect 33852 19346 34356 19348
rect 33852 19294 33854 19346
rect 33906 19294 34302 19346
rect 34354 19294 34356 19346
rect 33852 19292 34356 19294
rect 33852 19282 33908 19292
rect 34300 19282 34356 19292
rect 33740 19068 34132 19124
rect 33740 18228 33796 18238
rect 33964 18228 34020 18238
rect 33740 17780 33796 18172
rect 33740 17714 33796 17724
rect 33852 18226 34020 18228
rect 33852 18174 33966 18226
rect 34018 18174 34020 18226
rect 33852 18172 34020 18174
rect 33516 17614 33518 17666
rect 33570 17614 33572 17666
rect 33516 16884 33572 17614
rect 33516 16818 33572 16828
rect 33852 17556 33908 18172
rect 33964 18162 34020 18172
rect 33964 17780 34020 17790
rect 33964 17686 34020 17724
rect 33516 16660 33572 16670
rect 33516 16210 33572 16604
rect 33628 16324 33684 16334
rect 33852 16324 33908 17500
rect 33964 17108 34020 17118
rect 33964 17014 34020 17052
rect 34076 16884 34132 19068
rect 34300 18674 34356 18686
rect 34300 18622 34302 18674
rect 34354 18622 34356 18674
rect 34300 18452 34356 18622
rect 34300 18386 34356 18396
rect 34412 18340 34468 20524
rect 34412 18274 34468 18284
rect 34524 20020 34580 21534
rect 34188 18226 34244 18238
rect 34188 18174 34190 18226
rect 34242 18174 34244 18226
rect 34188 17892 34244 18174
rect 34300 18228 34356 18238
rect 34300 18134 34356 18172
rect 34188 17826 34244 17836
rect 34412 16996 34468 17006
rect 34412 16902 34468 16940
rect 33628 16322 33908 16324
rect 33628 16270 33630 16322
rect 33682 16270 33908 16322
rect 33628 16268 33908 16270
rect 33628 16258 33684 16268
rect 33516 16158 33518 16210
rect 33570 16158 33572 16210
rect 33516 16146 33572 16158
rect 33740 15540 33796 15550
rect 33740 15446 33796 15484
rect 33852 15426 33908 16268
rect 33852 15374 33854 15426
rect 33906 15374 33908 15426
rect 33852 15362 33908 15374
rect 33964 16828 34132 16884
rect 33516 15316 33572 15326
rect 33516 15222 33572 15260
rect 33404 8082 33460 8092
rect 33516 14308 33572 14318
rect 33516 5796 33572 14252
rect 33628 13972 33684 13982
rect 33628 13878 33684 13916
rect 33964 13860 34020 16828
rect 34524 16436 34580 19964
rect 34748 19796 34804 22316
rect 34972 22146 35028 22158
rect 34972 22094 34974 22146
rect 35026 22094 35028 22146
rect 34972 22036 35028 22094
rect 34972 21970 35028 21980
rect 34860 21026 34916 21038
rect 34860 20974 34862 21026
rect 34914 20974 34916 21026
rect 34860 20914 34916 20974
rect 34860 20862 34862 20914
rect 34914 20862 34916 20914
rect 34860 20850 34916 20862
rect 34860 20356 34916 20366
rect 34860 20132 34916 20300
rect 34860 20130 35028 20132
rect 34860 20078 34862 20130
rect 34914 20078 35028 20130
rect 34860 20076 35028 20078
rect 34860 20066 34916 20076
rect 34748 19730 34804 19740
rect 34748 19236 34804 19246
rect 34748 19142 34804 19180
rect 34860 19124 34916 19134
rect 34860 19030 34916 19068
rect 34860 18340 34916 18350
rect 34972 18340 35028 20076
rect 35084 19348 35140 22316
rect 35420 21810 35476 22540
rect 35420 21758 35422 21810
rect 35474 21758 35476 21810
rect 35420 21746 35476 21758
rect 35420 21586 35476 21598
rect 35420 21534 35422 21586
rect 35474 21534 35476 21586
rect 35420 21476 35476 21534
rect 35420 21410 35476 21420
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35420 21028 35476 21038
rect 35308 20578 35364 20590
rect 35308 20526 35310 20578
rect 35362 20526 35364 20578
rect 35308 20468 35364 20526
rect 35308 20402 35364 20412
rect 35196 20356 35252 20366
rect 35196 20130 35252 20300
rect 35196 20078 35198 20130
rect 35250 20078 35252 20130
rect 35196 20066 35252 20078
rect 35420 19796 35476 20972
rect 35532 20468 35588 22876
rect 35756 22596 35812 23100
rect 35868 23090 35924 23100
rect 35756 22502 35812 22540
rect 35868 22370 35924 22382
rect 35868 22318 35870 22370
rect 35922 22318 35924 22370
rect 35644 22148 35700 22158
rect 35644 20804 35700 22092
rect 35756 21364 35812 21374
rect 35756 21270 35812 21308
rect 35868 21028 35924 22318
rect 35980 21812 36036 24446
rect 36092 23380 36148 26012
rect 36204 25844 36260 25854
rect 36204 25508 36260 25788
rect 36316 25508 36372 26236
rect 36428 26198 36484 26236
rect 36428 25508 36484 25518
rect 36316 25452 36428 25508
rect 36204 24050 36260 25452
rect 36428 25376 36484 25452
rect 36428 24612 36484 24622
rect 36540 24612 36596 26572
rect 36652 26180 36708 26796
rect 36764 26404 36820 27580
rect 36764 26338 36820 26348
rect 36876 26180 36932 26190
rect 36652 26178 36932 26180
rect 36652 26126 36878 26178
rect 36930 26126 36932 26178
rect 36652 26124 36932 26126
rect 36652 25620 36708 25630
rect 36652 25394 36708 25564
rect 36652 25342 36654 25394
rect 36706 25342 36708 25394
rect 36652 25330 36708 25342
rect 36764 25394 36820 25406
rect 36764 25342 36766 25394
rect 36818 25342 36820 25394
rect 36428 24610 36596 24612
rect 36428 24558 36430 24610
rect 36482 24558 36596 24610
rect 36428 24556 36596 24558
rect 36652 25172 36708 25182
rect 36428 24498 36484 24556
rect 36428 24446 36430 24498
rect 36482 24446 36484 24498
rect 36428 24434 36484 24446
rect 36204 23998 36206 24050
rect 36258 23998 36260 24050
rect 36204 23986 36260 23998
rect 36540 23716 36596 23726
rect 36540 23622 36596 23660
rect 36428 23604 36484 23614
rect 36316 23492 36372 23502
rect 36204 23380 36260 23390
rect 36092 23378 36260 23380
rect 36092 23326 36206 23378
rect 36258 23326 36260 23378
rect 36092 23324 36260 23326
rect 36204 23314 36260 23324
rect 36316 23378 36372 23436
rect 36316 23326 36318 23378
rect 36370 23326 36372 23378
rect 36316 23314 36372 23326
rect 36092 23156 36148 23166
rect 36092 23062 36148 23100
rect 36428 22596 36484 23548
rect 35980 21746 36036 21756
rect 36092 22540 36484 22596
rect 36540 23154 36596 23166
rect 36540 23102 36542 23154
rect 36594 23102 36596 23154
rect 35868 20962 35924 20972
rect 35980 21588 36036 21598
rect 35868 20804 35924 20814
rect 35644 20802 35924 20804
rect 35644 20750 35870 20802
rect 35922 20750 35924 20802
rect 35644 20748 35924 20750
rect 35868 20738 35924 20748
rect 35980 20580 36036 21532
rect 35532 20402 35588 20412
rect 35756 20524 36036 20580
rect 35756 20356 35812 20524
rect 36092 20356 36148 22540
rect 36428 22372 36484 22382
rect 36316 22316 36428 22372
rect 36204 22148 36260 22158
rect 36204 22054 36260 22092
rect 36204 21700 36260 21710
rect 36316 21700 36372 22316
rect 36428 22278 36484 22316
rect 36540 22370 36596 23102
rect 36540 22318 36542 22370
rect 36594 22318 36596 22370
rect 36540 22306 36596 22318
rect 36652 22260 36708 25116
rect 36764 22932 36820 25342
rect 36764 22866 36820 22876
rect 36876 22820 36932 26124
rect 36988 25620 37044 29036
rect 37100 26628 37156 35644
rect 37436 35588 37492 35598
rect 37212 34130 37268 34142
rect 37212 34078 37214 34130
rect 37266 34078 37268 34130
rect 37212 29764 37268 34078
rect 37436 34020 37492 35532
rect 37548 34804 37604 34814
rect 37548 34690 37604 34748
rect 37548 34638 37550 34690
rect 37602 34638 37604 34690
rect 37548 34580 37604 34638
rect 37548 34514 37604 34524
rect 37548 34020 37604 34030
rect 37436 34018 37604 34020
rect 37436 33966 37550 34018
rect 37602 33966 37604 34018
rect 37436 33964 37604 33966
rect 37436 33572 37492 33582
rect 37548 33572 37604 33964
rect 37436 33570 37604 33572
rect 37436 33518 37438 33570
rect 37490 33518 37604 33570
rect 37436 33516 37604 33518
rect 37436 33458 37492 33516
rect 37436 33406 37438 33458
rect 37490 33406 37492 33458
rect 37436 33394 37492 33406
rect 37548 33012 37604 33022
rect 37436 32676 37492 32686
rect 37436 32562 37492 32620
rect 37548 32674 37604 32956
rect 37548 32622 37550 32674
rect 37602 32622 37604 32674
rect 37548 32610 37604 32622
rect 37436 32510 37438 32562
rect 37490 32510 37492 32562
rect 37436 32498 37492 32510
rect 37660 32340 37716 36990
rect 37884 36036 37940 38612
rect 38332 38052 38388 38670
rect 38332 37986 38388 37996
rect 38444 38668 38556 38724
rect 38332 37828 38388 37838
rect 38332 37490 38388 37772
rect 38332 37438 38334 37490
rect 38386 37438 38388 37490
rect 38332 37426 38388 37438
rect 38444 37826 38500 38668
rect 38556 38658 38612 38668
rect 39228 38724 39284 38762
rect 39676 38668 39732 40684
rect 40012 40290 40068 40302
rect 40012 40238 40014 40290
rect 40066 40238 40068 40290
rect 40012 39508 40068 40238
rect 40012 39442 40068 39452
rect 39900 39396 39956 39406
rect 39900 39302 39956 39340
rect 40236 39284 40292 41468
rect 40460 40626 40516 41804
rect 40572 41300 40628 41310
rect 40684 41300 40740 42028
rect 40572 41298 40740 41300
rect 40572 41246 40574 41298
rect 40626 41246 40740 41298
rect 40572 41244 40740 41246
rect 40572 41234 40628 41244
rect 40460 40574 40462 40626
rect 40514 40574 40516 40626
rect 40460 39732 40516 40574
rect 40460 39666 40516 39676
rect 40908 39620 40964 44940
rect 41132 44434 41188 45052
rect 41132 44382 41134 44434
rect 41186 44382 41188 44434
rect 41132 44370 41188 44382
rect 41244 44772 41300 45614
rect 41244 43764 41300 44716
rect 41244 43698 41300 43708
rect 41132 43652 41188 43662
rect 41020 43428 41076 43438
rect 41020 41300 41076 43372
rect 41132 42532 41188 43596
rect 41356 42756 41412 50540
rect 42028 50482 42084 50494
rect 42028 50430 42030 50482
rect 42082 50430 42084 50482
rect 41580 50372 41636 50382
rect 41468 50370 41636 50372
rect 41468 50318 41582 50370
rect 41634 50318 41636 50370
rect 41468 50316 41636 50318
rect 41468 49698 41524 50316
rect 41580 50306 41636 50316
rect 41468 49646 41470 49698
rect 41522 49646 41524 49698
rect 41468 49140 41524 49646
rect 41468 49084 41860 49140
rect 41692 48916 41748 48926
rect 41692 48822 41748 48860
rect 41692 48244 41748 48254
rect 41580 48130 41636 48142
rect 41580 48078 41582 48130
rect 41634 48078 41636 48130
rect 41580 47908 41636 48078
rect 41468 46564 41524 46574
rect 41468 46470 41524 46508
rect 41468 44994 41524 45006
rect 41468 44942 41470 44994
rect 41522 44942 41524 44994
rect 41468 43652 41524 44942
rect 41580 44436 41636 47852
rect 41692 47570 41748 48188
rect 41804 48132 41860 49084
rect 41916 48132 41972 48142
rect 41804 48130 41972 48132
rect 41804 48078 41918 48130
rect 41970 48078 41972 48130
rect 41804 48076 41972 48078
rect 41692 47518 41694 47570
rect 41746 47518 41748 47570
rect 41692 47460 41748 47518
rect 41692 47394 41748 47404
rect 41804 47124 41860 47134
rect 41692 46564 41748 46574
rect 41692 46002 41748 46508
rect 41692 45950 41694 46002
rect 41746 45950 41748 46002
rect 41692 45892 41748 45950
rect 41692 45826 41748 45836
rect 41804 45108 41860 47068
rect 41916 47012 41972 48076
rect 42028 47684 42084 50430
rect 42140 47796 42196 52220
rect 42476 52274 42532 53116
rect 42700 54292 42756 54302
rect 42700 53172 42756 54236
rect 42812 53844 42868 53854
rect 42812 53750 42868 53788
rect 42924 53732 42980 54460
rect 43260 54422 43316 54460
rect 43708 54514 43764 54572
rect 43708 54462 43710 54514
rect 43762 54462 43764 54514
rect 42924 53506 42980 53676
rect 43148 54404 43204 54414
rect 43148 53732 43204 54348
rect 43484 53732 43540 53742
rect 43708 53732 43764 54462
rect 43820 54514 43876 54526
rect 43820 54462 43822 54514
rect 43874 54462 43876 54514
rect 43820 54404 43876 54462
rect 43820 54338 43876 54348
rect 43932 54514 43988 54526
rect 43932 54462 43934 54514
rect 43986 54462 43988 54514
rect 43148 53730 43316 53732
rect 43148 53678 43150 53730
rect 43202 53678 43316 53730
rect 43148 53676 43316 53678
rect 43148 53666 43204 53676
rect 42924 53454 42926 53506
rect 42978 53454 42980 53506
rect 42924 53284 42980 53454
rect 42924 53228 43204 53284
rect 42812 53172 42868 53182
rect 42700 53170 42868 53172
rect 42700 53118 42814 53170
rect 42866 53118 42868 53170
rect 42700 53116 42868 53118
rect 42588 53058 42644 53116
rect 42812 53106 42868 53116
rect 42588 53006 42590 53058
rect 42642 53006 42644 53058
rect 42588 52994 42644 53006
rect 43036 53058 43092 53070
rect 43036 53006 43038 53058
rect 43090 53006 43092 53058
rect 42700 52836 42756 52846
rect 42700 52742 42756 52780
rect 42812 52388 42868 52398
rect 42812 52294 42868 52332
rect 43036 52388 43092 53006
rect 43036 52322 43092 52332
rect 42476 52222 42478 52274
rect 42530 52222 42532 52274
rect 42476 52210 42532 52222
rect 42252 52164 42308 52174
rect 42252 52070 42308 52108
rect 42588 52050 42644 52062
rect 42588 51998 42590 52050
rect 42642 51998 42644 52050
rect 42588 51940 42644 51998
rect 42588 51874 42644 51884
rect 43148 51602 43204 53228
rect 43260 52386 43316 53676
rect 43484 53730 43764 53732
rect 43484 53678 43486 53730
rect 43538 53678 43764 53730
rect 43484 53676 43764 53678
rect 43484 53666 43540 53676
rect 43596 53508 43652 53518
rect 43260 52334 43262 52386
rect 43314 52334 43316 52386
rect 43260 52322 43316 52334
rect 43372 53284 43428 53294
rect 43148 51550 43150 51602
rect 43202 51550 43204 51602
rect 43148 51538 43204 51550
rect 43260 51604 43316 51614
rect 43372 51604 43428 53228
rect 43596 53058 43652 53452
rect 43596 53006 43598 53058
rect 43650 53006 43652 53058
rect 43596 52276 43652 53006
rect 43708 52722 43764 53676
rect 43932 53732 43988 54462
rect 43932 53666 43988 53676
rect 43932 53506 43988 53518
rect 43932 53454 43934 53506
rect 43986 53454 43988 53506
rect 43708 52670 43710 52722
rect 43762 52670 43764 52722
rect 43708 52658 43764 52670
rect 43820 53396 43876 53406
rect 43820 53058 43876 53340
rect 43932 53284 43988 53454
rect 44380 53508 44436 53518
rect 44380 53414 44436 53452
rect 45388 53508 45444 53518
rect 43932 53218 43988 53228
rect 43820 53006 43822 53058
rect 43874 53006 43876 53058
rect 43708 52276 43764 52286
rect 43596 52220 43708 52276
rect 43708 52144 43764 52220
rect 43316 51548 43428 51604
rect 43260 51378 43316 51548
rect 43260 51326 43262 51378
rect 43314 51326 43316 51378
rect 43820 51492 43876 53006
rect 44380 53172 44436 53182
rect 44380 52948 44436 53116
rect 43932 52946 44436 52948
rect 43932 52894 44382 52946
rect 44434 52894 44436 52946
rect 43932 52892 44436 52894
rect 43932 52386 43988 52892
rect 44380 52882 44436 52892
rect 45052 52834 45108 52846
rect 45052 52782 45054 52834
rect 45106 52782 45108 52834
rect 43932 52334 43934 52386
rect 43986 52334 43988 52386
rect 43932 52164 43988 52334
rect 44156 52722 44212 52734
rect 44156 52670 44158 52722
rect 44210 52670 44212 52722
rect 44156 52276 44212 52670
rect 44156 52182 44212 52220
rect 43932 52098 43988 52108
rect 43820 51360 43876 51436
rect 44380 52050 44436 52062
rect 44380 51998 44382 52050
rect 44434 51998 44436 52050
rect 44380 51380 44436 51998
rect 43260 51314 43316 51326
rect 44380 51314 44436 51324
rect 45052 51716 45108 52782
rect 45388 52274 45444 53452
rect 47068 53172 47124 53182
rect 47068 53078 47124 53116
rect 46844 52946 46900 52958
rect 46844 52894 46846 52946
rect 46898 52894 46900 52946
rect 46396 52834 46452 52846
rect 46396 52782 46398 52834
rect 46450 52782 46452 52834
rect 45948 52388 46004 52398
rect 45948 52294 46004 52332
rect 45388 52222 45390 52274
rect 45442 52222 45444 52274
rect 45388 52210 45444 52222
rect 46060 51940 46116 51950
rect 46060 51846 46116 51884
rect 46284 51938 46340 51950
rect 46284 51886 46286 51938
rect 46338 51886 46340 51938
rect 42252 51268 42308 51278
rect 42252 49922 42308 51212
rect 42700 51268 42756 51278
rect 42700 51266 42868 51268
rect 42700 51214 42702 51266
rect 42754 51214 42868 51266
rect 42700 51212 42868 51214
rect 42700 51202 42756 51212
rect 42700 51044 42756 51054
rect 42476 50932 42532 50942
rect 42476 50706 42532 50876
rect 42476 50654 42478 50706
rect 42530 50654 42532 50706
rect 42476 50642 42532 50654
rect 42700 50596 42756 50988
rect 42700 50502 42756 50540
rect 42588 50484 42644 50494
rect 42364 50482 42644 50484
rect 42364 50430 42590 50482
rect 42642 50430 42644 50482
rect 42364 50428 42644 50430
rect 42364 50034 42420 50428
rect 42588 50418 42644 50428
rect 42364 49982 42366 50034
rect 42418 49982 42420 50034
rect 42364 49970 42420 49982
rect 42252 49870 42254 49922
rect 42306 49870 42308 49922
rect 42252 49858 42308 49870
rect 42476 48914 42532 48926
rect 42476 48862 42478 48914
rect 42530 48862 42532 48914
rect 42476 48804 42532 48862
rect 42476 48738 42532 48748
rect 42812 48802 42868 51212
rect 44828 51266 44884 51278
rect 44828 51214 44830 51266
rect 44882 51214 44884 51266
rect 43484 51156 43540 51166
rect 43372 51154 43540 51156
rect 43372 51102 43486 51154
rect 43538 51102 43540 51154
rect 43372 51100 43540 51102
rect 43372 50820 43428 51100
rect 43484 51090 43540 51100
rect 44044 51154 44100 51166
rect 44044 51102 44046 51154
rect 44098 51102 44100 51154
rect 43372 50764 43652 50820
rect 43260 50484 43316 50494
rect 42812 48750 42814 48802
rect 42866 48750 42868 48802
rect 42364 48132 42420 48142
rect 42364 48038 42420 48076
rect 42700 48020 42756 48030
rect 42140 47740 42420 47796
rect 42028 47618 42084 47628
rect 42252 47236 42308 47246
rect 41916 46946 41972 46956
rect 42028 47234 42308 47236
rect 42028 47182 42254 47234
rect 42306 47182 42308 47234
rect 42028 47180 42308 47182
rect 41804 45042 41860 45052
rect 41916 44996 41972 45006
rect 42028 44996 42084 47180
rect 42252 47170 42308 47180
rect 42252 46562 42308 46574
rect 42252 46510 42254 46562
rect 42306 46510 42308 46562
rect 42252 46452 42308 46510
rect 42252 46386 42308 46396
rect 42252 45666 42308 45678
rect 42252 45614 42254 45666
rect 42306 45614 42308 45666
rect 41916 44994 42196 44996
rect 41916 44942 41918 44994
rect 41970 44942 42196 44994
rect 41916 44940 42196 44942
rect 41916 44930 41972 44940
rect 41580 44370 41636 44380
rect 41692 44100 41748 44110
rect 41692 44098 41860 44100
rect 41692 44046 41694 44098
rect 41746 44046 41860 44098
rect 41692 44044 41860 44046
rect 41692 44034 41748 44044
rect 41468 43586 41524 43596
rect 41692 43538 41748 43550
rect 41692 43486 41694 43538
rect 41746 43486 41748 43538
rect 41580 43316 41636 43326
rect 41356 42700 41524 42756
rect 41132 42438 41188 42476
rect 41244 42530 41300 42542
rect 41244 42478 41246 42530
rect 41298 42478 41300 42530
rect 41244 42196 41300 42478
rect 41356 42532 41412 42542
rect 41356 42438 41412 42476
rect 41244 42130 41300 42140
rect 41020 41206 41076 41244
rect 40908 39554 40964 39564
rect 39228 38658 39284 38668
rect 39340 38612 39732 38668
rect 40012 39228 40292 39284
rect 40348 39394 40404 39406
rect 40348 39342 40350 39394
rect 40402 39342 40404 39394
rect 39340 38050 39396 38612
rect 39340 37998 39342 38050
rect 39394 37998 39396 38050
rect 39340 37986 39396 37998
rect 39004 37940 39060 37950
rect 39004 37846 39060 37884
rect 38444 37774 38446 37826
rect 38498 37774 38500 37826
rect 37996 37156 38052 37166
rect 37996 37154 38164 37156
rect 37996 37102 37998 37154
rect 38050 37102 38164 37154
rect 37996 37100 38164 37102
rect 37996 37090 38052 37100
rect 37996 36372 38052 36382
rect 37996 36278 38052 36316
rect 37884 35980 38052 36036
rect 37772 35812 37828 35822
rect 37772 34914 37828 35756
rect 37772 34862 37774 34914
rect 37826 34862 37828 34914
rect 37772 34850 37828 34862
rect 37996 34354 38052 35980
rect 38108 35700 38164 37100
rect 38444 37042 38500 37774
rect 39564 37492 39620 37502
rect 39564 37398 39620 37436
rect 39900 37378 39956 37390
rect 39900 37326 39902 37378
rect 39954 37326 39956 37378
rect 39900 37268 39956 37326
rect 39900 37202 39956 37212
rect 38444 36990 38446 37042
rect 38498 36990 38500 37042
rect 38444 36978 38500 36990
rect 38780 37154 38836 37166
rect 38780 37102 38782 37154
rect 38834 37102 38836 37154
rect 38780 37044 38836 37102
rect 38780 36978 38836 36988
rect 39676 37156 39732 37166
rect 39004 36932 39060 36942
rect 38668 36708 38724 36718
rect 38668 36706 38948 36708
rect 38668 36654 38670 36706
rect 38722 36654 38948 36706
rect 38668 36652 38948 36654
rect 38668 36642 38724 36652
rect 38780 36484 38836 36494
rect 38220 36372 38276 36382
rect 38220 35812 38276 36316
rect 38780 36370 38836 36428
rect 38780 36318 38782 36370
rect 38834 36318 38836 36370
rect 38668 36260 38724 36270
rect 38668 36166 38724 36204
rect 38556 36036 38612 36046
rect 38556 35922 38612 35980
rect 38556 35870 38558 35922
rect 38610 35870 38612 35922
rect 38556 35858 38612 35870
rect 38220 35680 38276 35756
rect 38444 35700 38500 35710
rect 38108 35634 38164 35644
rect 38444 35606 38500 35644
rect 38668 35698 38724 35710
rect 38668 35646 38670 35698
rect 38722 35646 38724 35698
rect 38668 35588 38724 35646
rect 38556 34916 38612 34926
rect 38668 34916 38724 35532
rect 38556 34914 38724 34916
rect 38556 34862 38558 34914
rect 38610 34862 38724 34914
rect 38556 34860 38724 34862
rect 38556 34850 38612 34860
rect 38780 34692 38836 36318
rect 38892 35700 38948 36652
rect 38892 35606 38948 35644
rect 39004 35026 39060 36876
rect 39676 36484 39732 37100
rect 39676 36390 39732 36428
rect 39004 34974 39006 35026
rect 39058 34974 39060 35026
rect 39004 34962 39060 34974
rect 39116 36260 39172 36270
rect 37996 34302 37998 34354
rect 38050 34302 38052 34354
rect 37996 34290 38052 34302
rect 38668 34690 38836 34692
rect 38668 34638 38782 34690
rect 38834 34638 38836 34690
rect 38668 34636 38836 34638
rect 38108 34242 38164 34254
rect 38108 34190 38110 34242
rect 38162 34190 38164 34242
rect 37212 29698 37268 29708
rect 37324 32284 37716 32340
rect 37772 33684 37828 33694
rect 37324 29540 37380 32284
rect 37436 31780 37492 31790
rect 37436 31686 37492 31724
rect 37772 31668 37828 33628
rect 38108 33684 38164 34190
rect 38108 33618 38164 33628
rect 38444 34130 38500 34142
rect 38444 34078 38446 34130
rect 38498 34078 38500 34130
rect 37884 33570 37940 33582
rect 37884 33518 37886 33570
rect 37938 33518 37940 33570
rect 37884 33122 37940 33518
rect 38444 33572 38500 34078
rect 38444 33506 38500 33516
rect 37884 33070 37886 33122
rect 37938 33070 37940 33122
rect 37884 32900 37940 33070
rect 38444 33122 38500 33134
rect 38444 33070 38446 33122
rect 38498 33070 38500 33122
rect 37884 32844 38276 32900
rect 38108 32452 38164 32462
rect 37996 32396 38108 32452
rect 37884 31668 37940 31678
rect 37772 31666 37940 31668
rect 37772 31614 37886 31666
rect 37938 31614 37940 31666
rect 37772 31612 37940 31614
rect 37660 31556 37716 31566
rect 37660 31462 37716 31500
rect 37884 30994 37940 31612
rect 37996 31444 38052 32396
rect 38108 32358 38164 32396
rect 37996 31378 38052 31388
rect 38108 31668 38164 31678
rect 38220 31668 38276 32844
rect 38108 31666 38276 31668
rect 38108 31614 38110 31666
rect 38162 31614 38276 31666
rect 38108 31612 38276 31614
rect 38444 32676 38500 33070
rect 38556 33012 38612 33022
rect 38556 32786 38612 32956
rect 38556 32734 38558 32786
rect 38610 32734 38612 32786
rect 38556 32722 38612 32734
rect 38444 31780 38500 32620
rect 37884 30942 37886 30994
rect 37938 30942 37940 30994
rect 37884 30930 37940 30942
rect 37884 30100 37940 30110
rect 37884 30098 38052 30100
rect 37884 30046 37886 30098
rect 37938 30046 38052 30098
rect 37884 30044 38052 30046
rect 37884 30034 37940 30044
rect 37548 29988 37604 29998
rect 37548 29986 37716 29988
rect 37548 29934 37550 29986
rect 37602 29934 37716 29986
rect 37548 29932 37716 29934
rect 37548 29922 37604 29932
rect 37212 29484 37380 29540
rect 37212 27636 37268 29484
rect 37548 28756 37604 28766
rect 37548 28662 37604 28700
rect 37548 27970 37604 27982
rect 37548 27918 37550 27970
rect 37602 27918 37604 27970
rect 37212 27570 37268 27580
rect 37324 27858 37380 27870
rect 37324 27806 37326 27858
rect 37378 27806 37380 27858
rect 37324 27188 37380 27806
rect 37436 27860 37492 27870
rect 37436 27412 37492 27804
rect 37548 27748 37604 27918
rect 37660 27860 37716 29932
rect 37772 29652 37828 29662
rect 37772 28530 37828 29596
rect 37772 28478 37774 28530
rect 37826 28478 37828 28530
rect 37772 28466 37828 28478
rect 37884 29540 37940 29550
rect 37884 28084 37940 29484
rect 37996 29538 38052 30044
rect 38108 29988 38164 31612
rect 38444 30548 38500 31724
rect 38556 31892 38612 31902
rect 38556 31554 38612 31836
rect 38556 31502 38558 31554
rect 38610 31502 38612 31554
rect 38556 31332 38612 31502
rect 38668 31556 38724 34636
rect 38780 34626 38836 34636
rect 39004 34804 39060 34814
rect 39004 34690 39060 34748
rect 39004 34638 39006 34690
rect 39058 34638 39060 34690
rect 39004 34580 39060 34638
rect 39004 34514 39060 34524
rect 38892 34018 38948 34030
rect 38892 33966 38894 34018
rect 38946 33966 38948 34018
rect 38892 32564 38948 33966
rect 38892 32498 38948 32508
rect 39116 31892 39172 36204
rect 39340 36258 39396 36270
rect 39340 36206 39342 36258
rect 39394 36206 39396 36258
rect 39228 34916 39284 34926
rect 39228 34822 39284 34860
rect 39340 34580 39396 36206
rect 39564 35700 39620 35710
rect 39564 35606 39620 35644
rect 39900 35698 39956 35710
rect 39900 35646 39902 35698
rect 39954 35646 39956 35698
rect 39340 34514 39396 34524
rect 39788 35588 39844 35598
rect 39788 33346 39844 35532
rect 39900 35252 39956 35646
rect 39900 33908 39956 35196
rect 40012 34468 40068 39228
rect 40124 38722 40180 38734
rect 40124 38670 40126 38722
rect 40178 38670 40180 38722
rect 40124 37492 40180 38670
rect 40348 38668 40404 39342
rect 40796 39396 40852 39406
rect 41244 39396 41300 39406
rect 40796 39394 41300 39396
rect 40796 39342 40798 39394
rect 40850 39342 41246 39394
rect 41298 39342 41300 39394
rect 40796 39340 41300 39342
rect 40572 39284 40628 39294
rect 40572 39058 40628 39228
rect 40572 39006 40574 39058
rect 40626 39006 40628 39058
rect 40572 38994 40628 39006
rect 40796 38668 40852 39340
rect 41244 39330 41300 39340
rect 41468 38948 41524 42700
rect 41580 42532 41636 43260
rect 41692 43204 41748 43486
rect 41692 43138 41748 43148
rect 41804 42868 41860 44044
rect 41916 43764 41972 43774
rect 41972 43708 42084 43764
rect 41916 43670 41972 43708
rect 41804 42774 41860 42812
rect 41580 42466 41636 42476
rect 41804 41972 41860 41982
rect 41804 41970 41972 41972
rect 41804 41918 41806 41970
rect 41858 41918 41972 41970
rect 41804 41916 41972 41918
rect 41804 41906 41860 41916
rect 41692 41860 41748 41870
rect 41580 40964 41636 40974
rect 41580 40870 41636 40908
rect 41692 40626 41748 41804
rect 41916 41748 41972 41916
rect 42028 41970 42084 43708
rect 42140 43428 42196 44940
rect 42252 44100 42308 45614
rect 42364 45330 42420 47740
rect 42700 46562 42756 47964
rect 42812 47124 42868 48750
rect 42924 49698 42980 49710
rect 42924 49646 42926 49698
rect 42978 49646 42980 49698
rect 42924 48132 42980 49646
rect 43148 48468 43204 48478
rect 43260 48468 43316 50428
rect 43372 50482 43428 50764
rect 43372 50430 43374 50482
rect 43426 50430 43428 50482
rect 43372 50418 43428 50430
rect 43484 50594 43540 50606
rect 43484 50542 43486 50594
rect 43538 50542 43540 50594
rect 43484 50036 43540 50542
rect 43596 50484 43652 50764
rect 44044 50596 44100 51102
rect 44044 50530 44100 50540
rect 44716 50594 44772 50606
rect 44716 50542 44718 50594
rect 44770 50542 44772 50594
rect 44716 50484 44772 50542
rect 43596 50428 43764 50484
rect 43596 50036 43652 50046
rect 43484 49980 43596 50036
rect 43596 49942 43652 49980
rect 43148 48466 43316 48468
rect 43148 48414 43150 48466
rect 43202 48414 43316 48466
rect 43148 48412 43316 48414
rect 43372 49700 43428 49710
rect 43372 48914 43428 49644
rect 43708 49138 43764 50428
rect 44716 50418 44772 50428
rect 44156 49700 44212 49710
rect 44604 49700 44660 49710
rect 44156 49698 44548 49700
rect 44156 49646 44158 49698
rect 44210 49646 44548 49698
rect 44156 49644 44548 49646
rect 44156 49634 44212 49644
rect 43708 49086 43710 49138
rect 43762 49086 43764 49138
rect 43708 49074 43764 49086
rect 43932 49586 43988 49598
rect 43932 49534 43934 49586
rect 43986 49534 43988 49586
rect 43932 49476 43988 49534
rect 43932 49026 43988 49420
rect 43932 48974 43934 49026
rect 43986 48974 43988 49026
rect 43932 48962 43988 48974
rect 43372 48862 43374 48914
rect 43426 48862 43428 48914
rect 43148 48402 43204 48412
rect 42924 48066 42980 48076
rect 43372 48020 43428 48862
rect 43596 48802 43652 48814
rect 43596 48750 43598 48802
rect 43650 48750 43652 48802
rect 43596 48692 43652 48750
rect 43820 48804 43876 48814
rect 43820 48710 43876 48748
rect 44380 48804 44436 48814
rect 43596 48132 43652 48636
rect 43708 48132 43764 48142
rect 43596 48130 43876 48132
rect 43596 48078 43710 48130
rect 43762 48078 43876 48130
rect 43596 48076 43876 48078
rect 43708 48066 43764 48076
rect 43484 48020 43540 48030
rect 43372 48018 43540 48020
rect 43372 47966 43486 48018
rect 43538 47966 43540 48018
rect 43372 47964 43540 47966
rect 43036 47908 43092 47918
rect 42812 47058 42868 47068
rect 42924 47460 42980 47470
rect 42700 46510 42702 46562
rect 42754 46510 42756 46562
rect 42700 46498 42756 46510
rect 42924 46786 42980 47404
rect 43036 47458 43092 47852
rect 43036 47406 43038 47458
rect 43090 47406 43092 47458
rect 43036 46900 43092 47406
rect 43260 46900 43316 46910
rect 43036 46898 43316 46900
rect 43036 46846 43262 46898
rect 43314 46846 43316 46898
rect 43036 46844 43316 46846
rect 42924 46734 42926 46786
rect 42978 46734 42980 46786
rect 42924 46002 42980 46734
rect 43036 46676 43092 46686
rect 43036 46582 43092 46620
rect 43260 46564 43316 46844
rect 42924 45950 42926 46002
rect 42978 45950 42980 46002
rect 42924 45938 42980 45950
rect 43148 46508 43316 46564
rect 42364 45278 42366 45330
rect 42418 45278 42420 45330
rect 42364 45266 42420 45278
rect 42700 45106 42756 45118
rect 42700 45054 42702 45106
rect 42754 45054 42756 45106
rect 42700 44546 42756 45054
rect 42700 44494 42702 44546
rect 42754 44494 42756 44546
rect 42700 44482 42756 44494
rect 42924 44322 42980 44334
rect 42924 44270 42926 44322
rect 42978 44270 42980 44322
rect 42252 44034 42308 44044
rect 42364 44098 42420 44110
rect 42364 44046 42366 44098
rect 42418 44046 42420 44098
rect 42364 43876 42420 44046
rect 42364 43810 42420 43820
rect 42588 44098 42644 44110
rect 42588 44046 42590 44098
rect 42642 44046 42644 44098
rect 42140 43362 42196 43372
rect 42476 43538 42532 43550
rect 42476 43486 42478 43538
rect 42530 43486 42532 43538
rect 42476 43428 42532 43486
rect 42476 42084 42532 43372
rect 42588 42532 42644 44046
rect 42812 43764 42868 43774
rect 42812 43538 42868 43708
rect 42812 43486 42814 43538
rect 42866 43486 42868 43538
rect 42812 42756 42868 43486
rect 42924 43428 42980 44270
rect 43036 43428 43092 43438
rect 42924 43372 43036 43428
rect 42812 42662 42868 42700
rect 43036 42754 43092 43372
rect 43148 43314 43204 46508
rect 43148 43262 43150 43314
rect 43202 43262 43204 43314
rect 43148 43250 43204 43262
rect 43260 44436 43316 44446
rect 43036 42702 43038 42754
rect 43090 42702 43092 42754
rect 43036 42690 43092 42702
rect 42924 42642 42980 42654
rect 42924 42590 42926 42642
rect 42978 42590 42980 42642
rect 42924 42532 42980 42590
rect 42588 42476 42980 42532
rect 42476 42018 42532 42028
rect 42812 42308 42868 42318
rect 42028 41918 42030 41970
rect 42082 41918 42084 41970
rect 42028 41906 42084 41918
rect 42252 41860 42308 41870
rect 41916 41692 42196 41748
rect 42140 41298 42196 41692
rect 42140 41246 42142 41298
rect 42194 41246 42196 41298
rect 41692 40574 41694 40626
rect 41746 40574 41748 40626
rect 41692 40562 41748 40574
rect 41916 40964 41972 40974
rect 41916 40514 41972 40908
rect 41916 40462 41918 40514
rect 41970 40462 41972 40514
rect 41916 40450 41972 40462
rect 42140 40514 42196 41246
rect 42140 40462 42142 40514
rect 42194 40462 42196 40514
rect 42140 40450 42196 40462
rect 42252 41186 42308 41804
rect 42252 41134 42254 41186
rect 42306 41134 42308 41186
rect 41580 40404 41636 40414
rect 41580 39508 41636 40348
rect 42252 40404 42308 41134
rect 42700 41188 42756 41198
rect 42700 41094 42756 41132
rect 42700 40404 42756 40414
rect 42252 40338 42308 40348
rect 42588 40402 42756 40404
rect 42588 40350 42702 40402
rect 42754 40350 42756 40402
rect 42588 40348 42756 40350
rect 41692 39732 41748 39742
rect 41692 39638 41748 39676
rect 42588 39618 42644 40348
rect 42700 40338 42756 40348
rect 42812 40292 42868 42252
rect 42924 40628 42980 42476
rect 42924 40562 42980 40572
rect 43036 41412 43092 41422
rect 43036 40626 43092 41356
rect 43036 40574 43038 40626
rect 43090 40574 43092 40626
rect 42924 40292 42980 40302
rect 42812 40290 42980 40292
rect 42812 40238 42926 40290
rect 42978 40238 42980 40290
rect 42812 40236 42980 40238
rect 42924 40226 42980 40236
rect 42588 39566 42590 39618
rect 42642 39566 42644 39618
rect 41580 39452 41748 39508
rect 40348 38612 40516 38668
rect 40124 37426 40180 37436
rect 40460 38050 40516 38612
rect 40460 37998 40462 38050
rect 40514 37998 40516 38050
rect 40460 37268 40516 37998
rect 40460 37202 40516 37212
rect 40572 38612 40852 38668
rect 41132 38892 41524 38948
rect 40572 38162 40628 38612
rect 40796 38276 40852 38286
rect 40796 38182 40852 38220
rect 40572 38110 40574 38162
rect 40626 38110 40628 38162
rect 40348 37154 40404 37166
rect 40348 37102 40350 37154
rect 40402 37102 40404 37154
rect 40236 36258 40292 36270
rect 40236 36206 40238 36258
rect 40290 36206 40292 36258
rect 40236 34916 40292 36206
rect 40348 36260 40404 37102
rect 40572 36596 40628 38110
rect 40908 37380 40964 37390
rect 40796 37156 40852 37166
rect 40796 37062 40852 37100
rect 40572 36530 40628 36540
rect 40572 36372 40628 36382
rect 40572 36278 40628 36316
rect 40348 36194 40404 36204
rect 40908 35698 40964 37324
rect 40908 35646 40910 35698
rect 40962 35646 40964 35698
rect 40908 35634 40964 35646
rect 41020 36258 41076 36270
rect 41020 36206 41022 36258
rect 41074 36206 41076 36258
rect 41020 35588 41076 36206
rect 41020 35522 41076 35532
rect 40684 35474 40740 35486
rect 40684 35422 40686 35474
rect 40738 35422 40740 35474
rect 40236 34850 40292 34860
rect 40572 34914 40628 34926
rect 40572 34862 40574 34914
rect 40626 34862 40628 34914
rect 40348 34580 40404 34590
rect 40012 34412 40180 34468
rect 40012 34244 40068 34254
rect 40012 34150 40068 34188
rect 39900 33842 39956 33852
rect 40012 33348 40068 33358
rect 39788 33294 39790 33346
rect 39842 33294 39844 33346
rect 39676 33234 39732 33246
rect 39676 33182 39678 33234
rect 39730 33182 39732 33234
rect 39228 33124 39284 33134
rect 39228 33030 39284 33068
rect 39676 32900 39732 33182
rect 39788 33236 39844 33294
rect 39788 33170 39844 33180
rect 39900 33292 40012 33348
rect 39676 32834 39732 32844
rect 39452 32788 39508 32798
rect 39788 32788 39844 32798
rect 39900 32788 39956 33292
rect 40012 33254 40068 33292
rect 39508 32732 39620 32788
rect 39452 32694 39508 32732
rect 38668 31490 38724 31500
rect 38780 31836 39172 31892
rect 38556 31266 38612 31276
rect 38444 30482 38500 30492
rect 38668 30772 38724 30782
rect 38108 29922 38164 29932
rect 38444 29988 38500 29998
rect 38332 29652 38388 29662
rect 38332 29558 38388 29596
rect 38444 29650 38500 29932
rect 38444 29598 38446 29650
rect 38498 29598 38500 29650
rect 38444 29586 38500 29598
rect 37996 29486 37998 29538
rect 38050 29486 38052 29538
rect 37996 28980 38052 29486
rect 38220 29540 38276 29550
rect 38220 29446 38276 29484
rect 37996 28914 38052 28924
rect 38556 28980 38612 28990
rect 38556 28644 38612 28924
rect 38556 28578 38612 28588
rect 37884 28018 37940 28028
rect 37996 28530 38052 28542
rect 37996 28478 37998 28530
rect 38050 28478 38052 28530
rect 37660 27804 37940 27860
rect 37548 27682 37604 27692
rect 37772 27636 37828 27646
rect 37436 27356 37604 27412
rect 37324 27122 37380 27132
rect 37548 26852 37604 27356
rect 37548 26850 37716 26852
rect 37548 26798 37550 26850
rect 37602 26798 37716 26850
rect 37548 26796 37716 26798
rect 37548 26786 37604 26796
rect 37100 26572 37604 26628
rect 36988 25554 37044 25564
rect 37436 26290 37492 26302
rect 37436 26238 37438 26290
rect 37490 26238 37492 26290
rect 37436 26180 37492 26238
rect 37100 25284 37156 25294
rect 36988 25060 37044 25070
rect 36988 23268 37044 25004
rect 37100 23716 37156 25228
rect 37212 25172 37268 25182
rect 37212 24722 37268 25116
rect 37324 25060 37380 25070
rect 37324 24946 37380 25004
rect 37324 24894 37326 24946
rect 37378 24894 37380 24946
rect 37324 24882 37380 24894
rect 37212 24670 37214 24722
rect 37266 24670 37268 24722
rect 37212 23940 37268 24670
rect 37212 23874 37268 23884
rect 37436 24050 37492 26124
rect 37548 25060 37604 26572
rect 37660 25956 37716 26796
rect 37772 26516 37828 27580
rect 37884 27188 37940 27804
rect 37996 27412 38052 28478
rect 38332 28530 38388 28542
rect 38332 28478 38334 28530
rect 38386 28478 38388 28530
rect 38108 28420 38164 28430
rect 38332 28420 38388 28478
rect 38556 28420 38612 28430
rect 38108 28418 38276 28420
rect 38108 28366 38110 28418
rect 38162 28366 38276 28418
rect 38108 28364 38276 28366
rect 38332 28364 38556 28420
rect 38108 28354 38164 28364
rect 37996 27346 38052 27356
rect 38220 27188 38276 28364
rect 38556 28354 38612 28364
rect 38444 28084 38500 28094
rect 38444 27412 38500 28028
rect 38668 28084 38724 30716
rect 38668 28018 38724 28028
rect 38556 27858 38612 27870
rect 38556 27806 38558 27858
rect 38610 27806 38612 27858
rect 38556 27636 38612 27806
rect 38556 27570 38612 27580
rect 38668 27860 38724 27870
rect 38668 27412 38724 27804
rect 38444 27356 38612 27412
rect 37884 27132 38164 27188
rect 37884 26964 37940 27002
rect 37884 26898 37940 26908
rect 37772 26460 37940 26516
rect 37772 26290 37828 26302
rect 37772 26238 37774 26290
rect 37826 26238 37828 26290
rect 37772 26068 37828 26238
rect 37884 26178 37940 26460
rect 37996 26404 38052 26442
rect 37996 26338 38052 26348
rect 37884 26126 37886 26178
rect 37938 26126 37940 26178
rect 37884 26114 37940 26126
rect 37996 26180 38052 26190
rect 37772 26002 37828 26012
rect 37660 25890 37716 25900
rect 37660 25732 37716 25742
rect 37660 25394 37716 25676
rect 37772 25508 37828 25518
rect 37772 25414 37828 25452
rect 37884 25508 37940 25518
rect 37996 25508 38052 26124
rect 37884 25506 38052 25508
rect 37884 25454 37886 25506
rect 37938 25454 38052 25506
rect 37884 25452 38052 25454
rect 37884 25442 37940 25452
rect 37660 25342 37662 25394
rect 37714 25342 37716 25394
rect 37660 25284 37716 25342
rect 37660 25218 37716 25228
rect 37548 25004 38052 25060
rect 37548 24724 37604 24734
rect 37548 24630 37604 24668
rect 37772 24722 37828 24734
rect 37772 24670 37774 24722
rect 37826 24670 37828 24722
rect 37660 24610 37716 24622
rect 37660 24558 37662 24610
rect 37714 24558 37716 24610
rect 37660 24162 37716 24558
rect 37772 24276 37828 24670
rect 37772 24210 37828 24220
rect 37660 24110 37662 24162
rect 37714 24110 37716 24162
rect 37660 24098 37716 24110
rect 37436 23998 37438 24050
rect 37490 23998 37492 24050
rect 37100 23660 37380 23716
rect 36988 23212 37268 23268
rect 36988 23044 37044 23054
rect 36988 22950 37044 22988
rect 36876 22754 36932 22764
rect 36652 22166 36708 22204
rect 36988 22708 37044 22718
rect 36204 21698 36372 21700
rect 36204 21646 36206 21698
rect 36258 21646 36372 21698
rect 36204 21644 36372 21646
rect 36652 21812 36708 21822
rect 36204 21634 36260 21644
rect 36652 21476 36708 21756
rect 36652 21410 36708 21420
rect 36764 21364 36820 21374
rect 36652 20916 36708 20926
rect 36540 20860 36652 20916
rect 35756 20242 35812 20300
rect 35756 20190 35758 20242
rect 35810 20190 35812 20242
rect 35756 20178 35812 20190
rect 35868 20300 36148 20356
rect 36204 20580 36260 20590
rect 35868 20020 35924 20300
rect 35644 19964 35924 20020
rect 36092 20018 36148 20030
rect 36092 19966 36094 20018
rect 36146 19966 36148 20018
rect 35420 19740 35588 19796
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35532 19460 35588 19740
rect 35308 19404 35588 19460
rect 35084 19292 35252 19348
rect 35084 19122 35140 19134
rect 35084 19070 35086 19122
rect 35138 19070 35140 19122
rect 35084 19012 35140 19070
rect 35084 18946 35140 18956
rect 34860 18338 35028 18340
rect 34860 18286 34862 18338
rect 34914 18286 35028 18338
rect 34860 18284 35028 18286
rect 34748 18228 34804 18238
rect 34636 17892 34692 17902
rect 34636 17778 34692 17836
rect 34636 17726 34638 17778
rect 34690 17726 34692 17778
rect 34636 17714 34692 17726
rect 34748 17106 34804 18172
rect 34860 17890 34916 18284
rect 35196 18228 35252 19292
rect 35308 19234 35364 19404
rect 35308 19182 35310 19234
rect 35362 19182 35364 19234
rect 35308 19170 35364 19182
rect 35532 19122 35588 19404
rect 35532 19070 35534 19122
rect 35586 19070 35588 19122
rect 35532 19058 35588 19070
rect 34860 17838 34862 17890
rect 34914 17838 34916 17890
rect 34860 17826 34916 17838
rect 34972 18172 35252 18228
rect 35532 18452 35588 18462
rect 34972 17556 35028 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 34748 17054 34750 17106
rect 34802 17054 34804 17106
rect 34748 17042 34804 17054
rect 34860 17500 35028 17556
rect 35084 17890 35140 17902
rect 35084 17838 35086 17890
rect 35138 17838 35140 17890
rect 34524 16380 34692 16436
rect 34524 16212 34580 16222
rect 34076 15988 34132 15998
rect 34076 15894 34132 15932
rect 34300 15540 34356 15550
rect 34300 15446 34356 15484
rect 34524 14644 34580 16156
rect 34636 16100 34692 16380
rect 34636 16034 34692 16044
rect 34860 15988 34916 17500
rect 35084 17444 35140 17838
rect 35532 17890 35588 18396
rect 35644 18450 35700 19964
rect 36092 19908 36148 19966
rect 35980 19458 36036 19470
rect 35980 19406 35982 19458
rect 36034 19406 36036 19458
rect 35644 18398 35646 18450
rect 35698 18398 35700 18450
rect 35644 18386 35700 18398
rect 35756 19122 35812 19134
rect 35756 19070 35758 19122
rect 35810 19070 35812 19122
rect 35532 17838 35534 17890
rect 35586 17838 35588 17890
rect 35532 17826 35588 17838
rect 35756 17892 35812 19070
rect 35868 19124 35924 19134
rect 35868 19030 35924 19068
rect 35980 18788 36036 19406
rect 36092 19234 36148 19852
rect 36092 19182 36094 19234
rect 36146 19182 36148 19234
rect 36092 19012 36148 19182
rect 36092 18946 36148 18956
rect 35868 18732 36036 18788
rect 35868 18674 35924 18732
rect 35868 18622 35870 18674
rect 35922 18622 35924 18674
rect 35868 18610 35924 18622
rect 36204 18676 36260 20524
rect 36428 19460 36484 19470
rect 36428 19366 36484 19404
rect 36204 18610 36260 18620
rect 36428 19012 36484 19022
rect 35980 18564 36036 18574
rect 35980 18470 36036 18508
rect 36092 17892 36148 17902
rect 35756 17890 36148 17892
rect 35756 17838 36094 17890
rect 36146 17838 36148 17890
rect 35756 17836 36148 17838
rect 36092 17826 36148 17836
rect 36428 17780 36484 18956
rect 34860 15538 34916 15932
rect 34972 17388 35140 17444
rect 35308 17666 35364 17678
rect 35308 17614 35310 17666
rect 35362 17614 35364 17666
rect 34972 15876 35028 17388
rect 35196 16996 35252 17006
rect 35308 16996 35364 17614
rect 35756 17668 35812 17678
rect 35756 17666 36372 17668
rect 35756 17614 35758 17666
rect 35810 17614 36372 17666
rect 36428 17648 36484 17724
rect 35756 17612 36372 17614
rect 35756 17602 35812 17612
rect 35420 17444 35476 17454
rect 35420 17350 35476 17388
rect 36092 17332 36148 17342
rect 35532 17108 35588 17118
rect 35308 16940 35476 16996
rect 35196 16884 35252 16940
rect 35196 16828 35364 16884
rect 35308 16770 35364 16828
rect 35308 16718 35310 16770
rect 35362 16718 35364 16770
rect 35308 16706 35364 16718
rect 35420 16772 35476 16940
rect 35532 16994 35588 17052
rect 35532 16942 35534 16994
rect 35586 16942 35588 16994
rect 35532 16930 35588 16942
rect 35868 17108 35924 17118
rect 35644 16884 35700 16894
rect 35644 16790 35700 16828
rect 35420 16716 35588 16772
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35308 16212 35364 16222
rect 35084 16100 35140 16110
rect 35308 16100 35364 16156
rect 35532 16210 35588 16716
rect 35532 16158 35534 16210
rect 35586 16158 35588 16210
rect 35532 16146 35588 16158
rect 35756 16100 35812 16110
rect 35140 16044 35252 16100
rect 35084 16006 35140 16044
rect 34972 15820 35140 15876
rect 34860 15486 34862 15538
rect 34914 15486 34916 15538
rect 34860 15474 34916 15486
rect 34972 15652 35028 15662
rect 34636 14644 34692 14654
rect 34524 14642 34692 14644
rect 34524 14590 34638 14642
rect 34690 14590 34692 14642
rect 34524 14588 34692 14590
rect 34636 14578 34692 14588
rect 34300 14308 34356 14318
rect 34300 14214 34356 14252
rect 34412 13972 34468 13982
rect 34468 13916 34692 13972
rect 34412 13878 34468 13916
rect 33964 13858 34244 13860
rect 33964 13806 33966 13858
rect 34018 13806 34244 13858
rect 33964 13804 34244 13806
rect 33964 13794 34020 13804
rect 33852 13524 33908 13534
rect 33628 12964 33684 12974
rect 33628 12870 33684 12908
rect 33740 12852 33796 12862
rect 33628 12738 33684 12750
rect 33628 12686 33630 12738
rect 33682 12686 33684 12738
rect 33628 7700 33684 12686
rect 33740 11620 33796 12796
rect 33852 12068 33908 13468
rect 33964 12852 34020 12862
rect 33964 12850 34132 12852
rect 33964 12798 33966 12850
rect 34018 12798 34132 12850
rect 33964 12796 34132 12798
rect 33964 12786 34020 12796
rect 33964 12292 34020 12302
rect 33964 12198 34020 12236
rect 33852 12012 34020 12068
rect 33852 11620 33908 11630
rect 33740 11618 33908 11620
rect 33740 11566 33854 11618
rect 33906 11566 33908 11618
rect 33740 11564 33908 11566
rect 33852 11554 33908 11564
rect 33964 9380 34020 12012
rect 34076 11506 34132 12796
rect 34188 12292 34244 13804
rect 34636 13076 34692 13916
rect 34524 12852 34580 12862
rect 34524 12758 34580 12796
rect 34636 12850 34692 13020
rect 34972 12964 35028 15596
rect 35084 15092 35140 15820
rect 35196 15540 35252 16044
rect 35308 16098 35476 16100
rect 35308 16046 35310 16098
rect 35362 16046 35476 16098
rect 35308 16044 35476 16046
rect 35308 16034 35364 16044
rect 35420 15988 35476 16044
rect 35756 16006 35812 16044
rect 35420 15932 35588 15988
rect 35420 15540 35476 15550
rect 35196 15538 35476 15540
rect 35196 15486 35422 15538
rect 35474 15486 35476 15538
rect 35196 15484 35476 15486
rect 35420 15474 35476 15484
rect 35084 14306 35140 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35532 14530 35588 15932
rect 35868 15428 35924 17052
rect 36092 16882 36148 17276
rect 36316 17106 36372 17612
rect 36316 17054 36318 17106
rect 36370 17054 36372 17106
rect 36316 17042 36372 17054
rect 36092 16830 36094 16882
rect 36146 16830 36148 16882
rect 36092 16818 36148 16830
rect 36428 16996 36484 17006
rect 35532 14478 35534 14530
rect 35586 14478 35588 14530
rect 35532 14466 35588 14478
rect 35756 15426 35924 15428
rect 35756 15374 35870 15426
rect 35922 15374 35924 15426
rect 35756 15372 35924 15374
rect 35084 14254 35086 14306
rect 35138 14254 35140 14306
rect 35084 13748 35140 14254
rect 35756 13970 35812 15372
rect 35868 15362 35924 15372
rect 35980 16100 36036 16110
rect 35756 13918 35758 13970
rect 35810 13918 35812 13970
rect 35756 13906 35812 13918
rect 35980 14530 36036 16044
rect 36316 15988 36372 15998
rect 36316 15894 36372 15932
rect 36428 15988 36484 16940
rect 36540 16212 36596 20860
rect 36652 20822 36708 20860
rect 36652 20692 36708 20702
rect 36652 19908 36708 20636
rect 36764 20580 36820 21308
rect 36764 20130 36820 20524
rect 36988 20356 37044 22652
rect 36764 20078 36766 20130
rect 36818 20078 36820 20130
rect 36764 20066 36820 20078
rect 36876 20300 37044 20356
rect 37100 21700 37156 21710
rect 37100 21474 37156 21644
rect 37100 21422 37102 21474
rect 37154 21422 37156 21474
rect 37100 20356 37156 21422
rect 37212 21476 37268 23212
rect 37212 21410 37268 21420
rect 37324 21362 37380 23660
rect 37436 22148 37492 23998
rect 37884 23828 37940 23838
rect 37772 23492 37828 23502
rect 37436 22082 37492 22092
rect 37548 23154 37604 23166
rect 37548 23102 37550 23154
rect 37602 23102 37604 23154
rect 37548 21812 37604 23102
rect 37660 23042 37716 23054
rect 37660 22990 37662 23042
rect 37714 22990 37716 23042
rect 37660 22372 37716 22990
rect 37660 22306 37716 22316
rect 37548 21746 37604 21756
rect 37660 21812 37716 21822
rect 37772 21812 37828 23436
rect 37884 23380 37940 23772
rect 37884 23314 37940 23324
rect 37884 23154 37940 23166
rect 37884 23102 37886 23154
rect 37938 23102 37940 23154
rect 37884 23044 37940 23102
rect 37884 22978 37940 22988
rect 37996 22482 38052 25004
rect 38108 24724 38164 27132
rect 38220 27122 38276 27132
rect 38444 27076 38500 27086
rect 38444 26908 38500 27020
rect 38332 26852 38500 26908
rect 38556 26852 38612 27356
rect 38668 26908 38724 27356
rect 38780 27076 38836 31836
rect 39228 31780 39284 31790
rect 39564 31780 39620 32732
rect 39788 32786 39956 32788
rect 39788 32734 39790 32786
rect 39842 32734 39956 32786
rect 39788 32732 39956 32734
rect 39788 32722 39844 32732
rect 39676 32564 39732 32574
rect 39676 32470 39732 32508
rect 39900 32562 39956 32574
rect 39900 32510 39902 32562
rect 39954 32510 39956 32562
rect 39676 31780 39732 31790
rect 39116 31778 39284 31780
rect 39116 31726 39230 31778
rect 39282 31726 39284 31778
rect 39116 31724 39284 31726
rect 38892 30324 38948 30334
rect 38892 28754 38948 30268
rect 39004 30212 39060 30222
rect 39116 30212 39172 31724
rect 39228 31714 39284 31724
rect 39452 31778 39732 31780
rect 39452 31726 39678 31778
rect 39730 31726 39732 31778
rect 39452 31724 39732 31726
rect 39004 30210 39172 30212
rect 39004 30158 39006 30210
rect 39058 30158 39172 30210
rect 39004 30156 39172 30158
rect 39004 30146 39060 30156
rect 39004 29652 39060 29662
rect 39004 29538 39060 29596
rect 39004 29486 39006 29538
rect 39058 29486 39060 29538
rect 39004 29474 39060 29486
rect 38892 28702 38894 28754
rect 38946 28702 38948 28754
rect 38892 28690 38948 28702
rect 39116 27972 39172 30156
rect 39340 29764 39396 29774
rect 39340 29650 39396 29708
rect 39340 29598 39342 29650
rect 39394 29598 39396 29650
rect 39340 29586 39396 29598
rect 39340 29426 39396 29438
rect 39340 29374 39342 29426
rect 39394 29374 39396 29426
rect 39340 28868 39396 29374
rect 39340 28802 39396 28812
rect 39228 28756 39284 28766
rect 39228 28662 39284 28700
rect 39116 27524 39172 27916
rect 39228 28084 39284 28094
rect 39228 27970 39284 28028
rect 39340 28084 39396 28094
rect 39452 28084 39508 31724
rect 39676 31714 39732 31724
rect 39788 31108 39844 31118
rect 39788 31014 39844 31052
rect 39676 30994 39732 31006
rect 39676 30942 39678 30994
rect 39730 30942 39732 30994
rect 39676 30436 39732 30942
rect 39900 30660 39956 32510
rect 40124 31780 40180 34412
rect 40124 31714 40180 31724
rect 40236 33684 40292 33694
rect 39900 30594 39956 30604
rect 40236 30436 40292 33628
rect 40348 32786 40404 34524
rect 40572 34354 40628 34862
rect 40684 34802 40740 35422
rect 41020 35140 41076 35150
rect 41132 35140 41188 38892
rect 41580 38836 41636 38846
rect 41580 38742 41636 38780
rect 41692 38668 41748 39452
rect 42140 39396 42196 39406
rect 41356 38612 41748 38668
rect 41804 39394 42196 39396
rect 41804 39342 42142 39394
rect 42194 39342 42196 39394
rect 41804 39340 42196 39342
rect 41804 39058 41860 39340
rect 42140 39330 42196 39340
rect 41804 39006 41806 39058
rect 41858 39006 41860 39058
rect 41020 35138 41188 35140
rect 41020 35086 41022 35138
rect 41074 35086 41188 35138
rect 41020 35084 41188 35086
rect 41244 37268 41300 37278
rect 41020 35074 41076 35084
rect 41244 35028 41300 37212
rect 40684 34750 40686 34802
rect 40738 34750 40740 34802
rect 40684 34738 40740 34750
rect 41132 34972 41300 35028
rect 40572 34302 40574 34354
rect 40626 34302 40628 34354
rect 40572 34290 40628 34302
rect 40348 32734 40350 32786
rect 40402 32734 40404 32786
rect 40348 32722 40404 32734
rect 40460 34242 40516 34254
rect 40460 34190 40462 34242
rect 40514 34190 40516 34242
rect 40460 33908 40516 34190
rect 40460 31892 40516 33852
rect 40796 34130 40852 34142
rect 40796 34078 40798 34130
rect 40850 34078 40852 34130
rect 40572 33572 40628 33582
rect 40572 33458 40628 33516
rect 40572 33406 40574 33458
rect 40626 33406 40628 33458
rect 40572 33394 40628 33406
rect 40796 33124 40852 34078
rect 41020 33236 41076 33246
rect 40460 31890 40740 31892
rect 40460 31838 40462 31890
rect 40514 31838 40740 31890
rect 40460 31836 40740 31838
rect 40460 31826 40516 31836
rect 39676 30380 40292 30436
rect 40236 30322 40292 30380
rect 40236 30270 40238 30322
rect 40290 30270 40292 30322
rect 40236 30258 40292 30270
rect 40348 30994 40404 31006
rect 40348 30942 40350 30994
rect 40402 30942 40404 30994
rect 40348 29988 40404 30942
rect 40572 30994 40628 31006
rect 40572 30942 40574 30994
rect 40626 30942 40628 30994
rect 40572 30436 40628 30942
rect 40684 30884 40740 31836
rect 40796 31780 40852 33068
rect 40908 33122 40964 33134
rect 40908 33070 40910 33122
rect 40962 33070 40964 33122
rect 40908 32900 40964 33070
rect 40908 32834 40964 32844
rect 40908 32676 40964 32686
rect 41020 32676 41076 33180
rect 40908 32674 41076 32676
rect 40908 32622 40910 32674
rect 40962 32622 41076 32674
rect 40908 32620 41076 32622
rect 40908 32610 40964 32620
rect 40796 31724 41076 31780
rect 40908 31556 40964 31566
rect 40908 31462 40964 31500
rect 40908 31220 40964 31230
rect 40908 31126 40964 31164
rect 40796 31108 40852 31118
rect 40796 31014 40852 31052
rect 40684 30828 40964 30884
rect 40572 30380 40740 30436
rect 40460 30212 40516 30222
rect 40460 30118 40516 30156
rect 40348 29932 40628 29988
rect 40012 29876 40068 29886
rect 39676 29428 39732 29438
rect 39676 29426 39844 29428
rect 39676 29374 39678 29426
rect 39730 29374 39844 29426
rect 39676 29372 39844 29374
rect 39676 29362 39732 29372
rect 39340 28082 39508 28084
rect 39340 28030 39342 28082
rect 39394 28030 39508 28082
rect 39340 28028 39508 28030
rect 39564 28756 39620 28766
rect 39340 28018 39396 28028
rect 39228 27918 39230 27970
rect 39282 27918 39284 27970
rect 39228 27906 39284 27918
rect 39116 27458 39172 27468
rect 39340 27634 39396 27646
rect 39340 27582 39342 27634
rect 39394 27582 39396 27634
rect 39116 27300 39172 27310
rect 39004 27188 39060 27198
rect 38780 27074 38948 27076
rect 38780 27022 38782 27074
rect 38834 27022 38948 27074
rect 38780 27020 38948 27022
rect 38780 27010 38836 27020
rect 38668 26852 38836 26908
rect 38332 26740 38388 26852
rect 38556 26720 38612 26796
rect 38332 26674 38388 26684
rect 38332 26404 38388 26414
rect 38108 23716 38164 24668
rect 38220 26290 38276 26302
rect 38220 26238 38222 26290
rect 38274 26238 38276 26290
rect 38220 24500 38276 26238
rect 38332 25730 38388 26348
rect 38668 26404 38724 26414
rect 38668 26290 38724 26348
rect 38668 26238 38670 26290
rect 38722 26238 38724 26290
rect 38668 26226 38724 26238
rect 38332 25678 38334 25730
rect 38386 25678 38388 25730
rect 38332 25666 38388 25678
rect 38444 25956 38500 25966
rect 38332 25172 38388 25182
rect 38332 24946 38388 25116
rect 38332 24894 38334 24946
rect 38386 24894 38388 24946
rect 38332 24882 38388 24894
rect 38220 24444 38388 24500
rect 38108 23650 38164 23660
rect 38220 24276 38276 24286
rect 38108 23154 38164 23166
rect 38108 23102 38110 23154
rect 38162 23102 38164 23154
rect 38108 22708 38164 23102
rect 38108 22642 38164 22652
rect 37996 22430 37998 22482
rect 38050 22430 38052 22482
rect 37996 22418 38052 22430
rect 37884 22372 37940 22382
rect 37884 22258 37940 22316
rect 37884 22206 37886 22258
rect 37938 22206 37940 22258
rect 37884 22194 37940 22206
rect 37996 22258 38052 22270
rect 37996 22206 37998 22258
rect 38050 22206 38052 22258
rect 37660 21810 37828 21812
rect 37660 21758 37662 21810
rect 37714 21758 37828 21810
rect 37660 21756 37828 21758
rect 37996 22148 38052 22206
rect 37660 21746 37716 21756
rect 37324 21310 37326 21362
rect 37378 21310 37380 21362
rect 37324 21298 37380 21310
rect 37772 21588 37828 21598
rect 37660 21028 37716 21038
rect 37660 20934 37716 20972
rect 37772 20802 37828 21532
rect 37996 21588 38052 22092
rect 38108 22146 38164 22158
rect 38108 22094 38110 22146
rect 38162 22094 38164 22146
rect 38108 21700 38164 22094
rect 38108 21634 38164 21644
rect 37996 21522 38052 21532
rect 38108 21476 38164 21486
rect 38108 21382 38164 21420
rect 37772 20750 37774 20802
rect 37826 20750 37828 20802
rect 37772 20738 37828 20750
rect 37884 21362 37940 21374
rect 37884 21310 37886 21362
rect 37938 21310 37940 21362
rect 37548 20692 37604 20702
rect 37548 20690 37716 20692
rect 37548 20638 37550 20690
rect 37602 20638 37716 20690
rect 37548 20636 37716 20638
rect 37548 20626 37604 20636
rect 36876 19908 36932 20300
rect 37100 20290 37156 20300
rect 36652 19852 36820 19908
rect 36652 19234 36708 19246
rect 36652 19182 36654 19234
rect 36706 19182 36708 19234
rect 36652 18788 36708 19182
rect 36652 18722 36708 18732
rect 36652 17890 36708 17902
rect 36652 17838 36654 17890
rect 36706 17838 36708 17890
rect 36652 17106 36708 17838
rect 36652 17054 36654 17106
rect 36706 17054 36708 17106
rect 36652 16436 36708 17054
rect 36652 16370 36708 16380
rect 36540 16146 36596 16156
rect 36652 15988 36708 15998
rect 36428 15986 36596 15988
rect 36428 15934 36430 15986
rect 36482 15934 36596 15986
rect 36428 15932 36596 15934
rect 36428 15922 36484 15932
rect 36204 15538 36260 15550
rect 36540 15540 36596 15932
rect 36652 15894 36708 15932
rect 36204 15486 36206 15538
rect 36258 15486 36260 15538
rect 36092 15314 36148 15326
rect 36092 15262 36094 15314
rect 36146 15262 36148 15314
rect 36092 15092 36148 15262
rect 36092 15026 36148 15036
rect 36092 14756 36148 14766
rect 36204 14756 36260 15486
rect 36428 15484 36596 15540
rect 36428 15148 36484 15484
rect 36540 15316 36596 15326
rect 36540 15222 36596 15260
rect 36428 15092 36708 15148
rect 36092 14754 36260 14756
rect 36092 14702 36094 14754
rect 36146 14702 36260 14754
rect 36092 14700 36260 14702
rect 36092 14690 36148 14700
rect 35980 14478 35982 14530
rect 36034 14478 36036 14530
rect 35308 13748 35364 13758
rect 35084 13692 35308 13748
rect 35980 13748 36036 14478
rect 36316 14532 36372 14542
rect 36652 14532 36708 15092
rect 36764 14756 36820 19852
rect 36876 19842 36932 19852
rect 36988 20130 37044 20142
rect 36988 20078 36990 20130
rect 37042 20078 37044 20130
rect 36876 18562 36932 18574
rect 36876 18510 36878 18562
rect 36930 18510 36932 18562
rect 36876 18340 36932 18510
rect 36876 18274 36932 18284
rect 36988 18116 37044 20078
rect 37548 20020 37604 20030
rect 37548 19926 37604 19964
rect 37100 19796 37156 19806
rect 37100 19794 37492 19796
rect 37100 19742 37102 19794
rect 37154 19742 37492 19794
rect 37100 19740 37492 19742
rect 37100 19730 37156 19740
rect 37212 19348 37268 19358
rect 37100 19012 37156 19022
rect 37100 18562 37156 18956
rect 37100 18510 37102 18562
rect 37154 18510 37156 18562
rect 37100 18498 37156 18510
rect 37212 18562 37268 19292
rect 37436 18674 37492 19740
rect 37660 19234 37716 20636
rect 37884 19348 37940 21310
rect 38220 21252 38276 24220
rect 38332 24162 38388 24444
rect 38332 24110 38334 24162
rect 38386 24110 38388 24162
rect 38332 24098 38388 24110
rect 38332 23716 38388 23726
rect 38332 23622 38388 23660
rect 38444 23604 38500 25900
rect 38556 25620 38612 25630
rect 38556 23716 38612 25564
rect 38780 25618 38836 26852
rect 38780 25566 38782 25618
rect 38834 25566 38836 25618
rect 38780 25554 38836 25566
rect 38892 26516 38948 27020
rect 38892 25284 38948 26460
rect 38892 25218 38948 25228
rect 38780 24948 38836 24958
rect 39004 24948 39060 27132
rect 39116 27186 39172 27244
rect 39116 27134 39118 27186
rect 39170 27134 39172 27186
rect 39116 27122 39172 27134
rect 39228 27076 39284 27086
rect 39116 26516 39172 26526
rect 39228 26516 39284 27020
rect 39116 26514 39284 26516
rect 39116 26462 39118 26514
rect 39170 26462 39284 26514
rect 39116 26460 39284 26462
rect 39116 26450 39172 26460
rect 39340 26404 39396 27582
rect 39564 26908 39620 28700
rect 39676 28644 39732 28654
rect 39676 28550 39732 28588
rect 39788 27636 39844 29372
rect 39788 27570 39844 27580
rect 40012 28082 40068 29820
rect 40572 29876 40628 29932
rect 40124 29426 40180 29438
rect 40124 29374 40126 29426
rect 40178 29374 40180 29426
rect 40124 28308 40180 29374
rect 40348 29428 40404 29438
rect 40348 29426 40516 29428
rect 40348 29374 40350 29426
rect 40402 29374 40516 29426
rect 40348 29372 40516 29374
rect 40348 29362 40404 29372
rect 40124 28242 40180 28252
rect 40236 29314 40292 29326
rect 40236 29262 40238 29314
rect 40290 29262 40292 29314
rect 40236 28084 40292 29262
rect 40012 28030 40014 28082
rect 40066 28030 40068 28082
rect 40012 26908 40068 28030
rect 39564 26852 39732 26908
rect 39340 26402 39620 26404
rect 39340 26350 39342 26402
rect 39394 26350 39620 26402
rect 39340 26348 39620 26350
rect 39340 26338 39396 26348
rect 38780 24946 39060 24948
rect 38780 24894 38782 24946
rect 38834 24894 39060 24946
rect 38780 24892 39060 24894
rect 39116 26292 39172 26302
rect 38780 24612 38836 24892
rect 38780 24546 38836 24556
rect 38892 23940 38948 23950
rect 38892 23846 38948 23884
rect 38556 23660 38724 23716
rect 38444 23538 38500 23548
rect 38668 23380 38724 23660
rect 39004 23380 39060 23390
rect 38668 23378 39060 23380
rect 38668 23326 39006 23378
rect 39058 23326 39060 23378
rect 38668 23324 39060 23326
rect 38556 23042 38612 23054
rect 38556 22990 38558 23042
rect 38610 22990 38612 23042
rect 38556 22932 38612 22990
rect 38556 22260 38612 22876
rect 38556 22194 38612 22204
rect 38668 22484 38724 23324
rect 39004 23314 39060 23324
rect 38220 21186 38276 21196
rect 38332 22146 38388 22158
rect 38332 22094 38334 22146
rect 38386 22094 38388 22146
rect 38332 22036 38388 22094
rect 38332 21028 38388 21980
rect 38556 21474 38612 21486
rect 38556 21422 38558 21474
rect 38610 21422 38612 21474
rect 38556 21362 38612 21422
rect 38556 21310 38558 21362
rect 38610 21310 38612 21362
rect 38556 21298 38612 21310
rect 38220 20972 38388 21028
rect 38556 21140 38612 21150
rect 38108 20804 38164 20814
rect 38108 20710 38164 20748
rect 37884 19282 37940 19292
rect 37996 19908 38052 19918
rect 37660 19182 37662 19234
rect 37714 19182 37716 19234
rect 37436 18622 37438 18674
rect 37490 18622 37492 18674
rect 37436 18610 37492 18622
rect 37548 18788 37604 18798
rect 37212 18510 37214 18562
rect 37266 18510 37268 18562
rect 37212 18340 37268 18510
rect 37324 18564 37380 18574
rect 37324 18470 37380 18508
rect 37548 18564 37604 18732
rect 37548 18498 37604 18508
rect 37212 18284 37380 18340
rect 36876 17780 36932 17790
rect 36876 17686 36932 17724
rect 36876 17220 36932 17230
rect 36876 15316 36932 17164
rect 36988 17108 37044 18060
rect 36988 17042 37044 17052
rect 37100 18228 37156 18238
rect 37100 17106 37156 18172
rect 37100 17054 37102 17106
rect 37154 17054 37156 17106
rect 36988 16100 37044 16110
rect 36988 15538 37044 16044
rect 37100 15764 37156 17054
rect 37100 15698 37156 15708
rect 36988 15486 36990 15538
rect 37042 15486 37044 15538
rect 36988 15474 37044 15486
rect 37100 15540 37156 15550
rect 36876 15260 37044 15316
rect 36764 14690 36820 14700
rect 36372 14476 36484 14532
rect 36652 14476 36820 14532
rect 36316 14438 36372 14476
rect 36316 13748 36372 13758
rect 35980 13746 36372 13748
rect 35980 13694 36318 13746
rect 36370 13694 36372 13746
rect 35980 13692 36372 13694
rect 35308 13654 35364 13692
rect 36316 13682 36372 13692
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 13076 35252 13086
rect 35196 12982 35252 13020
rect 36316 13076 36372 13086
rect 36428 13076 36484 14476
rect 36540 14420 36596 14430
rect 36540 14326 36596 14364
rect 36652 14306 36708 14318
rect 36652 14254 36654 14306
rect 36706 14254 36708 14306
rect 36540 13748 36596 13758
rect 36540 13654 36596 13692
rect 36316 13074 36484 13076
rect 36316 13022 36318 13074
rect 36370 13022 36484 13074
rect 36316 13020 36484 13022
rect 36316 13010 36372 13020
rect 34972 12908 35140 12964
rect 34636 12798 34638 12850
rect 34690 12798 34692 12850
rect 34636 12786 34692 12798
rect 34860 12738 34916 12750
rect 34860 12686 34862 12738
rect 34914 12686 34916 12738
rect 34412 12292 34468 12302
rect 34188 12290 34468 12292
rect 34188 12238 34414 12290
rect 34466 12238 34468 12290
rect 34188 12236 34468 12238
rect 34076 11454 34078 11506
rect 34130 11454 34132 11506
rect 34076 11442 34132 11454
rect 34412 11508 34468 12236
rect 34860 12292 34916 12686
rect 34860 12226 34916 12236
rect 34412 11442 34468 11452
rect 34636 11954 34692 11966
rect 34972 11956 35028 11966
rect 34636 11902 34638 11954
rect 34690 11902 34692 11954
rect 34076 11172 34132 11182
rect 34076 11078 34132 11116
rect 34636 11172 34692 11902
rect 34636 11078 34692 11116
rect 34748 11954 35028 11956
rect 34748 11902 34974 11954
rect 35026 11902 35028 11954
rect 34748 11900 35028 11902
rect 34748 10610 34804 11900
rect 34972 11890 35028 11900
rect 34748 10558 34750 10610
rect 34802 10558 34804 10610
rect 34748 10546 34804 10558
rect 34972 10722 35028 10734
rect 34972 10670 34974 10722
rect 35026 10670 35028 10722
rect 33964 9314 34020 9324
rect 34972 9044 35028 10670
rect 34972 8978 35028 8988
rect 33628 7634 33684 7644
rect 35084 6020 35140 12908
rect 35644 12738 35700 12750
rect 35644 12686 35646 12738
rect 35698 12686 35700 12738
rect 35644 12404 35700 12686
rect 35644 12338 35700 12348
rect 36092 12404 36148 12414
rect 36092 12178 36148 12348
rect 36316 12292 36372 12302
rect 36316 12198 36372 12236
rect 36092 12126 36094 12178
rect 36146 12126 36148 12178
rect 36092 12114 36148 12126
rect 35756 11956 35812 11966
rect 35756 11954 35924 11956
rect 35756 11902 35758 11954
rect 35810 11902 35924 11954
rect 35756 11900 35924 11902
rect 35756 11890 35812 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35756 11508 35812 11518
rect 35756 11414 35812 11452
rect 35308 11172 35364 11182
rect 35308 11078 35364 11116
rect 35868 10610 35924 11900
rect 36316 11172 36372 11182
rect 36204 11170 36372 11172
rect 36204 11118 36318 11170
rect 36370 11118 36372 11170
rect 36204 11116 36372 11118
rect 36204 11060 36260 11116
rect 36316 11106 36372 11116
rect 35868 10558 35870 10610
rect 35922 10558 35924 10610
rect 35868 10546 35924 10558
rect 36092 10722 36148 10734
rect 36092 10670 36094 10722
rect 36146 10670 36148 10722
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 36092 9828 36148 10670
rect 36092 9762 36148 9772
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35084 5954 35140 5964
rect 33516 5730 33572 5740
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 33852 5124 33908 5134
rect 33852 5030 33908 5068
rect 34636 5124 34692 5134
rect 34636 5030 34692 5068
rect 34188 4898 34244 4910
rect 34188 4846 34190 4898
rect 34242 4846 34244 4898
rect 34188 3556 34244 4846
rect 36204 4340 36260 11004
rect 36652 9716 36708 14254
rect 36764 13188 36820 14476
rect 36988 13972 37044 15260
rect 37100 15148 37156 15484
rect 37212 15316 37268 15354
rect 37212 15250 37268 15260
rect 37100 15092 37268 15148
rect 36988 13906 37044 13916
rect 37100 14980 37156 14990
rect 36764 13074 36820 13132
rect 36764 13022 36766 13074
rect 36818 13022 36820 13074
rect 36764 13010 36820 13022
rect 36876 12740 36932 12750
rect 36876 12290 36932 12684
rect 36876 12238 36878 12290
rect 36930 12238 36932 12290
rect 36876 12226 36932 12238
rect 36876 11844 36932 11854
rect 36876 11506 36932 11788
rect 36876 11454 36878 11506
rect 36930 11454 36932 11506
rect 36876 11442 36932 11454
rect 36652 9650 36708 9660
rect 36876 8932 36932 8942
rect 36876 8838 36932 8876
rect 36316 6132 36372 6142
rect 36316 6038 36372 6076
rect 36876 5794 36932 5806
rect 36876 5742 36878 5794
rect 36930 5742 36932 5794
rect 36428 5236 36484 5246
rect 36428 5142 36484 5180
rect 36876 5124 36932 5742
rect 36876 4898 36932 5068
rect 36876 4846 36878 4898
rect 36930 4846 36932 4898
rect 36876 4450 36932 4846
rect 36876 4398 36878 4450
rect 36930 4398 36932 4450
rect 36876 4386 36932 4398
rect 36204 4274 36260 4284
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 35196 3666 35252 3678
rect 35196 3614 35198 3666
rect 35250 3614 35252 3666
rect 34524 3556 34580 3566
rect 34188 3554 34580 3556
rect 34188 3502 34526 3554
rect 34578 3502 34580 3554
rect 34188 3500 34580 3502
rect 34524 3490 34580 3500
rect 35196 3388 35252 3614
rect 32844 2706 32900 2716
rect 35084 3332 35252 3388
rect 29148 1250 29204 1260
rect 34300 924 34692 980
rect 34300 800 34356 924
rect 17164 700 17668 756
rect 22848 200 22960 800
rect 28224 200 28336 800
rect 34272 200 34384 800
rect 34636 756 34692 924
rect 35084 756 35140 3332
rect 37100 2884 37156 14924
rect 37212 14420 37268 15092
rect 37324 14644 37380 18284
rect 37660 18228 37716 19182
rect 37884 19124 37940 19134
rect 37884 19030 37940 19068
rect 37772 19012 37828 19022
rect 37772 18918 37828 18956
rect 37996 18900 38052 19852
rect 37660 18162 37716 18172
rect 37884 18844 38052 18900
rect 37436 17780 37492 17818
rect 37436 17714 37492 17724
rect 37324 14578 37380 14588
rect 37436 17556 37492 17566
rect 37212 14364 37380 14420
rect 37212 13636 37268 13646
rect 37212 13542 37268 13580
rect 37324 13412 37380 14364
rect 37212 13356 37380 13412
rect 37212 7812 37268 13356
rect 37324 13188 37380 13198
rect 37324 10834 37380 13132
rect 37324 10782 37326 10834
rect 37378 10782 37380 10834
rect 37324 10770 37380 10782
rect 37436 9716 37492 17500
rect 37548 17108 37604 17118
rect 37548 17014 37604 17052
rect 37884 16212 37940 18844
rect 38220 18674 38276 20972
rect 38332 20802 38388 20814
rect 38332 20750 38334 20802
rect 38386 20750 38388 20802
rect 38332 20692 38388 20750
rect 38332 20626 38388 20636
rect 38444 20580 38500 20590
rect 38444 20242 38500 20524
rect 38444 20190 38446 20242
rect 38498 20190 38500 20242
rect 38444 20178 38500 20190
rect 38332 19236 38388 19246
rect 38556 19236 38612 21084
rect 38332 19234 38612 19236
rect 38332 19182 38334 19234
rect 38386 19182 38612 19234
rect 38332 19180 38612 19182
rect 38332 19170 38388 19180
rect 38220 18622 38222 18674
rect 38274 18622 38276 18674
rect 38220 18610 38276 18622
rect 37996 18340 38052 18350
rect 37996 16884 38052 18284
rect 38108 18228 38164 18238
rect 38108 17666 38164 18172
rect 38108 17614 38110 17666
rect 38162 17614 38164 17666
rect 38108 17602 38164 17614
rect 38444 17554 38500 17566
rect 38444 17502 38446 17554
rect 38498 17502 38500 17554
rect 38332 17444 38388 17454
rect 37996 16790 38052 16828
rect 38220 17388 38332 17444
rect 37884 16146 37940 16156
rect 37996 16324 38052 16334
rect 37996 16098 38052 16268
rect 37996 16046 37998 16098
rect 38050 16046 38052 16098
rect 37996 16034 38052 16046
rect 38108 16100 38164 16110
rect 38108 16006 38164 16044
rect 37660 15988 37716 15998
rect 37660 15894 37716 15932
rect 37884 15988 37940 15998
rect 37548 15876 37604 15886
rect 37548 14418 37604 15820
rect 37772 15874 37828 15886
rect 37772 15822 37774 15874
rect 37826 15822 37828 15874
rect 37772 15540 37828 15822
rect 37772 15474 37828 15484
rect 37884 15426 37940 15932
rect 38108 15540 38164 15550
rect 38108 15446 38164 15484
rect 37884 15374 37886 15426
rect 37938 15374 37940 15426
rect 37884 15362 37940 15374
rect 37996 15316 38052 15326
rect 37996 15222 38052 15260
rect 37548 14366 37550 14418
rect 37602 14366 37604 14418
rect 37548 13858 37604 14366
rect 37884 14420 37940 14430
rect 37884 14326 37940 14364
rect 37660 13972 37716 13982
rect 37660 13878 37716 13916
rect 38220 13970 38276 17388
rect 38332 17312 38388 17388
rect 38444 16996 38500 17502
rect 38332 16940 38500 16996
rect 38332 15540 38388 16940
rect 38444 16548 38500 16558
rect 38444 16098 38500 16492
rect 38444 16046 38446 16098
rect 38498 16046 38500 16098
rect 38444 16034 38500 16046
rect 38332 15474 38388 15484
rect 38444 15876 38500 15886
rect 38444 15148 38500 15820
rect 38556 15540 38612 19180
rect 38668 18340 38724 22428
rect 39004 23044 39060 23054
rect 39116 23044 39172 26236
rect 39228 26178 39284 26190
rect 39228 26126 39230 26178
rect 39282 26126 39284 26178
rect 39228 26068 39284 26126
rect 39228 26002 39284 26012
rect 39564 25956 39620 26348
rect 39564 25890 39620 25900
rect 39564 25508 39620 25518
rect 39564 25414 39620 25452
rect 39452 25282 39508 25294
rect 39452 25230 39454 25282
rect 39506 25230 39508 25282
rect 39452 25172 39508 25230
rect 39452 25106 39508 25116
rect 39340 25060 39396 25070
rect 39676 25060 39732 26852
rect 39900 26852 40068 26908
rect 40124 28028 40292 28084
rect 40348 28308 40404 28318
rect 39900 25508 39956 26852
rect 40012 26290 40068 26302
rect 40012 26238 40014 26290
rect 40066 26238 40068 26290
rect 40012 26180 40068 26238
rect 40012 26114 40068 26124
rect 40124 25732 40180 28028
rect 40348 27188 40404 28252
rect 40460 27300 40516 29372
rect 40572 29092 40628 29820
rect 40684 29764 40740 30380
rect 40796 30212 40852 30222
rect 40796 30098 40852 30156
rect 40796 30046 40798 30098
rect 40850 30046 40852 30098
rect 40796 29988 40852 30046
rect 40796 29922 40852 29932
rect 40684 29698 40740 29708
rect 40796 29426 40852 29438
rect 40796 29374 40798 29426
rect 40850 29374 40852 29426
rect 40796 29204 40852 29374
rect 40796 29138 40852 29148
rect 40572 29026 40628 29036
rect 40796 28980 40852 28990
rect 40684 28642 40740 28654
rect 40684 28590 40686 28642
rect 40738 28590 40740 28642
rect 40572 28530 40628 28542
rect 40572 28478 40574 28530
rect 40626 28478 40628 28530
rect 40572 28196 40628 28478
rect 40572 28130 40628 28140
rect 40572 27972 40628 27982
rect 40572 27878 40628 27916
rect 40460 27244 40628 27300
rect 40236 27076 40292 27086
rect 40348 27076 40404 27132
rect 40236 27074 40404 27076
rect 40236 27022 40238 27074
rect 40290 27022 40404 27074
rect 40236 27020 40404 27022
rect 40572 27076 40628 27244
rect 40684 27298 40740 28590
rect 40796 28418 40852 28924
rect 40796 28366 40798 28418
rect 40850 28366 40852 28418
rect 40796 28354 40852 28366
rect 40908 27748 40964 30828
rect 40908 27682 40964 27692
rect 40684 27246 40686 27298
rect 40738 27246 40740 27298
rect 40684 27234 40740 27246
rect 40684 27076 40740 27086
rect 40572 27074 40740 27076
rect 40572 27022 40686 27074
rect 40738 27022 40740 27074
rect 40572 27020 40740 27022
rect 40236 27010 40292 27020
rect 40460 26964 40516 26974
rect 39340 24052 39396 25004
rect 39564 25004 39732 25060
rect 39788 25452 39956 25508
rect 40012 25676 40180 25732
rect 40236 26852 40292 26862
rect 40236 26514 40292 26796
rect 40236 26462 40238 26514
rect 40290 26462 40292 26514
rect 39452 24948 39508 24958
rect 39564 24948 39620 25004
rect 39452 24946 39620 24948
rect 39452 24894 39454 24946
rect 39506 24894 39620 24946
rect 39452 24892 39620 24894
rect 39452 24882 39508 24892
rect 39340 23986 39396 23996
rect 39788 23940 39844 25452
rect 39900 25284 39956 25294
rect 39900 24722 39956 25228
rect 39900 24670 39902 24722
rect 39954 24670 39956 24722
rect 39900 24658 39956 24670
rect 39676 23884 39844 23940
rect 39340 23828 39396 23838
rect 39060 22988 39172 23044
rect 39228 23716 39284 23726
rect 39004 22484 39060 22988
rect 39004 22482 39172 22484
rect 39004 22430 39006 22482
rect 39058 22430 39172 22482
rect 39004 22428 39172 22430
rect 39004 22418 39060 22428
rect 39004 21476 39060 21486
rect 39004 21382 39060 21420
rect 38892 21252 38948 21262
rect 38892 20914 38948 21196
rect 38892 20862 38894 20914
rect 38946 20862 38948 20914
rect 38892 20850 38948 20862
rect 39116 20244 39172 22428
rect 39116 20178 39172 20188
rect 39116 20018 39172 20030
rect 39116 19966 39118 20018
rect 39170 19966 39172 20018
rect 38892 19234 38948 19246
rect 38892 19182 38894 19234
rect 38946 19182 38948 19234
rect 38780 18676 38836 18686
rect 38780 18582 38836 18620
rect 38892 18564 38948 19182
rect 39116 19122 39172 19966
rect 39228 19906 39284 23660
rect 39340 21476 39396 23772
rect 39452 22148 39508 22158
rect 39452 22054 39508 22092
rect 39340 21410 39396 21420
rect 39452 21474 39508 21486
rect 39452 21422 39454 21474
rect 39506 21422 39508 21474
rect 39452 21364 39508 21422
rect 39340 20580 39396 20590
rect 39452 20580 39508 21308
rect 39340 20578 39508 20580
rect 39340 20526 39342 20578
rect 39394 20526 39508 20578
rect 39340 20524 39508 20526
rect 39340 20514 39396 20524
rect 39228 19854 39230 19906
rect 39282 19854 39284 19906
rect 39228 19842 39284 19854
rect 39340 20018 39396 20030
rect 39340 19966 39342 20018
rect 39394 19966 39396 20018
rect 39116 19070 39118 19122
rect 39170 19070 39172 19122
rect 39116 19012 39172 19070
rect 39116 18946 39172 18956
rect 39228 19124 39284 19134
rect 39340 19124 39396 19966
rect 39452 19908 39508 20524
rect 39564 20916 39620 20926
rect 39564 20242 39620 20860
rect 39676 20468 39732 23884
rect 39788 23714 39844 23726
rect 39788 23662 39790 23714
rect 39842 23662 39844 23714
rect 39788 23604 39844 23662
rect 40012 23604 40068 25676
rect 40124 25508 40180 25518
rect 40236 25508 40292 26462
rect 40124 25506 40292 25508
rect 40124 25454 40126 25506
rect 40178 25454 40292 25506
rect 40124 25452 40292 25454
rect 40348 26628 40404 26638
rect 40124 25442 40180 25452
rect 40348 25394 40404 26572
rect 40460 26290 40516 26908
rect 40684 26852 40740 27020
rect 40684 26786 40740 26796
rect 41020 26404 41076 31724
rect 41132 28308 41188 34972
rect 41244 34804 41300 34814
rect 41244 34244 41300 34748
rect 41244 33236 41300 34188
rect 41244 33170 41300 33180
rect 41244 30100 41300 30110
rect 41244 30006 41300 30044
rect 41356 28980 41412 38612
rect 41692 38052 41748 38062
rect 41580 38050 41748 38052
rect 41580 37998 41694 38050
rect 41746 37998 41748 38050
rect 41580 37996 41748 37998
rect 41468 37940 41524 37950
rect 41468 37846 41524 37884
rect 41580 36596 41636 37996
rect 41692 37986 41748 37996
rect 41692 37380 41748 37390
rect 41692 37286 41748 37324
rect 41804 37266 41860 39006
rect 42028 38948 42084 38958
rect 42028 38854 42084 38892
rect 42476 38836 42532 38846
rect 41916 38724 41972 38762
rect 41916 38658 41972 38668
rect 42028 38500 42084 38510
rect 42028 38274 42084 38444
rect 42028 38222 42030 38274
rect 42082 38222 42084 38274
rect 42028 38210 42084 38222
rect 41804 37214 41806 37266
rect 41858 37214 41860 37266
rect 41804 37044 41860 37214
rect 41916 37268 41972 37278
rect 41916 37174 41972 37212
rect 42476 37268 42532 38780
rect 42588 38724 42644 39566
rect 42812 40068 42868 40078
rect 42812 39508 42868 40012
rect 43036 39508 43092 40574
rect 43260 41076 43316 44380
rect 43372 43204 43428 47964
rect 43484 47954 43540 47964
rect 43708 47796 43764 47806
rect 43484 47458 43540 47470
rect 43484 47406 43486 47458
rect 43538 47406 43540 47458
rect 43484 46676 43540 47406
rect 43708 47346 43764 47740
rect 43708 47294 43710 47346
rect 43762 47294 43764 47346
rect 43708 47282 43764 47294
rect 43708 46676 43764 46686
rect 43484 46674 43652 46676
rect 43484 46622 43486 46674
rect 43538 46622 43652 46674
rect 43484 46620 43652 46622
rect 43484 46610 43540 46620
rect 43484 45892 43540 45902
rect 43484 45798 43540 45836
rect 43596 44884 43652 46620
rect 43708 46002 43764 46620
rect 43708 45950 43710 46002
rect 43762 45950 43764 46002
rect 43708 45938 43764 45950
rect 43820 45332 43876 48076
rect 44156 48130 44212 48142
rect 44156 48078 44158 48130
rect 44210 48078 44212 48130
rect 44156 47684 44212 48078
rect 44156 47618 44212 47628
rect 44044 47460 44100 47470
rect 44044 47366 44100 47404
rect 44380 47346 44436 48748
rect 44380 47294 44382 47346
rect 44434 47294 44436 47346
rect 44380 47282 44436 47294
rect 44492 48802 44548 49644
rect 44604 49606 44660 49644
rect 44492 48750 44494 48802
rect 44546 48750 44548 48802
rect 44492 47124 44548 48750
rect 44604 48130 44660 48142
rect 44604 48078 44606 48130
rect 44658 48078 44660 48130
rect 44604 48020 44660 48078
rect 44604 47954 44660 47964
rect 44828 47908 44884 51214
rect 45052 51044 45108 51660
rect 46284 51604 46340 51886
rect 46284 51538 46340 51548
rect 46396 51492 46452 52782
rect 46508 52052 46564 52062
rect 46508 51958 46564 51996
rect 46844 51604 46900 52894
rect 47180 52946 47236 52958
rect 47180 52894 47182 52946
rect 47234 52894 47236 52946
rect 47068 52276 47124 52286
rect 47068 52182 47124 52220
rect 47180 51940 47236 52894
rect 47404 52948 47460 52958
rect 47404 52946 47572 52948
rect 47404 52894 47406 52946
rect 47458 52894 47572 52946
rect 47404 52892 47572 52894
rect 47404 52882 47460 52892
rect 47180 51874 47236 51884
rect 47516 52052 47572 52892
rect 47964 52836 48020 52846
rect 47852 52834 48020 52836
rect 47852 52782 47966 52834
rect 48018 52782 48020 52834
rect 47852 52780 48020 52782
rect 46844 51538 46900 51548
rect 46396 51426 46452 51436
rect 47292 51492 47348 51502
rect 47292 51378 47348 51436
rect 47292 51326 47294 51378
rect 47346 51326 47348 51378
rect 47292 51314 47348 51326
rect 45052 50978 45108 50988
rect 45164 51266 45220 51278
rect 45164 51214 45166 51266
rect 45218 51214 45220 51266
rect 45164 50428 45220 51214
rect 45724 51268 45780 51278
rect 46172 51268 46228 51278
rect 46508 51268 46564 51278
rect 45724 51266 46228 51268
rect 45724 51214 45726 51266
rect 45778 51214 46174 51266
rect 46226 51214 46228 51266
rect 45724 51212 46228 51214
rect 45724 51202 45780 51212
rect 45388 50596 45444 50606
rect 45388 50502 45444 50540
rect 45052 50372 45220 50428
rect 45724 50484 45780 50494
rect 45724 50390 45780 50428
rect 45052 49700 45108 50372
rect 45612 50370 45668 50382
rect 45612 50318 45614 50370
rect 45666 50318 45668 50370
rect 45612 50036 45668 50318
rect 45612 49970 45668 49980
rect 45052 49634 45108 49644
rect 45164 49698 45220 49710
rect 45164 49646 45166 49698
rect 45218 49646 45220 49698
rect 44828 47842 44884 47852
rect 45052 48130 45108 48142
rect 45052 48078 45054 48130
rect 45106 48078 45108 48130
rect 44604 47124 44660 47134
rect 44492 47068 44604 47124
rect 44268 46900 44324 46910
rect 44268 46806 44324 46844
rect 44492 46900 44548 46910
rect 44044 46676 44100 46686
rect 44044 46582 44100 46620
rect 44156 46562 44212 46574
rect 44156 46510 44158 46562
rect 44210 46510 44212 46562
rect 44156 45668 44212 46510
rect 44492 45892 44548 46844
rect 44604 46674 44660 47068
rect 45052 46788 45108 48078
rect 45052 46694 45108 46732
rect 44604 46622 44606 46674
rect 44658 46622 44660 46674
rect 44604 46610 44660 46622
rect 44716 46676 44772 46686
rect 43820 45266 43876 45276
rect 43932 45612 44212 45668
rect 44380 45666 44436 45678
rect 44380 45614 44382 45666
rect 44434 45614 44436 45666
rect 43932 45218 43988 45612
rect 44380 45556 44436 45614
rect 43932 45166 43934 45218
rect 43986 45166 43988 45218
rect 43932 45154 43988 45166
rect 44044 45500 44436 45556
rect 43372 43138 43428 43148
rect 43484 44828 43652 44884
rect 43820 45106 43876 45118
rect 43820 45054 43822 45106
rect 43874 45054 43876 45106
rect 43484 42978 43540 44828
rect 43484 42926 43486 42978
rect 43538 42926 43540 42978
rect 43484 42914 43540 42926
rect 43596 44098 43652 44110
rect 43596 44046 43598 44098
rect 43650 44046 43652 44098
rect 43596 41412 43652 44046
rect 43820 43540 43876 45054
rect 43932 44436 43988 44446
rect 43932 44342 43988 44380
rect 43708 43426 43764 43438
rect 43708 43374 43710 43426
rect 43762 43374 43764 43426
rect 43708 43092 43764 43374
rect 43708 42532 43764 43036
rect 43820 42980 43876 43484
rect 43820 42914 43876 42924
rect 44044 43876 44100 45500
rect 44044 42642 44100 43820
rect 44044 42590 44046 42642
rect 44098 42590 44100 42642
rect 44044 42578 44100 42590
rect 44156 45332 44212 45342
rect 43708 42466 43764 42476
rect 43820 41970 43876 41982
rect 43820 41918 43822 41970
rect 43874 41918 43876 41970
rect 43820 41860 43876 41918
rect 43820 41794 43876 41804
rect 43596 41346 43652 41356
rect 44044 41300 44100 41310
rect 43260 40626 43316 41020
rect 43596 41186 43652 41198
rect 43596 41134 43598 41186
rect 43650 41134 43652 41186
rect 43596 40852 43652 41134
rect 43596 40786 43652 40796
rect 43820 40962 43876 40974
rect 43820 40910 43822 40962
rect 43874 40910 43876 40962
rect 43260 40574 43262 40626
rect 43314 40574 43316 40626
rect 42812 39442 42868 39452
rect 42924 39506 43092 39508
rect 42924 39454 43038 39506
rect 43090 39454 43092 39506
rect 42924 39452 43092 39454
rect 42588 38658 42644 38668
rect 42476 37202 42532 37212
rect 42812 37268 42868 37278
rect 42812 37174 42868 37212
rect 42028 37156 42084 37166
rect 42028 37044 42084 37100
rect 41804 36988 42084 37044
rect 41580 36530 41636 36540
rect 41580 36258 41636 36270
rect 41580 36206 41582 36258
rect 41634 36206 41636 36258
rect 41468 35588 41524 35626
rect 41468 35522 41524 35532
rect 41468 35364 41524 35374
rect 41468 33124 41524 35308
rect 41580 34804 41636 36206
rect 41916 36258 41972 36270
rect 41916 36206 41918 36258
rect 41970 36206 41972 36258
rect 41916 35586 41972 36206
rect 41916 35534 41918 35586
rect 41970 35534 41972 35586
rect 41916 35252 41972 35534
rect 42028 35476 42084 36988
rect 42364 37044 42420 37054
rect 42588 37044 42644 37054
rect 42364 37042 42644 37044
rect 42364 36990 42366 37042
rect 42418 36990 42590 37042
rect 42642 36990 42644 37042
rect 42364 36988 42644 36990
rect 42364 36978 42420 36988
rect 42588 36978 42644 36988
rect 42476 36260 42532 36270
rect 42476 36166 42532 36204
rect 42924 36036 42980 39452
rect 43036 39442 43092 39452
rect 43148 40516 43204 40526
rect 43148 39506 43204 40460
rect 43260 40404 43316 40574
rect 43260 40348 43428 40404
rect 43260 39732 43316 39770
rect 43260 39666 43316 39676
rect 43372 39620 43428 40348
rect 43372 39618 43540 39620
rect 43372 39566 43374 39618
rect 43426 39566 43540 39618
rect 43372 39564 43540 39566
rect 43372 39554 43428 39564
rect 43148 39454 43150 39506
rect 43202 39454 43204 39506
rect 43148 39442 43204 39454
rect 43260 39508 43316 39518
rect 43148 39060 43204 39070
rect 43148 38946 43204 39004
rect 43148 38894 43150 38946
rect 43202 38894 43204 38946
rect 43148 37938 43204 38894
rect 43148 37886 43150 37938
rect 43202 37886 43204 37938
rect 43148 37604 43204 37886
rect 43260 37938 43316 39452
rect 43372 38164 43428 38174
rect 43372 38070 43428 38108
rect 43260 37886 43262 37938
rect 43314 37886 43316 37938
rect 43260 37874 43316 37886
rect 43148 37538 43204 37548
rect 43372 37826 43428 37838
rect 43372 37774 43374 37826
rect 43426 37774 43428 37826
rect 43036 37380 43092 37390
rect 43036 36370 43092 37324
rect 43260 37156 43316 37166
rect 43260 37062 43316 37100
rect 43372 37044 43428 37774
rect 43372 36978 43428 36988
rect 43036 36318 43038 36370
rect 43090 36318 43092 36370
rect 43036 36306 43092 36318
rect 43260 36370 43316 36382
rect 43260 36318 43262 36370
rect 43314 36318 43316 36370
rect 42812 35980 42980 36036
rect 43148 36258 43204 36270
rect 43148 36206 43150 36258
rect 43202 36206 43204 36258
rect 42028 35420 42532 35476
rect 41916 35186 41972 35196
rect 42140 35026 42196 35038
rect 42140 34974 42142 35026
rect 42194 34974 42196 35026
rect 41580 34738 41636 34748
rect 42028 34914 42084 34926
rect 42028 34862 42030 34914
rect 42082 34862 42084 34914
rect 41692 34130 41748 34142
rect 41692 34078 41694 34130
rect 41746 34078 41748 34130
rect 41580 33348 41636 33358
rect 41692 33348 41748 34078
rect 41916 34130 41972 34142
rect 41916 34078 41918 34130
rect 41970 34078 41972 34130
rect 41916 33460 41972 34078
rect 42028 33684 42084 34862
rect 42140 34242 42196 34974
rect 42140 34190 42142 34242
rect 42194 34190 42196 34242
rect 42140 34178 42196 34190
rect 42252 34692 42308 34702
rect 42028 33618 42084 33628
rect 41636 33292 41748 33348
rect 41804 33404 41972 33460
rect 41580 33216 41636 33292
rect 41804 33234 41860 33404
rect 42028 33348 42084 33358
rect 41804 33182 41806 33234
rect 41858 33182 41860 33234
rect 41692 33124 41748 33134
rect 41468 33122 41748 33124
rect 41468 33070 41694 33122
rect 41746 33070 41748 33122
rect 41468 33068 41748 33070
rect 41692 33058 41748 33068
rect 41692 32900 41748 32910
rect 41468 32562 41524 32574
rect 41468 32510 41470 32562
rect 41522 32510 41524 32562
rect 41468 32452 41524 32510
rect 41468 32386 41524 32396
rect 41580 32116 41636 32126
rect 41468 31780 41524 31790
rect 41468 31686 41524 31724
rect 41468 30882 41524 30894
rect 41468 30830 41470 30882
rect 41522 30830 41524 30882
rect 41468 30660 41524 30830
rect 41468 30594 41524 30604
rect 41580 30436 41636 32060
rect 41468 30380 41636 30436
rect 41468 29204 41524 30380
rect 41692 29652 41748 32844
rect 41804 32786 41860 33182
rect 41916 33236 41972 33246
rect 41916 33142 41972 33180
rect 42028 33234 42084 33292
rect 42028 33182 42030 33234
rect 42082 33182 42084 33234
rect 41804 32734 41806 32786
rect 41858 32734 41860 32786
rect 41804 32722 41860 32734
rect 41916 32562 41972 32574
rect 41916 32510 41918 32562
rect 41970 32510 41972 32562
rect 41916 32004 41972 32510
rect 41916 31938 41972 31948
rect 42028 31780 42084 33182
rect 42252 32788 42308 34636
rect 42140 32732 42308 32788
rect 42140 32674 42196 32732
rect 42140 32622 42142 32674
rect 42194 32622 42196 32674
rect 42140 32610 42196 32622
rect 41692 29586 41748 29596
rect 41804 31724 42084 31780
rect 42252 32564 42308 32574
rect 41580 29540 41636 29550
rect 41580 29446 41636 29484
rect 41468 29138 41524 29148
rect 41356 28914 41412 28924
rect 41804 28644 41860 31724
rect 42028 31554 42084 31566
rect 42028 31502 42030 31554
rect 42082 31502 42084 31554
rect 42028 31332 42084 31502
rect 42028 31266 42084 31276
rect 42252 30996 42308 32508
rect 42028 30940 42308 30996
rect 42028 30210 42084 30940
rect 42140 30772 42196 30782
rect 42364 30772 42420 30782
rect 42140 30678 42196 30716
rect 42252 30770 42420 30772
rect 42252 30718 42366 30770
rect 42418 30718 42420 30770
rect 42252 30716 42420 30718
rect 42028 30158 42030 30210
rect 42082 30158 42084 30210
rect 41916 29428 41972 29438
rect 41916 29334 41972 29372
rect 41804 28578 41860 28588
rect 41580 28532 41636 28542
rect 41132 28252 41412 28308
rect 41244 27748 41300 27758
rect 41132 27636 41188 27646
rect 41132 26964 41188 27580
rect 41132 26898 41188 26908
rect 40908 26348 41076 26404
rect 40460 26238 40462 26290
rect 40514 26238 40516 26290
rect 40460 26226 40516 26238
rect 40572 26292 40628 26302
rect 40572 25730 40628 26236
rect 40572 25678 40574 25730
rect 40626 25678 40628 25730
rect 40572 25666 40628 25678
rect 40684 26290 40740 26302
rect 40684 26238 40686 26290
rect 40738 26238 40740 26290
rect 40684 25620 40740 26238
rect 40796 26180 40852 26190
rect 40796 26086 40852 26124
rect 40684 25554 40740 25564
rect 40348 25342 40350 25394
rect 40402 25342 40404 25394
rect 40236 25172 40292 25182
rect 39788 23538 39844 23548
rect 39900 23548 40068 23604
rect 40124 24498 40180 24510
rect 40124 24446 40126 24498
rect 40178 24446 40180 24498
rect 39900 23380 39956 23548
rect 39900 23314 39956 23324
rect 40012 23380 40068 23390
rect 40124 23380 40180 24446
rect 40236 24498 40292 25116
rect 40236 24446 40238 24498
rect 40290 24446 40292 24498
rect 40236 24276 40292 24446
rect 40348 24500 40404 25342
rect 40796 25506 40852 25518
rect 40796 25454 40798 25506
rect 40850 25454 40852 25506
rect 40460 25284 40516 25294
rect 40460 25190 40516 25228
rect 40796 24836 40852 25454
rect 40348 24434 40404 24444
rect 40572 24780 40852 24836
rect 40236 24220 40404 24276
rect 40236 24052 40292 24062
rect 40236 23958 40292 23996
rect 40348 23828 40404 24220
rect 40012 23378 40180 23380
rect 40012 23326 40014 23378
rect 40066 23326 40180 23378
rect 40012 23324 40180 23326
rect 40236 23772 40404 23828
rect 40012 23314 40068 23324
rect 39788 23156 39844 23166
rect 39788 23154 39956 23156
rect 39788 23102 39790 23154
rect 39842 23102 39956 23154
rect 39788 23100 39956 23102
rect 39788 23090 39844 23100
rect 39900 21812 39956 23100
rect 40124 23154 40180 23166
rect 40124 23102 40126 23154
rect 40178 23102 40180 23154
rect 40124 22482 40180 23102
rect 40124 22430 40126 22482
rect 40178 22430 40180 22482
rect 40124 22418 40180 22430
rect 40236 22484 40292 23772
rect 40348 23268 40404 23278
rect 40348 23174 40404 23212
rect 40236 22418 40292 22428
rect 40012 22372 40068 22382
rect 40012 22278 40068 22316
rect 40348 22372 40404 22382
rect 40236 22148 40292 22158
rect 40236 22054 40292 22092
rect 40348 21924 40404 22316
rect 40460 22260 40516 22270
rect 40460 22166 40516 22204
rect 40236 21868 40404 21924
rect 40572 21924 40628 24780
rect 40796 24610 40852 24622
rect 40796 24558 40798 24610
rect 40850 24558 40852 24610
rect 40684 24052 40740 24062
rect 40684 23958 40740 23996
rect 40796 23828 40852 24558
rect 40684 23772 40852 23828
rect 40684 23044 40740 23772
rect 40908 23548 40964 26348
rect 41020 25394 41076 25406
rect 41020 25342 41022 25394
rect 41074 25342 41076 25394
rect 41020 25284 41076 25342
rect 41020 25218 41076 25228
rect 40684 22978 40740 22988
rect 40796 23492 40964 23548
rect 41020 24388 41076 24398
rect 40124 21812 40180 21822
rect 39900 21810 40180 21812
rect 39900 21758 40126 21810
rect 40178 21758 40180 21810
rect 39900 21756 40180 21758
rect 40124 21746 40180 21756
rect 40012 21586 40068 21598
rect 40012 21534 40014 21586
rect 40066 21534 40068 21586
rect 40012 21028 40068 21534
rect 40012 20962 40068 20972
rect 40124 21588 40180 21598
rect 40124 20802 40180 21532
rect 40124 20750 40126 20802
rect 40178 20750 40180 20802
rect 40124 20738 40180 20750
rect 39900 20692 39956 20702
rect 39900 20598 39956 20636
rect 39676 20412 40068 20468
rect 39564 20190 39566 20242
rect 39618 20190 39620 20242
rect 39564 20178 39620 20190
rect 39452 19852 39620 19908
rect 39452 19124 39508 19134
rect 39340 19068 39452 19124
rect 39116 18564 39172 18574
rect 38892 18508 39116 18564
rect 39116 18470 39172 18508
rect 38668 18284 39060 18340
rect 39004 17778 39060 18284
rect 39004 17726 39006 17778
rect 39058 17726 39060 17778
rect 39004 17108 39060 17726
rect 39116 17108 39172 17118
rect 39004 17106 39172 17108
rect 39004 17054 39118 17106
rect 39170 17054 39172 17106
rect 39004 17052 39172 17054
rect 38892 16884 38948 16894
rect 38892 16882 39060 16884
rect 38892 16830 38894 16882
rect 38946 16830 39060 16882
rect 38892 16828 39060 16830
rect 38892 16818 38948 16828
rect 39004 16100 39060 16828
rect 39116 16324 39172 17052
rect 39116 16258 39172 16268
rect 39228 16212 39284 19068
rect 39452 19058 39508 19068
rect 39564 18674 39620 19852
rect 40012 19236 40068 20412
rect 40124 20244 40180 20254
rect 40124 20150 40180 20188
rect 39676 19124 39732 19162
rect 40012 19142 40068 19180
rect 39676 19058 39732 19068
rect 39900 19012 39956 19022
rect 39564 18622 39566 18674
rect 39618 18622 39620 18674
rect 39564 18610 39620 18622
rect 39676 18900 39732 18910
rect 39676 17778 39732 18844
rect 39676 17726 39678 17778
rect 39730 17726 39732 17778
rect 39228 16146 39284 16156
rect 39340 16324 39396 16334
rect 39676 16324 39732 17726
rect 39900 16660 39956 18956
rect 40236 18900 40292 21868
rect 40572 21858 40628 21868
rect 40348 21588 40404 21598
rect 40348 21494 40404 21532
rect 40572 21586 40628 21598
rect 40572 21534 40574 21586
rect 40626 21534 40628 21586
rect 40572 21476 40628 21534
rect 40572 21410 40628 21420
rect 40460 21028 40516 21038
rect 40796 21028 40852 23492
rect 40908 23380 40964 23390
rect 40908 23286 40964 23324
rect 41020 22820 41076 24332
rect 40908 22764 41076 22820
rect 41132 24162 41188 24174
rect 41132 24110 41134 24162
rect 41186 24110 41188 24162
rect 40908 22372 40964 22764
rect 41020 22484 41076 22494
rect 41132 22484 41188 24110
rect 41244 24050 41300 27692
rect 41356 26180 41412 28252
rect 41580 28084 41636 28476
rect 41580 27990 41636 28028
rect 41916 27634 41972 27646
rect 41916 27582 41918 27634
rect 41970 27582 41972 27634
rect 41468 27524 41524 27534
rect 41468 27074 41524 27468
rect 41916 27412 41972 27582
rect 41916 27346 41972 27356
rect 41804 27188 41860 27198
rect 41468 27022 41470 27074
rect 41522 27022 41524 27074
rect 41468 27010 41524 27022
rect 41692 27132 41804 27188
rect 41692 27074 41748 27132
rect 41804 27122 41860 27132
rect 41692 27022 41694 27074
rect 41746 27022 41748 27074
rect 41580 26628 41636 26638
rect 41356 26114 41412 26124
rect 41468 26516 41524 26526
rect 41468 25618 41524 26460
rect 41580 26402 41636 26572
rect 41580 26350 41582 26402
rect 41634 26350 41636 26402
rect 41580 26338 41636 26350
rect 41468 25566 41470 25618
rect 41522 25566 41524 25618
rect 41468 25554 41524 25566
rect 41580 24948 41636 24958
rect 41580 24854 41636 24892
rect 41692 24276 41748 27022
rect 42028 26908 42084 30158
rect 42140 30100 42196 30110
rect 42140 30006 42196 30044
rect 42252 28084 42308 30716
rect 42364 30706 42420 30716
rect 42476 30324 42532 35420
rect 42588 32900 42644 32910
rect 42588 32450 42644 32844
rect 42588 32398 42590 32450
rect 42642 32398 42644 32450
rect 42588 32228 42644 32398
rect 42588 32162 42644 32172
rect 42700 32004 42756 32014
rect 42700 31778 42756 31948
rect 42700 31726 42702 31778
rect 42754 31726 42756 31778
rect 42700 31668 42756 31726
rect 42812 31668 42868 35980
rect 42924 35810 42980 35822
rect 42924 35758 42926 35810
rect 42978 35758 42980 35810
rect 42924 35364 42980 35758
rect 43148 35698 43204 36206
rect 43148 35646 43150 35698
rect 43202 35646 43204 35698
rect 43148 35634 43204 35646
rect 43260 36260 43316 36318
rect 42924 35298 42980 35308
rect 43036 34356 43092 34366
rect 43036 34130 43092 34300
rect 43036 34078 43038 34130
rect 43090 34078 43092 34130
rect 43036 34066 43092 34078
rect 43260 34020 43316 36204
rect 43260 33954 43316 33964
rect 43372 35812 43428 35822
rect 42924 33122 42980 33134
rect 42924 33070 42926 33122
rect 42978 33070 42980 33122
rect 42924 32900 42980 33070
rect 43260 33124 43316 33134
rect 43260 33030 43316 33068
rect 42924 32834 42980 32844
rect 43036 32564 43092 32574
rect 43036 32470 43092 32508
rect 43372 32116 43428 35756
rect 43484 35586 43540 39564
rect 43820 39508 43876 40910
rect 44044 40402 44100 41244
rect 44156 40852 44212 45276
rect 44492 45106 44548 45836
rect 44716 45892 44772 46620
rect 45164 46676 45220 49646
rect 45500 49698 45556 49710
rect 45500 49646 45502 49698
rect 45554 49646 45556 49698
rect 45388 48916 45444 48926
rect 45388 48822 45444 48860
rect 45500 48692 45556 49646
rect 45836 49476 45892 51212
rect 46172 51202 46228 51212
rect 46284 51266 46564 51268
rect 46284 51214 46510 51266
rect 46562 51214 46564 51266
rect 46284 51212 46564 51214
rect 46172 50372 46228 50382
rect 45836 49410 45892 49420
rect 46060 50370 46228 50372
rect 46060 50318 46174 50370
rect 46226 50318 46228 50370
rect 46060 50316 46228 50318
rect 45500 48626 45556 48636
rect 46060 48692 46116 50316
rect 46172 50306 46228 50316
rect 46284 49924 46340 51212
rect 46508 51202 46564 51212
rect 47516 51154 47572 51996
rect 47628 52162 47684 52174
rect 47628 52110 47630 52162
rect 47682 52110 47684 52162
rect 47628 51604 47684 52110
rect 47740 52052 47796 52062
rect 47740 51958 47796 51996
rect 47628 51538 47684 51548
rect 47740 51828 47796 51838
rect 47516 51102 47518 51154
rect 47570 51102 47572 51154
rect 47516 51090 47572 51102
rect 47404 50820 47460 50830
rect 47292 50818 47460 50820
rect 47292 50766 47406 50818
rect 47458 50766 47460 50818
rect 47292 50764 47460 50766
rect 47180 50484 47236 50494
rect 46844 50370 46900 50382
rect 46844 50318 46846 50370
rect 46898 50318 46900 50370
rect 46060 48626 46116 48636
rect 46172 49868 46340 49924
rect 46508 50036 46564 50046
rect 46172 49250 46228 49868
rect 46172 49198 46174 49250
rect 46226 49198 46228 49250
rect 45500 48130 45556 48142
rect 46060 48132 46116 48142
rect 45500 48078 45502 48130
rect 45554 48078 45556 48130
rect 45500 47908 45556 48078
rect 45500 47842 45556 47852
rect 45948 48130 46116 48132
rect 45948 48078 46062 48130
rect 46114 48078 46116 48130
rect 45948 48076 46116 48078
rect 45500 47684 45556 47694
rect 45388 47234 45444 47246
rect 45388 47182 45390 47234
rect 45442 47182 45444 47234
rect 45388 46900 45444 47182
rect 45388 46834 45444 46844
rect 45164 46610 45220 46620
rect 44604 45220 44660 45230
rect 44716 45220 44772 45836
rect 44604 45218 44772 45220
rect 44604 45166 44606 45218
rect 44658 45166 44772 45218
rect 44604 45164 44772 45166
rect 45500 45218 45556 47628
rect 45948 46900 46004 48076
rect 46060 48066 46116 48076
rect 46060 47572 46116 47582
rect 46060 47234 46116 47516
rect 46060 47182 46062 47234
rect 46114 47182 46116 47234
rect 46060 47170 46116 47182
rect 45612 46562 45668 46574
rect 45612 46510 45614 46562
rect 45666 46510 45668 46562
rect 45612 46452 45668 46510
rect 45948 46562 46004 46844
rect 45948 46510 45950 46562
rect 46002 46510 46004 46562
rect 45668 46396 45892 46452
rect 45612 46386 45668 46396
rect 45724 45780 45780 45790
rect 45724 45686 45780 45724
rect 45500 45166 45502 45218
rect 45554 45166 45556 45218
rect 44604 45154 44660 45164
rect 45500 45154 45556 45166
rect 45612 45666 45668 45678
rect 45612 45614 45614 45666
rect 45666 45614 45668 45666
rect 44492 45054 44494 45106
rect 44546 45054 44548 45106
rect 44492 45042 44548 45054
rect 45612 45106 45668 45614
rect 45612 45054 45614 45106
rect 45666 45054 45668 45106
rect 45612 45042 45668 45054
rect 45836 45668 45892 46396
rect 45388 44994 45444 45006
rect 45388 44942 45390 44994
rect 45442 44942 45444 44994
rect 44492 44098 44548 44110
rect 44492 44046 44494 44098
rect 44546 44046 44548 44098
rect 44380 43652 44436 43662
rect 44268 42756 44324 42766
rect 44268 42662 44324 42700
rect 44380 41188 44436 43596
rect 44492 42532 44548 44046
rect 45388 43764 45444 44942
rect 45836 44210 45892 45612
rect 45948 45556 46004 46510
rect 46172 46564 46228 49198
rect 46284 49698 46340 49710
rect 46284 49646 46286 49698
rect 46338 49646 46340 49698
rect 46284 48804 46340 49646
rect 46396 49140 46452 49178
rect 46396 49074 46452 49084
rect 46396 48916 46452 48926
rect 46508 48916 46564 49980
rect 46844 50036 46900 50318
rect 47180 50370 47236 50428
rect 47180 50318 47182 50370
rect 47234 50318 47236 50370
rect 47180 50306 47236 50318
rect 46844 49970 46900 49980
rect 46844 49810 46900 49822
rect 46844 49758 46846 49810
rect 46898 49758 46900 49810
rect 46844 49700 46900 49758
rect 46732 49028 46788 49038
rect 46732 48934 46788 48972
rect 46396 48914 46564 48916
rect 46396 48862 46398 48914
rect 46450 48862 46564 48914
rect 46396 48860 46564 48862
rect 46844 48916 46900 49644
rect 46956 49140 47012 49150
rect 47012 49084 47124 49140
rect 46956 49046 47012 49084
rect 46396 48850 46452 48860
rect 46844 48850 46900 48860
rect 46284 48738 46340 48748
rect 47068 48466 47124 49084
rect 47068 48414 47070 48466
rect 47122 48414 47124 48466
rect 47068 48402 47124 48414
rect 47180 48468 47236 48478
rect 47180 48374 47236 48412
rect 46732 48242 46788 48254
rect 46956 48244 47012 48254
rect 46732 48190 46734 48242
rect 46786 48190 46788 48242
rect 46508 47460 46564 47470
rect 46732 47460 46788 48190
rect 46508 47458 46788 47460
rect 46508 47406 46510 47458
rect 46562 47406 46788 47458
rect 46508 47404 46788 47406
rect 46508 47394 46564 47404
rect 46732 46786 46788 47404
rect 46732 46734 46734 46786
rect 46786 46734 46788 46786
rect 46732 46722 46788 46734
rect 46844 48242 47012 48244
rect 46844 48190 46958 48242
rect 47010 48190 47012 48242
rect 46844 48188 47012 48190
rect 46844 47346 46900 48188
rect 46956 48178 47012 48188
rect 46844 47294 46846 47346
rect 46898 47294 46900 47346
rect 46172 46498 46228 46508
rect 45948 45490 46004 45500
rect 46620 45890 46676 45902
rect 46620 45838 46622 45890
rect 46674 45838 46676 45890
rect 46060 45220 46116 45230
rect 46060 44322 46116 45164
rect 46284 45106 46340 45118
rect 46284 45054 46286 45106
rect 46338 45054 46340 45106
rect 46172 44548 46228 44558
rect 46284 44548 46340 45054
rect 46172 44546 46340 44548
rect 46172 44494 46174 44546
rect 46226 44494 46340 44546
rect 46172 44492 46340 44494
rect 46396 45108 46452 45118
rect 46172 44482 46228 44492
rect 46060 44270 46062 44322
rect 46114 44270 46116 44322
rect 46060 44258 46116 44270
rect 46396 44322 46452 45052
rect 46396 44270 46398 44322
rect 46450 44270 46452 44322
rect 46396 44258 46452 44270
rect 46508 45106 46564 45118
rect 46508 45054 46510 45106
rect 46562 45054 46564 45106
rect 45836 44158 45838 44210
rect 45890 44158 45892 44210
rect 45836 44146 45892 44158
rect 46508 43988 46564 45054
rect 46620 44212 46676 45838
rect 46844 45220 46900 47294
rect 47180 48020 47236 48030
rect 46956 46002 47012 46014
rect 46956 45950 46958 46002
rect 47010 45950 47012 46002
rect 46956 45780 47012 45950
rect 47180 46002 47236 47964
rect 47292 46900 47348 50764
rect 47404 50754 47460 50764
rect 47740 50428 47796 51772
rect 47852 51716 47908 52780
rect 47964 52770 48020 52780
rect 49308 52276 49364 55580
rect 52332 55524 52388 55534
rect 56700 55468 56756 56030
rect 50556 54908 50820 54918
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50556 54842 50820 54852
rect 50556 53340 50820 53350
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50556 53274 50820 53284
rect 48748 52164 48804 52174
rect 48636 52162 48804 52164
rect 48636 52110 48750 52162
rect 48802 52110 48804 52162
rect 49308 52144 49364 52220
rect 50876 52276 50932 52286
rect 48636 52108 48804 52110
rect 48412 51938 48468 51950
rect 48412 51886 48414 51938
rect 48466 51886 48468 51938
rect 48412 51828 48468 51886
rect 48412 51762 48468 51772
rect 47852 51156 47908 51660
rect 48412 51492 48468 51502
rect 47964 51378 48020 51390
rect 47964 51326 47966 51378
rect 48018 51326 48020 51378
rect 47964 51268 48020 51326
rect 47964 51212 48244 51268
rect 47852 51100 48132 51156
rect 47628 50372 47796 50428
rect 48076 50484 48132 51100
rect 47516 50036 47572 50046
rect 47516 49942 47572 49980
rect 47516 49812 47572 49822
rect 47404 49700 47460 49710
rect 47404 49606 47460 49644
rect 47516 48916 47572 49756
rect 47404 48580 47460 48590
rect 47404 48242 47460 48524
rect 47404 48190 47406 48242
rect 47458 48190 47460 48242
rect 47404 48178 47460 48190
rect 47292 46844 47460 46900
rect 47292 46676 47348 46686
rect 47292 46582 47348 46620
rect 47180 45950 47182 46002
rect 47234 45950 47236 46002
rect 47180 45938 47236 45950
rect 47404 46562 47460 46844
rect 47516 46676 47572 48860
rect 47628 48692 47684 50372
rect 47852 50370 47908 50382
rect 47852 50318 47854 50370
rect 47906 50318 47908 50370
rect 47852 49812 47908 50318
rect 47852 49746 47908 49756
rect 47964 49698 48020 49710
rect 47964 49646 47966 49698
rect 48018 49646 48020 49698
rect 47740 49140 47796 49150
rect 47740 49046 47796 49084
rect 47852 49028 47908 49038
rect 47852 48934 47908 48972
rect 47684 48636 47796 48692
rect 47628 48626 47684 48636
rect 47516 46610 47572 46620
rect 47404 46510 47406 46562
rect 47458 46510 47460 46562
rect 47404 46228 47460 46510
rect 46956 45444 47012 45724
rect 46956 45388 47348 45444
rect 46844 45164 47012 45220
rect 46620 44146 46676 44156
rect 45164 43708 45444 43764
rect 46172 43932 46564 43988
rect 46732 44098 46788 44110
rect 46732 44046 46734 44098
rect 46786 44046 46788 44098
rect 44716 43652 44772 43662
rect 44716 43558 44772 43596
rect 45052 43652 45108 43662
rect 45164 43652 45220 43708
rect 45052 43650 45220 43652
rect 45052 43598 45054 43650
rect 45106 43598 45220 43650
rect 45052 43596 45220 43598
rect 45052 43586 45108 43596
rect 44828 43538 44884 43550
rect 44828 43486 44830 43538
rect 44882 43486 44884 43538
rect 44828 43204 44884 43486
rect 44940 43428 44996 43438
rect 44940 43334 44996 43372
rect 44828 43148 45108 43204
rect 44492 41860 44548 42476
rect 44828 42084 44884 42094
rect 44828 41990 44884 42028
rect 44492 41794 44548 41804
rect 44380 41074 44436 41132
rect 44380 41022 44382 41074
rect 44434 41022 44436 41074
rect 44380 41010 44436 41022
rect 44716 40964 44772 40974
rect 44716 40962 44884 40964
rect 44716 40910 44718 40962
rect 44770 40910 44884 40962
rect 44716 40908 44884 40910
rect 44716 40898 44772 40908
rect 44828 40852 44884 40908
rect 44940 40852 44996 40862
rect 44156 40796 44436 40852
rect 44828 40796 44940 40852
rect 44044 40350 44046 40402
rect 44098 40350 44100 40402
rect 44044 39842 44100 40350
rect 44044 39790 44046 39842
rect 44098 39790 44100 39842
rect 44044 39778 44100 39790
rect 44268 40402 44324 40414
rect 44268 40350 44270 40402
rect 44322 40350 44324 40402
rect 43820 39442 43876 39452
rect 44044 39508 44100 39518
rect 44044 39414 44100 39452
rect 44156 38834 44212 38846
rect 44156 38782 44158 38834
rect 44210 38782 44212 38834
rect 43596 38610 43652 38622
rect 43596 38558 43598 38610
rect 43650 38558 43652 38610
rect 43596 37826 43652 38558
rect 44044 37940 44100 37950
rect 44044 37846 44100 37884
rect 43596 37774 43598 37826
rect 43650 37774 43652 37826
rect 43596 37042 43652 37774
rect 44156 37828 44212 38782
rect 44156 37762 44212 37772
rect 44044 37604 44100 37614
rect 43932 37268 43988 37278
rect 43932 37174 43988 37212
rect 43596 36990 43598 37042
rect 43650 36990 43652 37042
rect 43596 36978 43652 36990
rect 43820 36370 43876 36382
rect 43820 36318 43822 36370
rect 43874 36318 43876 36370
rect 43708 35812 43764 35822
rect 43708 35718 43764 35756
rect 43484 35534 43486 35586
rect 43538 35534 43540 35586
rect 43484 35522 43540 35534
rect 43596 35698 43652 35710
rect 43596 35646 43598 35698
rect 43650 35646 43652 35698
rect 43372 32050 43428 32060
rect 43484 34356 43540 34366
rect 43148 31892 43204 31902
rect 43036 31780 43092 31790
rect 42812 31612 42980 31668
rect 42588 30884 42644 30894
rect 42700 30884 42756 31612
rect 42924 31218 42980 31612
rect 42924 31166 42926 31218
rect 42978 31166 42980 31218
rect 42924 31154 42980 31166
rect 43036 31218 43092 31724
rect 43036 31166 43038 31218
rect 43090 31166 43092 31218
rect 43036 31154 43092 31166
rect 43148 31778 43204 31836
rect 43148 31726 43150 31778
rect 43202 31726 43204 31778
rect 42812 31106 42868 31118
rect 42812 31054 42814 31106
rect 42866 31054 42868 31106
rect 42812 30996 42868 31054
rect 43148 31108 43204 31726
rect 43484 31780 43540 34300
rect 43596 34132 43652 35646
rect 43596 34066 43652 34076
rect 43708 35588 43764 35598
rect 43708 33348 43764 35532
rect 43820 33684 43876 36318
rect 43932 34692 43988 34702
rect 43932 34598 43988 34636
rect 43820 33618 43876 33628
rect 43932 34018 43988 34030
rect 43932 33966 43934 34018
rect 43986 33966 43988 34018
rect 43708 33292 43876 33348
rect 43708 33124 43764 33134
rect 43708 33030 43764 33068
rect 43820 32788 43876 33292
rect 43932 33124 43988 33966
rect 44044 33906 44100 37548
rect 44156 37492 44212 37502
rect 44268 37492 44324 40350
rect 44380 40292 44436 40796
rect 44716 40740 44772 40750
rect 44604 40628 44660 40638
rect 44604 40534 44660 40572
rect 44716 40626 44772 40684
rect 44716 40574 44718 40626
rect 44770 40574 44772 40626
rect 44716 40562 44772 40574
rect 44492 40516 44548 40526
rect 44492 40422 44548 40460
rect 44380 40236 44772 40292
rect 44604 39842 44660 39854
rect 44604 39790 44606 39842
rect 44658 39790 44660 39842
rect 44156 37490 44324 37492
rect 44156 37438 44158 37490
rect 44210 37438 44324 37490
rect 44156 37436 44324 37438
rect 44380 39508 44436 39518
rect 44156 37426 44212 37436
rect 44156 37266 44212 37278
rect 44156 37214 44158 37266
rect 44210 37214 44212 37266
rect 44156 37156 44212 37214
rect 44156 36372 44212 37100
rect 44156 36278 44212 36316
rect 44268 37044 44324 37054
rect 44268 34468 44324 36988
rect 44380 36036 44436 39452
rect 44492 39394 44548 39406
rect 44492 39342 44494 39394
rect 44546 39342 44548 39394
rect 44492 39060 44548 39342
rect 44492 38994 44548 39004
rect 44604 38946 44660 39790
rect 44604 38894 44606 38946
rect 44658 38894 44660 38946
rect 44604 38882 44660 38894
rect 44716 38164 44772 40236
rect 44940 38834 44996 40796
rect 44940 38782 44942 38834
rect 44994 38782 44996 38834
rect 44940 38770 44996 38782
rect 44716 38098 44772 38108
rect 44492 37828 44548 37838
rect 44548 37772 44660 37828
rect 44492 37696 44548 37772
rect 44492 37266 44548 37278
rect 44492 37214 44494 37266
rect 44546 37214 44548 37266
rect 44492 36484 44548 37214
rect 44604 37044 44660 37772
rect 44604 36978 44660 36988
rect 44940 37154 44996 37166
rect 44940 37102 44942 37154
rect 44994 37102 44996 37154
rect 44492 36418 44548 36428
rect 44604 36372 44660 36382
rect 44604 36260 44660 36316
rect 44380 35970 44436 35980
rect 44492 36258 44660 36260
rect 44492 36206 44606 36258
rect 44658 36206 44660 36258
rect 44492 36204 44660 36206
rect 44492 35588 44548 36204
rect 44604 36194 44660 36204
rect 44604 35812 44660 35822
rect 44604 35718 44660 35756
rect 44492 35522 44548 35532
rect 44940 35476 44996 37102
rect 45052 36708 45108 43148
rect 45164 42308 45220 43596
rect 46172 43652 46228 43932
rect 46620 43876 46676 43886
rect 46284 43764 46340 43774
rect 46284 43762 46452 43764
rect 46284 43710 46286 43762
rect 46338 43710 46452 43762
rect 46284 43708 46452 43710
rect 46284 43698 46340 43708
rect 45276 43540 45332 43550
rect 45276 43446 45332 43484
rect 45836 43540 45892 43550
rect 45836 43446 45892 43484
rect 46172 43538 46228 43596
rect 46172 43486 46174 43538
rect 46226 43486 46228 43538
rect 46172 43474 46228 43486
rect 46284 43316 46340 43326
rect 45836 43314 46340 43316
rect 45836 43262 46286 43314
rect 46338 43262 46340 43314
rect 45836 43260 46340 43262
rect 45724 42980 45780 42990
rect 45724 42886 45780 42924
rect 45164 42242 45220 42252
rect 45388 42420 45444 42430
rect 45276 42196 45332 42206
rect 45276 42102 45332 42140
rect 45164 41860 45220 41870
rect 45164 40626 45220 41804
rect 45388 41636 45444 42364
rect 45388 41570 45444 41580
rect 45612 41412 45668 41422
rect 45388 41076 45444 41086
rect 45388 40982 45444 41020
rect 45164 40574 45166 40626
rect 45218 40574 45220 40626
rect 45164 40562 45220 40574
rect 45612 40626 45668 41356
rect 45612 40574 45614 40626
rect 45666 40574 45668 40626
rect 45612 40562 45668 40574
rect 45276 39396 45332 39406
rect 45276 37268 45332 39340
rect 45500 39396 45556 39406
rect 45500 39302 45556 39340
rect 45724 38948 45780 38958
rect 45500 38722 45556 38734
rect 45500 38670 45502 38722
rect 45554 38670 45556 38722
rect 45500 38668 45556 38670
rect 45500 38612 45668 38668
rect 45612 38500 45668 38612
rect 45500 37940 45556 37950
rect 45500 37846 45556 37884
rect 45612 37826 45668 38444
rect 45724 38610 45780 38892
rect 45724 38558 45726 38610
rect 45778 38558 45780 38610
rect 45724 37940 45780 38558
rect 45836 38050 45892 43260
rect 46284 43250 46340 43260
rect 46284 42980 46340 42990
rect 46396 42980 46452 43708
rect 46620 43540 46676 43820
rect 46620 43408 46676 43484
rect 46732 42980 46788 44046
rect 46284 42978 46676 42980
rect 46284 42926 46286 42978
rect 46338 42926 46676 42978
rect 46284 42924 46676 42926
rect 46284 42914 46340 42924
rect 45948 42756 46004 42766
rect 46508 42756 46564 42766
rect 45948 42662 46004 42700
rect 46396 42754 46564 42756
rect 46396 42702 46510 42754
rect 46562 42702 46564 42754
rect 46396 42700 46564 42702
rect 46060 42644 46116 42654
rect 46060 42550 46116 42588
rect 45948 41972 46004 41982
rect 45948 41878 46004 41916
rect 46396 41748 46452 42700
rect 46508 42690 46564 42700
rect 46620 41970 46676 42924
rect 46732 42914 46788 42924
rect 46844 43652 46900 43662
rect 46620 41918 46622 41970
rect 46674 41918 46676 41970
rect 46620 41906 46676 41918
rect 46844 42756 46900 43596
rect 46844 41970 46900 42700
rect 46844 41918 46846 41970
rect 46898 41918 46900 41970
rect 46844 41906 46900 41918
rect 46172 41746 46452 41748
rect 46172 41694 46398 41746
rect 46450 41694 46452 41746
rect 46172 41692 46452 41694
rect 46060 40740 46116 40750
rect 46060 39618 46116 40684
rect 46172 39730 46228 41692
rect 46396 41682 46452 41692
rect 46508 41186 46564 41198
rect 46508 41134 46510 41186
rect 46562 41134 46564 41186
rect 46284 41074 46340 41086
rect 46284 41022 46286 41074
rect 46338 41022 46340 41074
rect 46284 40740 46340 41022
rect 46396 40964 46452 40974
rect 46396 40870 46452 40908
rect 46284 40674 46340 40684
rect 46508 40516 46564 41134
rect 46844 41076 46900 41086
rect 46844 40982 46900 41020
rect 46732 40964 46788 40974
rect 46172 39678 46174 39730
rect 46226 39678 46228 39730
rect 46172 39666 46228 39678
rect 46396 40460 46564 40516
rect 46620 40516 46676 40526
rect 46396 40404 46452 40460
rect 46060 39566 46062 39618
rect 46114 39566 46116 39618
rect 46060 39554 46116 39566
rect 46396 39618 46452 40348
rect 46620 40402 46676 40460
rect 46620 40350 46622 40402
rect 46674 40350 46676 40402
rect 46620 40338 46676 40350
rect 46396 39566 46398 39618
rect 46450 39566 46452 39618
rect 46396 39554 46452 39566
rect 46508 39618 46564 39630
rect 46508 39566 46510 39618
rect 46562 39566 46564 39618
rect 46508 39172 46564 39566
rect 46732 39618 46788 40908
rect 46844 40740 46900 40750
rect 46844 40290 46900 40684
rect 46956 40514 47012 45164
rect 47180 44324 47236 44334
rect 47180 44230 47236 44268
rect 47292 43650 47348 45388
rect 47404 44546 47460 46172
rect 47516 45890 47572 45902
rect 47516 45838 47518 45890
rect 47570 45838 47572 45890
rect 47516 45330 47572 45838
rect 47516 45278 47518 45330
rect 47570 45278 47572 45330
rect 47516 45266 47572 45278
rect 47404 44494 47406 44546
rect 47458 44494 47460 44546
rect 47404 43876 47460 44494
rect 47628 44322 47684 44334
rect 47628 44270 47630 44322
rect 47682 44270 47684 44322
rect 47404 43810 47460 43820
rect 47516 44212 47572 44222
rect 47516 43652 47572 44156
rect 47292 43598 47294 43650
rect 47346 43598 47348 43650
rect 47292 43586 47348 43598
rect 47404 43650 47572 43652
rect 47404 43598 47518 43650
rect 47570 43598 47572 43650
rect 47404 43596 47572 43598
rect 47068 42978 47124 42990
rect 47068 42926 47070 42978
rect 47122 42926 47124 42978
rect 47068 42866 47124 42926
rect 47068 42814 47070 42866
rect 47122 42814 47124 42866
rect 47068 41300 47124 42814
rect 47068 41234 47124 41244
rect 47404 40964 47460 43596
rect 47516 43586 47572 43596
rect 47628 43426 47684 44270
rect 47628 43374 47630 43426
rect 47682 43374 47684 43426
rect 47628 43362 47684 43374
rect 47740 42978 47796 48636
rect 47852 48244 47908 48254
rect 47852 48150 47908 48188
rect 47852 47908 47908 47918
rect 47964 47908 48020 49646
rect 48076 49250 48132 50428
rect 48188 50428 48244 51212
rect 48300 50818 48356 50830
rect 48300 50766 48302 50818
rect 48354 50766 48356 50818
rect 48300 50706 48356 50766
rect 48300 50654 48302 50706
rect 48354 50654 48356 50706
rect 48300 50642 48356 50654
rect 48188 50372 48356 50428
rect 48076 49198 48078 49250
rect 48130 49198 48132 49250
rect 48076 49186 48132 49198
rect 48188 49252 48244 49262
rect 48188 49158 48244 49196
rect 48076 48804 48132 48814
rect 48076 48466 48132 48748
rect 48076 48414 48078 48466
rect 48130 48414 48132 48466
rect 48076 48402 48132 48414
rect 48188 48244 48244 48254
rect 48188 48150 48244 48188
rect 47908 47852 48020 47908
rect 47852 47458 47908 47852
rect 47852 47406 47854 47458
rect 47906 47406 47908 47458
rect 47852 47394 47908 47406
rect 48300 46898 48356 50372
rect 48412 48356 48468 51436
rect 48636 50372 48692 52108
rect 48748 52098 48804 52108
rect 49196 52052 49252 52062
rect 48748 51266 48804 51278
rect 48748 51214 48750 51266
rect 48802 51214 48804 51266
rect 48748 50428 48804 51214
rect 49196 50818 49252 51996
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 49868 51604 49924 51614
rect 49868 51510 49924 51548
rect 49532 51380 49588 51390
rect 49196 50766 49198 50818
rect 49250 50766 49252 50818
rect 49196 50754 49252 50766
rect 49420 51378 49588 51380
rect 49420 51326 49534 51378
rect 49586 51326 49588 51378
rect 49420 51324 49588 51326
rect 48748 50372 49028 50428
rect 48524 50370 48692 50372
rect 48524 50318 48638 50370
rect 48690 50318 48692 50370
rect 48524 50316 48692 50318
rect 48524 49700 48580 50316
rect 48636 50306 48692 50316
rect 48524 49634 48580 49644
rect 48636 49698 48692 49710
rect 48636 49646 48638 49698
rect 48690 49646 48692 49698
rect 48636 49364 48692 49646
rect 48692 49308 48804 49364
rect 48636 49298 48692 49308
rect 48636 48916 48692 48926
rect 48636 48822 48692 48860
rect 48636 48356 48692 48366
rect 48412 48354 48692 48356
rect 48412 48302 48638 48354
rect 48690 48302 48692 48354
rect 48412 48300 48692 48302
rect 48300 46846 48302 46898
rect 48354 46846 48356 46898
rect 48300 46834 48356 46846
rect 48076 46674 48132 46686
rect 48076 46622 48078 46674
rect 48130 46622 48132 46674
rect 47964 45778 48020 45790
rect 47964 45726 47966 45778
rect 48018 45726 48020 45778
rect 47852 45668 47908 45678
rect 47852 44884 47908 45612
rect 47964 45556 48020 45726
rect 48076 45780 48132 46622
rect 48412 46676 48468 46686
rect 48412 46582 48468 46620
rect 48412 45892 48468 45902
rect 48412 45798 48468 45836
rect 48076 45714 48132 45724
rect 48524 45556 48580 48300
rect 48636 48290 48692 48300
rect 47964 45500 48580 45556
rect 48748 46004 48804 49308
rect 48860 48804 48916 48814
rect 48860 47458 48916 48748
rect 48972 48468 49028 50372
rect 49420 50036 49476 51324
rect 49532 51314 49588 51324
rect 49756 51378 49812 51390
rect 49756 51326 49758 51378
rect 49810 51326 49812 51378
rect 49532 50932 49588 50942
rect 49532 50818 49588 50876
rect 49532 50766 49534 50818
rect 49586 50766 49588 50818
rect 49532 50754 49588 50766
rect 49420 49970 49476 49980
rect 49756 50482 49812 51326
rect 50204 51378 50260 51390
rect 50204 51326 50206 51378
rect 50258 51326 50260 51378
rect 50204 50932 50260 51326
rect 50764 51268 50820 51278
rect 50204 50820 50260 50876
rect 50428 51266 50820 51268
rect 50428 51214 50766 51266
rect 50818 51214 50820 51266
rect 50428 51212 50820 51214
rect 50316 50820 50372 50830
rect 50204 50818 50372 50820
rect 50204 50766 50318 50818
rect 50370 50766 50372 50818
rect 50204 50764 50372 50766
rect 50316 50754 50372 50764
rect 50428 50706 50484 51212
rect 50764 50818 50820 51212
rect 50764 50766 50766 50818
rect 50818 50766 50820 50818
rect 50764 50754 50820 50766
rect 50428 50654 50430 50706
rect 50482 50654 50484 50706
rect 50428 50642 50484 50654
rect 50876 50706 50932 52220
rect 50876 50654 50878 50706
rect 50930 50654 50932 50706
rect 49756 50430 49758 50482
rect 49810 50430 49812 50482
rect 49756 50036 49812 50430
rect 50876 50428 50932 50654
rect 49756 49970 49812 49980
rect 50428 50372 50932 50428
rect 51324 50818 51380 50830
rect 51324 50766 51326 50818
rect 51378 50766 51380 50818
rect 51324 50706 51380 50766
rect 51324 50654 51326 50706
rect 51378 50654 51380 50706
rect 49532 49698 49588 49710
rect 49532 49646 49534 49698
rect 49586 49646 49588 49698
rect 48972 48402 49028 48412
rect 49420 49586 49476 49598
rect 49420 49534 49422 49586
rect 49474 49534 49476 49586
rect 48860 47406 48862 47458
rect 48914 47406 48916 47458
rect 48860 47394 48916 47406
rect 49308 46564 49364 46574
rect 48972 46340 49028 46350
rect 48860 46004 48916 46014
rect 48748 46002 48916 46004
rect 48748 45950 48862 46002
rect 48914 45950 48916 46002
rect 48748 45948 48916 45950
rect 48076 45220 48132 45230
rect 48076 45126 48132 45164
rect 47964 45108 48020 45118
rect 47964 45014 48020 45052
rect 48188 45106 48244 45118
rect 48188 45054 48190 45106
rect 48242 45054 48244 45106
rect 48188 44884 48244 45054
rect 47852 44828 48244 44884
rect 47852 44434 47908 44828
rect 47852 44382 47854 44434
rect 47906 44382 47908 44434
rect 47852 44370 47908 44382
rect 48300 43876 48356 45500
rect 48748 45220 48804 45948
rect 48860 45938 48916 45948
rect 48636 45164 48748 45220
rect 48636 44322 48692 45164
rect 48748 45154 48804 45164
rect 48972 45892 49028 46284
rect 48748 44996 48804 45006
rect 48972 44996 49028 45836
rect 48748 44994 49028 44996
rect 48748 44942 48750 44994
rect 48802 44942 49028 44994
rect 48748 44940 49028 44942
rect 49084 45108 49140 45118
rect 48748 44930 48804 44940
rect 48636 44270 48638 44322
rect 48690 44270 48692 44322
rect 48412 44212 48468 44222
rect 48412 44118 48468 44156
rect 47740 42926 47742 42978
rect 47794 42926 47796 42978
rect 47516 42532 47572 42542
rect 47516 42438 47572 42476
rect 47628 42084 47684 42094
rect 47404 40898 47460 40908
rect 47516 42082 47684 42084
rect 47516 42030 47630 42082
rect 47682 42030 47684 42082
rect 47516 42028 47684 42030
rect 46956 40462 46958 40514
rect 47010 40462 47012 40514
rect 46956 40450 47012 40462
rect 47516 40852 47572 42028
rect 47628 42018 47684 42028
rect 47740 41858 47796 42926
rect 47852 43820 48356 43876
rect 47852 42866 47908 43820
rect 48636 43764 48692 44270
rect 48860 44324 48916 44334
rect 48860 44230 48916 44268
rect 49084 44322 49140 45052
rect 49084 44270 49086 44322
rect 49138 44270 49140 44322
rect 48636 43698 48692 43708
rect 48076 43652 48132 43662
rect 48076 43558 48132 43596
rect 48412 43652 48468 43662
rect 47852 42814 47854 42866
rect 47906 42814 47908 42866
rect 47852 42802 47908 42814
rect 48188 43428 48244 43438
rect 48076 42530 48132 42542
rect 48076 42478 48078 42530
rect 48130 42478 48132 42530
rect 47740 41806 47742 41858
rect 47794 41806 47796 41858
rect 47740 41300 47796 41806
rect 47740 41234 47796 41244
rect 47852 42084 47908 42094
rect 46844 40238 46846 40290
rect 46898 40238 46900 40290
rect 46844 40226 46900 40238
rect 47404 40404 47460 40414
rect 46732 39566 46734 39618
rect 46786 39566 46788 39618
rect 46732 39554 46788 39566
rect 46060 39116 46564 39172
rect 46620 39396 46676 39406
rect 46060 39058 46116 39116
rect 46060 39006 46062 39058
rect 46114 39006 46116 39058
rect 46060 38994 46116 39006
rect 46508 38948 46564 38958
rect 46620 38948 46676 39340
rect 46564 38892 46676 38948
rect 47292 38948 47348 38958
rect 46508 38816 46564 38892
rect 47068 38722 47124 38734
rect 47068 38670 47070 38722
rect 47122 38670 47124 38722
rect 47068 38500 47124 38670
rect 47068 38434 47124 38444
rect 45836 37998 45838 38050
rect 45890 37998 45892 38050
rect 45836 37986 45892 37998
rect 45724 37874 45780 37884
rect 46172 37828 46228 37838
rect 45612 37774 45614 37826
rect 45666 37774 45668 37826
rect 45612 37716 45668 37774
rect 45612 37650 45668 37660
rect 46060 37826 46228 37828
rect 46060 37774 46174 37826
rect 46226 37774 46228 37826
rect 46060 37772 46228 37774
rect 45276 37202 45332 37212
rect 46060 37492 46116 37772
rect 46172 37762 46228 37772
rect 46620 37826 46676 37838
rect 46620 37774 46622 37826
rect 46674 37774 46676 37826
rect 45500 37156 45556 37166
rect 45948 37156 46004 37166
rect 45052 36642 45108 36652
rect 45388 37154 46004 37156
rect 45388 37102 45502 37154
rect 45554 37102 45950 37154
rect 46002 37102 46004 37154
rect 45388 37100 46004 37102
rect 45276 36484 45332 36494
rect 45164 36260 45220 36270
rect 45164 35812 45220 36204
rect 45164 35698 45220 35756
rect 45164 35646 45166 35698
rect 45218 35646 45220 35698
rect 45164 35634 45220 35646
rect 44940 35420 45220 35476
rect 44380 34804 44436 34814
rect 44380 34710 44436 34748
rect 44828 34692 44884 34702
rect 44716 34690 44884 34692
rect 44716 34638 44830 34690
rect 44882 34638 44884 34690
rect 44716 34636 44884 34638
rect 44268 34412 44436 34468
rect 44044 33854 44046 33906
rect 44098 33854 44100 33906
rect 44044 33842 44100 33854
rect 44268 34130 44324 34142
rect 44268 34078 44270 34130
rect 44322 34078 44324 34130
rect 44268 33908 44324 34078
rect 44268 33842 44324 33852
rect 44156 33348 44212 33358
rect 44156 33254 44212 33292
rect 43932 33068 44212 33124
rect 43820 32732 43988 32788
rect 43484 31714 43540 31724
rect 43596 32562 43652 32574
rect 43820 32564 43876 32574
rect 43596 32510 43598 32562
rect 43650 32510 43652 32562
rect 43148 31042 43204 31052
rect 43260 31556 43316 31566
rect 43036 30996 43092 31006
rect 42812 30940 43036 30996
rect 43036 30930 43092 30940
rect 43148 30884 43204 30894
rect 42700 30828 42868 30884
rect 42588 30790 42644 30828
rect 42476 30258 42532 30268
rect 42364 30098 42420 30110
rect 42364 30046 42366 30098
rect 42418 30046 42420 30098
rect 42364 29540 42420 30046
rect 42588 30098 42644 30110
rect 42588 30046 42590 30098
rect 42642 30046 42644 30098
rect 42588 29988 42644 30046
rect 42588 29922 42644 29932
rect 42364 29474 42420 29484
rect 42812 29540 42868 30828
rect 42364 29316 42420 29326
rect 42364 29314 42756 29316
rect 42364 29262 42366 29314
rect 42418 29262 42756 29314
rect 42364 29260 42756 29262
rect 42364 29250 42420 29260
rect 42700 29204 42756 29260
rect 42700 29138 42756 29148
rect 42252 28018 42308 28028
rect 42364 29092 42420 29102
rect 42140 27746 42196 27758
rect 42140 27694 42142 27746
rect 42194 27694 42196 27746
rect 42140 27076 42196 27694
rect 42252 27748 42308 27758
rect 42252 27186 42308 27692
rect 42252 27134 42254 27186
rect 42306 27134 42308 27186
rect 42252 27122 42308 27134
rect 42140 27010 42196 27020
rect 41916 26852 42084 26908
rect 42364 26908 42420 29036
rect 42812 29092 42868 29484
rect 42812 29026 42868 29036
rect 42924 30660 42980 30670
rect 42924 28868 42980 30604
rect 43036 29986 43092 29998
rect 43036 29934 43038 29986
rect 43090 29934 43092 29986
rect 43036 29876 43092 29934
rect 43036 29810 43092 29820
rect 42588 28812 42980 28868
rect 42364 26852 42532 26908
rect 41804 26404 41860 26414
rect 41804 26290 41860 26348
rect 41804 26238 41806 26290
rect 41858 26238 41860 26290
rect 41804 26226 41860 26238
rect 41916 25620 41972 26852
rect 42140 26740 42196 26750
rect 41804 25618 41972 25620
rect 41804 25566 41918 25618
rect 41970 25566 41972 25618
rect 41804 25564 41972 25566
rect 41804 24388 41860 25564
rect 41916 25554 41972 25564
rect 42028 26068 42084 26078
rect 41916 24610 41972 24622
rect 41916 24558 41918 24610
rect 41970 24558 41972 24610
rect 41916 24500 41972 24558
rect 41916 24434 41972 24444
rect 41804 24322 41860 24332
rect 41244 23998 41246 24050
rect 41298 23998 41300 24050
rect 41244 23986 41300 23998
rect 41580 24220 41748 24276
rect 41468 23828 41524 23838
rect 41020 22482 41412 22484
rect 41020 22430 41022 22482
rect 41074 22430 41412 22482
rect 41020 22428 41412 22430
rect 41020 22418 41076 22428
rect 40908 22306 40964 22316
rect 40460 21026 40852 21028
rect 40460 20974 40462 21026
rect 40514 20974 40852 21026
rect 40460 20972 40852 20974
rect 41132 22260 41188 22270
rect 41356 22260 41412 22428
rect 41468 22482 41524 23772
rect 41580 23548 41636 24220
rect 42028 24162 42084 26012
rect 42140 26066 42196 26684
rect 42140 26014 42142 26066
rect 42194 26014 42196 26066
rect 42140 25844 42196 26014
rect 42140 25778 42196 25788
rect 42364 26628 42420 26638
rect 42364 26068 42420 26572
rect 42364 25284 42420 26012
rect 42364 25218 42420 25228
rect 42364 24388 42420 24398
rect 42028 24110 42030 24162
rect 42082 24110 42084 24162
rect 41692 24052 41748 24062
rect 41692 23958 41748 23996
rect 42028 24050 42084 24110
rect 42028 23998 42030 24050
rect 42082 23998 42084 24050
rect 42028 23986 42084 23998
rect 42140 24164 42196 24174
rect 41580 23492 41972 23548
rect 41692 23268 41748 23278
rect 41692 23266 41860 23268
rect 41692 23214 41694 23266
rect 41746 23214 41860 23266
rect 41692 23212 41860 23214
rect 41692 23202 41748 23212
rect 41580 23156 41636 23166
rect 41580 23042 41636 23100
rect 41580 22990 41582 23042
rect 41634 22990 41636 23042
rect 41580 22978 41636 22990
rect 41468 22430 41470 22482
rect 41522 22430 41524 22482
rect 41468 22418 41524 22430
rect 41356 22204 41636 22260
rect 40460 20962 40516 20972
rect 40348 20580 40404 20590
rect 40348 20356 40404 20524
rect 40348 20290 40404 20300
rect 40796 20580 40852 20590
rect 40796 20244 40852 20524
rect 40572 19908 40628 19918
rect 40572 19814 40628 19852
rect 40236 18834 40292 18844
rect 40348 19124 40404 19134
rect 40460 19124 40516 19134
rect 40404 19122 40516 19124
rect 40404 19070 40462 19122
rect 40514 19070 40516 19122
rect 40404 19068 40516 19070
rect 40124 18450 40180 18462
rect 40124 18398 40126 18450
rect 40178 18398 40180 18450
rect 40012 16996 40068 17006
rect 40012 16882 40068 16940
rect 40012 16830 40014 16882
rect 40066 16830 40068 16882
rect 40012 16818 40068 16830
rect 40124 16884 40180 18398
rect 40348 18116 40404 19068
rect 40460 19058 40516 19068
rect 40796 19122 40852 20188
rect 40796 19070 40798 19122
rect 40850 19070 40852 19122
rect 40796 19058 40852 19070
rect 40684 18900 40740 18910
rect 40684 18674 40740 18844
rect 40684 18622 40686 18674
rect 40738 18622 40740 18674
rect 40684 18610 40740 18622
rect 40572 18564 40628 18574
rect 40572 18470 40628 18508
rect 40796 18564 40852 18574
rect 41020 18564 41076 18574
rect 40796 18562 41076 18564
rect 40796 18510 40798 18562
rect 40850 18510 41022 18562
rect 41074 18510 41076 18562
rect 40796 18508 41076 18510
rect 40796 18498 40852 18508
rect 41020 18498 41076 18508
rect 41020 18338 41076 18350
rect 41020 18286 41022 18338
rect 41074 18286 41076 18338
rect 40348 18060 40516 18116
rect 40348 17892 40404 17902
rect 40348 17108 40404 17836
rect 40348 17042 40404 17052
rect 39900 16604 40068 16660
rect 39116 16100 39172 16110
rect 39004 16098 39172 16100
rect 39004 16046 39118 16098
rect 39170 16046 39172 16098
rect 39004 16044 39172 16046
rect 38556 15474 38612 15484
rect 38668 15764 38724 15774
rect 38668 15538 38724 15708
rect 38668 15486 38670 15538
rect 38722 15486 38724 15538
rect 38220 13918 38222 13970
rect 38274 13918 38276 13970
rect 38220 13906 38276 13918
rect 38332 15092 38500 15148
rect 37548 13806 37550 13858
rect 37602 13806 37604 13858
rect 37548 13794 37604 13806
rect 37772 13636 37828 13646
rect 37548 13522 37604 13534
rect 37548 13470 37550 13522
rect 37602 13470 37604 13522
rect 37548 12402 37604 13470
rect 37772 12962 37828 13580
rect 38332 13188 38388 15092
rect 38668 14868 38724 15486
rect 38668 14802 38724 14812
rect 38892 14756 38948 14766
rect 38444 14644 38500 14654
rect 38444 14550 38500 14588
rect 38668 14532 38724 14542
rect 38668 13746 38724 14476
rect 38668 13694 38670 13746
rect 38722 13694 38724 13746
rect 38668 13524 38724 13694
rect 38892 13746 38948 14700
rect 39004 14420 39060 14458
rect 39004 14354 39060 14364
rect 38892 13694 38894 13746
rect 38946 13694 38948 13746
rect 38780 13636 38836 13646
rect 38780 13542 38836 13580
rect 38668 13458 38724 13468
rect 37772 12910 37774 12962
rect 37826 12910 37828 12962
rect 37772 12898 37828 12910
rect 37884 13132 38388 13188
rect 38556 13412 38612 13422
rect 37548 12350 37550 12402
rect 37602 12350 37604 12402
rect 37548 12338 37604 12350
rect 37772 11508 37828 11518
rect 37772 11414 37828 11452
rect 37212 7746 37268 7756
rect 37324 9660 37492 9716
rect 37660 10498 37716 10510
rect 37660 10446 37662 10498
rect 37714 10446 37716 10498
rect 37324 3892 37380 9660
rect 37548 9604 37604 9614
rect 37660 9604 37716 10446
rect 37436 9602 37716 9604
rect 37436 9550 37550 9602
rect 37602 9550 37716 9602
rect 37436 9548 37716 9550
rect 37436 9042 37492 9548
rect 37548 9538 37604 9548
rect 37436 8990 37438 9042
rect 37490 8990 37492 9042
rect 37436 8932 37492 8990
rect 37772 9044 37828 9054
rect 37772 8950 37828 8988
rect 37436 8036 37492 8876
rect 37660 8036 37716 8046
rect 37436 8034 37716 8036
rect 37436 7982 37662 8034
rect 37714 7982 37716 8034
rect 37436 7980 37716 7982
rect 37660 6468 37716 7980
rect 37772 6692 37828 6702
rect 37772 6468 37828 6636
rect 37660 6466 37828 6468
rect 37660 6414 37774 6466
rect 37826 6414 37828 6466
rect 37660 6412 37828 6414
rect 37436 5908 37492 5918
rect 37660 5908 37716 6412
rect 37772 6402 37828 6412
rect 37436 5906 37716 5908
rect 37436 5854 37438 5906
rect 37490 5854 37716 5906
rect 37436 5852 37716 5854
rect 37772 6132 37828 6142
rect 37772 5906 37828 6076
rect 37772 5854 37774 5906
rect 37826 5854 37828 5906
rect 37436 5124 37492 5852
rect 37772 5842 37828 5854
rect 37436 5030 37492 5068
rect 37324 3826 37380 3836
rect 37660 3332 37716 3342
rect 37660 3238 37716 3276
rect 37100 2818 37156 2828
rect 37884 1540 37940 13132
rect 38556 13076 38612 13356
rect 38332 13074 38612 13076
rect 38332 13022 38558 13074
rect 38610 13022 38612 13074
rect 38332 13020 38612 13022
rect 37996 12740 38052 12750
rect 37996 12738 38276 12740
rect 37996 12686 37998 12738
rect 38050 12686 38276 12738
rect 37996 12684 38276 12686
rect 37996 12674 38052 12684
rect 37996 11396 38052 11406
rect 37996 10500 38052 11340
rect 37996 10434 38052 10444
rect 38108 11394 38164 11406
rect 38108 11342 38110 11394
rect 38162 11342 38164 11394
rect 38108 9828 38164 11342
rect 38220 10724 38276 12684
rect 38332 12402 38388 13020
rect 38556 13010 38612 13020
rect 38332 12350 38334 12402
rect 38386 12350 38388 12402
rect 38332 12338 38388 12350
rect 38668 12628 38724 12638
rect 38668 12402 38724 12572
rect 38668 12350 38670 12402
rect 38722 12350 38724 12402
rect 38668 12338 38724 12350
rect 38780 11844 38836 11854
rect 38668 11396 38724 11406
rect 38668 11302 38724 11340
rect 38668 10836 38724 10846
rect 38780 10836 38836 11788
rect 38892 11508 38948 13694
rect 38892 11442 38948 11452
rect 39004 14196 39060 14206
rect 38668 10834 38836 10836
rect 38668 10782 38670 10834
rect 38722 10782 38836 10834
rect 38668 10780 38836 10782
rect 39004 10836 39060 14140
rect 39116 13412 39172 16044
rect 39228 15540 39284 15550
rect 39228 15446 39284 15484
rect 39340 15148 39396 16268
rect 39452 16268 39676 16324
rect 39452 15986 39508 16268
rect 39676 16258 39732 16268
rect 39452 15934 39454 15986
rect 39506 15934 39508 15986
rect 39452 15922 39508 15934
rect 39900 15876 39956 15886
rect 39900 15782 39956 15820
rect 39564 15540 39620 15550
rect 39564 15446 39620 15484
rect 40012 15538 40068 16604
rect 40012 15486 40014 15538
rect 40066 15486 40068 15538
rect 40012 15474 40068 15486
rect 40124 15148 40180 16828
rect 40236 16996 40292 17006
rect 40236 16660 40292 16940
rect 40348 16884 40404 16894
rect 40348 16790 40404 16828
rect 40236 16604 40404 16660
rect 39116 13346 39172 13356
rect 39228 15092 39396 15148
rect 40012 15092 40180 15148
rect 39116 12964 39172 12974
rect 39116 11844 39172 12908
rect 39228 12402 39284 15092
rect 39788 14644 39844 14654
rect 39788 14550 39844 14588
rect 39340 14306 39396 14318
rect 39340 14254 39342 14306
rect 39394 14254 39396 14306
rect 39340 14196 39396 14254
rect 39340 14130 39396 14140
rect 39340 13748 39396 13758
rect 39340 13746 39956 13748
rect 39340 13694 39342 13746
rect 39394 13694 39956 13746
rect 39340 13692 39956 13694
rect 39340 13682 39396 13692
rect 39788 13524 39844 13534
rect 39676 13412 39732 13422
rect 39676 13076 39732 13356
rect 39676 13010 39732 13020
rect 39228 12350 39230 12402
rect 39282 12350 39284 12402
rect 39228 12338 39284 12350
rect 39452 12852 39508 12862
rect 39116 11778 39172 11788
rect 39452 11844 39508 12796
rect 39452 11778 39508 11788
rect 39116 10836 39172 10846
rect 39004 10834 39172 10836
rect 39004 10782 39118 10834
rect 39170 10782 39172 10834
rect 39004 10780 39172 10782
rect 38668 10770 38724 10780
rect 39116 10770 39172 10780
rect 38220 10668 38500 10724
rect 38220 10500 38276 10510
rect 38220 10406 38276 10444
rect 38220 9828 38276 9838
rect 38108 9826 38276 9828
rect 38108 9774 38222 9826
rect 38274 9774 38276 9826
rect 38108 9772 38276 9774
rect 38220 8258 38276 9772
rect 38220 8206 38222 8258
rect 38274 8206 38276 8258
rect 37996 7700 38052 7710
rect 37996 7606 38052 7644
rect 38220 6692 38276 8206
rect 38332 8260 38388 8270
rect 38332 7698 38388 8204
rect 38332 7646 38334 7698
rect 38386 7646 38388 7698
rect 38332 7364 38388 7646
rect 38332 7298 38388 7308
rect 38220 6598 38276 6636
rect 38444 6692 38500 10668
rect 39452 10500 39508 10510
rect 39452 10406 39508 10444
rect 39788 10500 39844 13468
rect 39900 12962 39956 13692
rect 39900 12910 39902 12962
rect 39954 12910 39956 12962
rect 39900 12898 39956 12910
rect 40012 12402 40068 15092
rect 40124 14196 40180 14206
rect 40124 13970 40180 14140
rect 40124 13918 40126 13970
rect 40178 13918 40180 13970
rect 40124 13906 40180 13918
rect 40348 13970 40404 16604
rect 40460 16548 40516 18060
rect 40796 17780 40852 17790
rect 40796 17686 40852 17724
rect 41020 17778 41076 18286
rect 41020 17726 41022 17778
rect 41074 17726 41076 17778
rect 41020 17714 41076 17726
rect 40572 17666 40628 17678
rect 40572 17614 40574 17666
rect 40626 17614 40628 17666
rect 40572 16772 40628 17614
rect 41020 17556 41076 17566
rect 41020 17462 41076 17500
rect 40572 16706 40628 16716
rect 41020 16884 41076 16894
rect 40572 16548 40628 16558
rect 40460 16492 40572 16548
rect 40460 16324 40516 16334
rect 40460 15316 40516 16268
rect 40460 15250 40516 15260
rect 40460 14532 40516 14542
rect 40460 14438 40516 14476
rect 40348 13918 40350 13970
rect 40402 13918 40404 13970
rect 40236 13634 40292 13646
rect 40236 13582 40238 13634
rect 40290 13582 40292 13634
rect 40236 13188 40292 13582
rect 40348 13524 40404 13918
rect 40572 13860 40628 16492
rect 40908 16324 40964 16362
rect 40908 16258 40964 16268
rect 41020 16322 41076 16828
rect 41020 16270 41022 16322
rect 41074 16270 41076 16322
rect 41020 15988 41076 16270
rect 40684 15540 40740 15578
rect 40684 15474 40740 15484
rect 40348 13458 40404 13468
rect 40460 13804 40628 13860
rect 40684 15316 40740 15326
rect 40236 13132 40404 13188
rect 40236 12964 40292 12974
rect 40236 12870 40292 12908
rect 40124 12740 40180 12750
rect 40348 12740 40404 13132
rect 40124 12646 40180 12684
rect 40236 12684 40404 12740
rect 40012 12350 40014 12402
rect 40066 12350 40068 12402
rect 40012 12338 40068 12350
rect 40124 11844 40180 11854
rect 40124 10834 40180 11788
rect 40124 10782 40126 10834
rect 40178 10782 40180 10834
rect 40124 10770 40180 10782
rect 39788 10434 39844 10444
rect 38668 9828 38724 9838
rect 38668 9734 38724 9772
rect 39116 8596 39172 8606
rect 38668 8258 38724 8270
rect 38668 8206 38670 8258
rect 38722 8206 38724 8258
rect 38668 7700 38724 8206
rect 38668 7634 38724 7644
rect 39116 7698 39172 8540
rect 39116 7646 39118 7698
rect 39170 7646 39172 7698
rect 39116 7634 39172 7646
rect 39564 8260 39620 8270
rect 39564 7812 39620 8204
rect 39564 7698 39620 7756
rect 39564 7646 39566 7698
rect 39618 7646 39620 7698
rect 39564 7634 39620 7646
rect 38444 6626 38500 6636
rect 38780 7364 38836 7374
rect 38780 6690 38836 7308
rect 40012 7364 40068 7374
rect 40012 7270 40068 7308
rect 38780 6638 38782 6690
rect 38834 6638 38836 6690
rect 38780 6626 38836 6638
rect 40236 5908 40292 12684
rect 40460 12404 40516 13804
rect 40572 13634 40628 13646
rect 40572 13582 40574 13634
rect 40626 13582 40628 13634
rect 40572 13412 40628 13582
rect 40572 13346 40628 13356
rect 40572 12404 40628 12414
rect 40460 12348 40572 12404
rect 40572 12272 40628 12348
rect 40572 10836 40628 10846
rect 40684 10836 40740 15260
rect 41020 15148 41076 15932
rect 41132 16772 41188 22204
rect 41468 21924 41524 21934
rect 41468 21810 41524 21868
rect 41468 21758 41470 21810
rect 41522 21758 41524 21810
rect 41468 21746 41524 21758
rect 41468 21362 41524 21374
rect 41468 21310 41470 21362
rect 41522 21310 41524 21362
rect 41468 21026 41524 21310
rect 41468 20974 41470 21026
rect 41522 20974 41524 21026
rect 41468 20962 41524 20974
rect 41244 20804 41300 20814
rect 41244 20710 41300 20748
rect 41580 20130 41636 22204
rect 41804 21588 41860 23212
rect 41916 23266 41972 23492
rect 41916 23214 41918 23266
rect 41970 23214 41972 23266
rect 41916 22484 41972 23214
rect 42140 23044 42196 24108
rect 42140 22978 42196 22988
rect 41916 22418 41972 22428
rect 42252 22258 42308 22270
rect 42252 22206 42254 22258
rect 42306 22206 42308 22258
rect 41916 21812 41972 21822
rect 41916 21718 41972 21756
rect 41804 21532 41972 21588
rect 41916 21362 41972 21532
rect 41916 21310 41918 21362
rect 41970 21310 41972 21362
rect 41804 21028 41860 21038
rect 41804 20934 41860 20972
rect 41580 20078 41582 20130
rect 41634 20078 41636 20130
rect 41468 19348 41524 19358
rect 41468 19254 41524 19292
rect 41580 18676 41636 20078
rect 41804 20244 41860 20254
rect 41804 20018 41860 20188
rect 41804 19966 41806 20018
rect 41858 19966 41860 20018
rect 41692 19906 41748 19918
rect 41692 19854 41694 19906
rect 41746 19854 41748 19906
rect 41692 19460 41748 19854
rect 41692 19394 41748 19404
rect 41804 19236 41860 19966
rect 41580 18610 41636 18620
rect 41692 19180 41860 19236
rect 41692 18452 41748 19180
rect 41916 19124 41972 21310
rect 42140 21476 42196 21486
rect 41916 19058 41972 19068
rect 42028 20018 42084 20030
rect 42028 19966 42030 20018
rect 42082 19966 42084 20018
rect 42028 19908 42084 19966
rect 42140 20020 42196 21420
rect 42252 21028 42308 22206
rect 42252 20962 42308 20972
rect 42364 20916 42420 24332
rect 42476 23716 42532 26852
rect 42588 25506 42644 28812
rect 42812 28642 42868 28654
rect 42812 28590 42814 28642
rect 42866 28590 42868 28642
rect 42812 28082 42868 28590
rect 42812 28030 42814 28082
rect 42866 28030 42868 28082
rect 42812 28018 42868 28030
rect 42700 27858 42756 27870
rect 42700 27806 42702 27858
rect 42754 27806 42756 27858
rect 42700 26402 42756 27806
rect 42924 27860 42980 27870
rect 42924 27766 42980 27804
rect 43036 27636 43092 27646
rect 42700 26350 42702 26402
rect 42754 26350 42756 26402
rect 42700 26338 42756 26350
rect 42812 26740 42868 26750
rect 42812 26290 42868 26684
rect 42812 26238 42814 26290
rect 42866 26238 42868 26290
rect 42812 26226 42868 26238
rect 43036 26292 43092 27580
rect 43148 26852 43204 30828
rect 43260 29204 43316 31500
rect 43596 30100 43652 32510
rect 43708 32562 43876 32564
rect 43708 32510 43822 32562
rect 43874 32510 43876 32562
rect 43708 32508 43876 32510
rect 43708 32004 43764 32508
rect 43820 32498 43876 32508
rect 43708 31938 43764 31948
rect 43820 32340 43876 32350
rect 43820 31668 43876 32284
rect 43932 31668 43988 32732
rect 44044 32562 44100 32574
rect 44044 32510 44046 32562
rect 44098 32510 44100 32562
rect 44044 31892 44100 32510
rect 44156 32450 44212 33068
rect 44268 32564 44324 32574
rect 44268 32470 44324 32508
rect 44156 32398 44158 32450
rect 44210 32398 44212 32450
rect 44156 32386 44212 32398
rect 44044 31826 44100 31836
rect 44156 31780 44212 31790
rect 44156 31686 44212 31724
rect 43932 31612 44100 31668
rect 43820 31602 43876 31612
rect 43932 31444 43988 31454
rect 43820 31218 43876 31230
rect 43820 31166 43822 31218
rect 43874 31166 43876 31218
rect 43820 30996 43876 31166
rect 43820 30930 43876 30940
rect 43932 30994 43988 31388
rect 43932 30942 43934 30994
rect 43986 30942 43988 30994
rect 43596 30034 43652 30044
rect 43820 30770 43876 30782
rect 43820 30718 43822 30770
rect 43874 30718 43876 30770
rect 43820 30100 43876 30718
rect 43932 30660 43988 30942
rect 44044 30996 44100 31612
rect 44268 31556 44324 31566
rect 44268 31220 44324 31500
rect 44268 31154 44324 31164
rect 44380 31108 44436 34412
rect 44604 33124 44660 33134
rect 44716 33124 44772 34636
rect 44828 34626 44884 34636
rect 45164 34580 45220 35420
rect 45052 34468 45108 34478
rect 45052 34356 45108 34412
rect 44940 34300 45108 34356
rect 44940 34130 44996 34300
rect 44940 34078 44942 34130
rect 44994 34078 44996 34130
rect 44940 33684 44996 34078
rect 45164 34130 45220 34524
rect 45164 34078 45166 34130
rect 45218 34078 45220 34130
rect 45052 34020 45108 34030
rect 45052 33926 45108 33964
rect 45164 33684 45220 34078
rect 44940 33628 45108 33684
rect 44604 33122 44772 33124
rect 44604 33070 44606 33122
rect 44658 33070 44772 33122
rect 44604 33068 44772 33070
rect 44492 32900 44548 32910
rect 44492 32004 44548 32844
rect 44604 32340 44660 33068
rect 44604 32274 44660 32284
rect 44716 32562 44772 32574
rect 44716 32510 44718 32562
rect 44770 32510 44772 32562
rect 44492 31778 44548 31948
rect 44604 32004 44660 32014
rect 44716 32004 44772 32510
rect 44604 32002 44772 32004
rect 44604 31950 44606 32002
rect 44658 31950 44772 32002
rect 44604 31948 44772 31950
rect 44828 32452 44884 32462
rect 44604 31938 44660 31948
rect 44492 31726 44494 31778
rect 44546 31726 44548 31778
rect 44492 31714 44548 31726
rect 44716 31666 44772 31678
rect 44716 31614 44718 31666
rect 44770 31614 44772 31666
rect 44380 31052 44548 31108
rect 44156 30996 44212 31006
rect 44044 30994 44212 30996
rect 44044 30942 44158 30994
rect 44210 30942 44212 30994
rect 44044 30940 44212 30942
rect 43932 30594 43988 30604
rect 44044 30212 44100 30222
rect 43820 30034 43876 30044
rect 43932 30210 44100 30212
rect 43932 30158 44046 30210
rect 44098 30158 44100 30210
rect 43932 30156 44100 30158
rect 43484 29986 43540 29998
rect 43484 29934 43486 29986
rect 43538 29934 43540 29986
rect 43484 29764 43540 29934
rect 43260 29138 43316 29148
rect 43372 29426 43428 29438
rect 43372 29374 43374 29426
rect 43426 29374 43428 29426
rect 43260 27858 43316 27870
rect 43260 27806 43262 27858
rect 43314 27806 43316 27858
rect 43260 27076 43316 27806
rect 43372 27298 43428 29374
rect 43372 27246 43374 27298
rect 43426 27246 43428 27298
rect 43372 27234 43428 27246
rect 43260 27010 43316 27020
rect 43372 27074 43428 27086
rect 43372 27022 43374 27074
rect 43426 27022 43428 27074
rect 43372 26964 43428 27022
rect 43372 26898 43428 26908
rect 43484 26908 43540 29708
rect 43820 29652 43876 29662
rect 43596 29204 43652 29214
rect 43596 28644 43652 29148
rect 43596 28588 43764 28644
rect 43596 28308 43652 28318
rect 43596 27748 43652 28252
rect 43596 27076 43652 27692
rect 43596 27010 43652 27020
rect 43708 27524 43764 28588
rect 43708 27074 43764 27468
rect 43708 27022 43710 27074
rect 43762 27022 43764 27074
rect 43708 27010 43764 27022
rect 43484 26852 43652 26908
rect 43148 26796 43316 26852
rect 43148 26292 43204 26302
rect 43036 26290 43204 26292
rect 43036 26238 43150 26290
rect 43202 26238 43204 26290
rect 43036 26236 43204 26238
rect 43148 26226 43204 26236
rect 43036 26066 43092 26078
rect 43036 26014 43038 26066
rect 43090 26014 43092 26066
rect 43036 25620 43092 26014
rect 42588 25454 42590 25506
rect 42642 25454 42644 25506
rect 42588 24052 42644 25454
rect 42700 25564 43092 25620
rect 43260 25732 43316 26796
rect 42700 24388 42756 25564
rect 42924 25396 42980 25406
rect 42812 25284 42868 25322
rect 42924 25302 42980 25340
rect 42812 25218 42868 25228
rect 43036 25284 43092 25294
rect 43036 25190 43092 25228
rect 43148 25282 43204 25294
rect 43148 25230 43150 25282
rect 43202 25230 43204 25282
rect 43036 25060 43092 25070
rect 42812 24834 42868 24846
rect 42812 24782 42814 24834
rect 42866 24782 42868 24834
rect 42812 24612 42868 24782
rect 42812 24546 42868 24556
rect 42700 24332 42980 24388
rect 42588 23986 42644 23996
rect 42700 24164 42756 24174
rect 42700 24050 42756 24108
rect 42700 23998 42702 24050
rect 42754 23998 42756 24050
rect 42700 23986 42756 23998
rect 42812 23716 42868 23726
rect 42476 23660 42644 23716
rect 42476 23492 42532 23502
rect 42476 23378 42532 23436
rect 42476 23326 42478 23378
rect 42530 23326 42532 23378
rect 42476 23314 42532 23326
rect 42476 23156 42532 23166
rect 42476 22372 42532 23100
rect 42588 22596 42644 23660
rect 42588 22530 42644 22540
rect 42812 22594 42868 23660
rect 42812 22542 42814 22594
rect 42866 22542 42868 22594
rect 42812 22530 42868 22542
rect 42476 22370 42644 22372
rect 42476 22318 42478 22370
rect 42530 22318 42644 22370
rect 42476 22316 42644 22318
rect 42476 22306 42532 22316
rect 42364 20850 42420 20860
rect 42476 21698 42532 21710
rect 42476 21646 42478 21698
rect 42530 21646 42532 21698
rect 42476 21588 42532 21646
rect 42476 21026 42532 21532
rect 42588 21700 42644 22316
rect 42588 21476 42644 21644
rect 42588 21410 42644 21420
rect 42700 21586 42756 21598
rect 42700 21534 42702 21586
rect 42754 21534 42756 21586
rect 42476 20974 42478 21026
rect 42530 20974 42532 21026
rect 42476 20468 42532 20974
rect 42700 20692 42756 21534
rect 42812 20804 42868 20814
rect 42812 20710 42868 20748
rect 42700 20626 42756 20636
rect 42476 20402 42532 20412
rect 42812 20244 42868 20254
rect 42812 20130 42868 20188
rect 42812 20078 42814 20130
rect 42866 20078 42868 20130
rect 42812 20066 42868 20078
rect 42588 20020 42644 20030
rect 42140 19964 42308 20020
rect 42028 19234 42084 19852
rect 42252 19572 42308 19964
rect 42252 19516 42420 19572
rect 42028 19182 42030 19234
rect 42082 19182 42084 19234
rect 42028 18674 42084 19182
rect 42028 18622 42030 18674
rect 42082 18622 42084 18674
rect 42028 18610 42084 18622
rect 42252 18562 42308 18574
rect 42252 18510 42254 18562
rect 42306 18510 42308 18562
rect 41580 18396 41748 18452
rect 41804 18450 41860 18462
rect 41804 18398 41806 18450
rect 41858 18398 41860 18450
rect 41468 17668 41524 17678
rect 41244 17444 41300 17454
rect 41468 17444 41524 17612
rect 41244 17442 41524 17444
rect 41244 17390 41246 17442
rect 41298 17390 41524 17442
rect 41244 17388 41524 17390
rect 41244 17378 41300 17388
rect 41132 15876 41188 16716
rect 41356 16322 41412 17388
rect 41468 16882 41524 16894
rect 41468 16830 41470 16882
rect 41522 16830 41524 16882
rect 41468 16772 41524 16830
rect 41468 16706 41524 16716
rect 41580 16884 41636 18396
rect 41804 18116 41860 18398
rect 42252 18452 42308 18510
rect 42252 18386 42308 18396
rect 41916 18228 41972 18238
rect 41916 18134 41972 18172
rect 42252 18228 42308 18238
rect 41692 18060 41804 18116
rect 41692 16996 41748 18060
rect 41804 18050 41860 18060
rect 41692 16930 41748 16940
rect 41804 17780 41860 17790
rect 41356 16270 41358 16322
rect 41410 16270 41412 16322
rect 41356 16258 41412 16270
rect 41132 15810 41188 15820
rect 41244 16098 41300 16110
rect 41244 16046 41246 16098
rect 41298 16046 41300 16098
rect 41244 15316 41300 16046
rect 41580 15538 41636 16828
rect 41580 15486 41582 15538
rect 41634 15486 41636 15538
rect 41580 15474 41636 15486
rect 41244 15250 41300 15260
rect 40796 15092 40852 15102
rect 41020 15092 41300 15148
rect 40796 14308 40852 15036
rect 41244 14642 41300 15092
rect 41244 14590 41246 14642
rect 41298 14590 41300 14642
rect 41132 14420 41188 14430
rect 40796 14306 40964 14308
rect 40796 14254 40798 14306
rect 40850 14254 40964 14306
rect 40796 14252 40964 14254
rect 40796 14242 40852 14252
rect 40796 13522 40852 13534
rect 40796 13470 40798 13522
rect 40850 13470 40852 13522
rect 40796 13188 40852 13470
rect 40908 13412 40964 14252
rect 40908 13346 40964 13356
rect 40908 13188 40964 13198
rect 40796 13186 40964 13188
rect 40796 13134 40910 13186
rect 40962 13134 40964 13186
rect 40796 13132 40964 13134
rect 40908 13122 40964 13132
rect 41020 12964 41076 12974
rect 40908 12852 40964 12862
rect 40908 12758 40964 12796
rect 41020 12292 41076 12908
rect 41132 12852 41188 14364
rect 41132 12786 41188 12796
rect 41020 12226 41076 12236
rect 40572 10834 40740 10836
rect 40572 10782 40574 10834
rect 40626 10782 40740 10834
rect 40572 10780 40740 10782
rect 40908 11172 40964 11182
rect 40572 10770 40628 10780
rect 40348 9604 40404 9614
rect 40348 9266 40404 9548
rect 40348 9214 40350 9266
rect 40402 9214 40404 9266
rect 40348 9202 40404 9214
rect 40908 9266 40964 11116
rect 40908 9214 40910 9266
rect 40962 9214 40964 9266
rect 40908 9202 40964 9214
rect 41020 11170 41076 11182
rect 41020 11118 41022 11170
rect 41074 11118 41076 11170
rect 41020 9604 41076 11118
rect 41244 10052 41300 14590
rect 41692 14420 41748 14430
rect 41692 14326 41748 14364
rect 41804 14084 41860 17724
rect 42140 17780 42196 17790
rect 42252 17780 42308 18172
rect 42140 17778 42308 17780
rect 42140 17726 42142 17778
rect 42194 17726 42308 17778
rect 42140 17724 42308 17726
rect 41916 17668 41972 17678
rect 41916 17574 41972 17612
rect 42140 17556 42196 17724
rect 42140 17490 42196 17500
rect 41916 17108 41972 17118
rect 41916 17014 41972 17052
rect 42364 17106 42420 19516
rect 42588 19346 42644 19964
rect 42700 19794 42756 19806
rect 42700 19742 42702 19794
rect 42754 19742 42756 19794
rect 42700 19684 42756 19742
rect 42700 19618 42756 19628
rect 42924 19684 42980 24332
rect 43036 22370 43092 25004
rect 43148 24722 43204 25230
rect 43148 24670 43150 24722
rect 43202 24670 43204 24722
rect 43148 23940 43204 24670
rect 43260 24052 43316 25676
rect 43372 26628 43428 26638
rect 43372 25060 43428 26572
rect 43372 24994 43428 25004
rect 43596 24388 43652 26852
rect 43708 26852 43764 26862
rect 43708 26514 43764 26796
rect 43820 26628 43876 29596
rect 43932 27858 43988 30156
rect 44044 30146 44100 30156
rect 44156 29876 44212 30940
rect 44156 29810 44212 29820
rect 44268 30322 44324 30334
rect 44268 30270 44270 30322
rect 44322 30270 44324 30322
rect 43932 27806 43934 27858
rect 43986 27806 43988 27858
rect 43932 26852 43988 27806
rect 44044 29538 44100 29550
rect 44044 29486 44046 29538
rect 44098 29486 44100 29538
rect 44044 27746 44100 29486
rect 44044 27694 44046 27746
rect 44098 27694 44100 27746
rect 44044 27682 44100 27694
rect 44156 28980 44212 28990
rect 43932 26786 43988 26796
rect 43820 26572 43988 26628
rect 43708 26462 43710 26514
rect 43762 26462 43764 26514
rect 43708 26450 43764 26462
rect 43820 26404 43876 26414
rect 43820 25844 43876 26348
rect 43820 25778 43876 25788
rect 43932 25730 43988 26572
rect 44044 26516 44100 26526
rect 44044 26422 44100 26460
rect 43932 25678 43934 25730
rect 43986 25678 43988 25730
rect 43932 25666 43988 25678
rect 44156 25620 44212 28924
rect 44268 27300 44324 30270
rect 44492 29652 44548 31052
rect 44604 30660 44660 30670
rect 44604 30434 44660 30604
rect 44604 30382 44606 30434
rect 44658 30382 44660 30434
rect 44604 30370 44660 30382
rect 44716 30212 44772 31614
rect 44828 31218 44884 32396
rect 45052 32116 45108 33628
rect 45164 33618 45220 33628
rect 45276 32786 45332 36428
rect 45388 35474 45444 37100
rect 45500 37090 45556 37100
rect 45948 37090 46004 37100
rect 46060 36932 46116 37436
rect 46396 37380 46452 37390
rect 46396 37286 46452 37324
rect 46284 37268 46340 37278
rect 45948 36876 46116 36932
rect 46172 37044 46228 37054
rect 45500 36708 45556 36718
rect 45500 36614 45556 36652
rect 45836 36484 45892 36494
rect 45836 36390 45892 36428
rect 45948 36260 46004 36876
rect 45948 36194 46004 36204
rect 46060 36370 46116 36382
rect 46060 36318 46062 36370
rect 46114 36318 46116 36370
rect 45724 35924 45780 35934
rect 46060 35924 46116 36318
rect 45724 35922 46116 35924
rect 45724 35870 45726 35922
rect 45778 35870 46116 35922
rect 45724 35868 46116 35870
rect 45724 35858 45780 35868
rect 45388 35422 45390 35474
rect 45442 35422 45444 35474
rect 45388 33460 45444 35422
rect 46060 35476 46116 35486
rect 46060 34802 46116 35420
rect 46060 34750 46062 34802
rect 46114 34750 46116 34802
rect 46060 34738 46116 34750
rect 45500 34690 45556 34702
rect 45500 34638 45502 34690
rect 45554 34638 45556 34690
rect 45500 33684 45556 34638
rect 45500 33618 45556 33628
rect 45612 34692 45668 34702
rect 45612 33460 45668 34636
rect 45388 33394 45444 33404
rect 45500 33404 45668 33460
rect 45276 32734 45278 32786
rect 45330 32734 45332 32786
rect 45276 32722 45332 32734
rect 45500 33234 45556 33404
rect 45500 33182 45502 33234
rect 45554 33182 45556 33234
rect 45052 32050 45108 32060
rect 45164 32562 45220 32574
rect 45164 32510 45166 32562
rect 45218 32510 45220 32562
rect 45052 31892 45108 31902
rect 44828 31166 44830 31218
rect 44882 31166 44884 31218
rect 44828 31108 44884 31166
rect 44940 31220 44996 31230
rect 44940 31126 44996 31164
rect 45052 31218 45108 31836
rect 45052 31166 45054 31218
rect 45106 31166 45108 31218
rect 45052 31154 45108 31166
rect 44828 31042 44884 31052
rect 45164 30660 45220 32510
rect 45388 32562 45444 32574
rect 45388 32510 45390 32562
rect 45442 32510 45444 32562
rect 45164 30594 45220 30604
rect 45276 32004 45332 32014
rect 44716 30156 45220 30212
rect 44940 29876 44996 29886
rect 44716 29652 44772 29662
rect 44492 29650 44772 29652
rect 44492 29598 44718 29650
rect 44770 29598 44772 29650
rect 44492 29596 44772 29598
rect 44716 29586 44772 29596
rect 44940 29426 44996 29820
rect 44940 29374 44942 29426
rect 44994 29374 44996 29426
rect 44940 29362 44996 29374
rect 44380 28644 44436 28654
rect 44380 28550 44436 28588
rect 44716 28530 44772 28542
rect 44716 28478 44718 28530
rect 44770 28478 44772 28530
rect 44268 27186 44324 27244
rect 44268 27134 44270 27186
rect 44322 27134 44324 27186
rect 44268 27122 44324 27134
rect 44492 27746 44548 27758
rect 44492 27694 44494 27746
rect 44546 27694 44548 27746
rect 44492 27188 44548 27694
rect 44716 27748 44772 28478
rect 44716 27682 44772 27692
rect 44828 27972 44884 27982
rect 44492 27122 44548 27132
rect 44268 26628 44324 26638
rect 44268 26402 44324 26572
rect 44380 26516 44436 26526
rect 44436 26460 44660 26516
rect 44380 26450 44436 26460
rect 44268 26350 44270 26402
rect 44322 26350 44324 26402
rect 44268 26338 44324 26350
rect 44044 25564 44212 25620
rect 44492 25732 44548 25742
rect 44492 25618 44548 25676
rect 44492 25566 44494 25618
rect 44546 25566 44548 25618
rect 44044 25508 44100 25564
rect 44492 25554 44548 25566
rect 43820 25452 44100 25508
rect 43596 24322 43652 24332
rect 43708 25172 43764 25182
rect 43596 24052 43652 24062
rect 43260 24050 43652 24052
rect 43260 23998 43598 24050
rect 43650 23998 43652 24050
rect 43260 23996 43652 23998
rect 43596 23986 43652 23996
rect 43708 23940 43764 25116
rect 43148 23884 43428 23940
rect 43148 23716 43204 23726
rect 43148 23622 43204 23660
rect 43036 22318 43038 22370
rect 43090 22318 43092 22370
rect 43036 21252 43092 22318
rect 43148 23154 43204 23166
rect 43148 23102 43150 23154
rect 43202 23102 43204 23154
rect 43148 22146 43204 23102
rect 43260 23042 43316 23054
rect 43260 22990 43262 23042
rect 43314 22990 43316 23042
rect 43260 22820 43316 22990
rect 43260 22754 43316 22764
rect 43372 22596 43428 23884
rect 43708 23874 43764 23884
rect 43484 23156 43540 23166
rect 43484 23062 43540 23100
rect 43708 23156 43764 23166
rect 43820 23156 43876 25452
rect 44156 25396 44212 25406
rect 44044 25340 44156 25396
rect 44044 25338 44100 25340
rect 43708 23154 43876 23156
rect 43708 23102 43710 23154
rect 43762 23102 43876 23154
rect 43708 23100 43876 23102
rect 43708 23090 43764 23100
rect 43148 22094 43150 22146
rect 43202 22094 43204 22146
rect 43148 22082 43204 22094
rect 43260 22540 43428 22596
rect 43708 22596 43764 22606
rect 43036 21196 43204 21252
rect 43036 20804 43092 20814
rect 43036 20710 43092 20748
rect 43036 20468 43092 20478
rect 43036 20130 43092 20412
rect 43036 20078 43038 20130
rect 43090 20078 43092 20130
rect 43036 20066 43092 20078
rect 42924 19618 42980 19628
rect 42588 19294 42590 19346
rect 42642 19294 42644 19346
rect 42588 19282 42644 19294
rect 42812 19572 42868 19582
rect 42812 19348 42868 19516
rect 42924 19348 42980 19358
rect 42812 19346 42980 19348
rect 42812 19294 42926 19346
rect 42978 19294 42980 19346
rect 42812 19292 42980 19294
rect 42924 19282 42980 19292
rect 42924 19124 42980 19134
rect 42476 18788 42532 18798
rect 42476 18562 42532 18732
rect 42476 18510 42478 18562
rect 42530 18510 42532 18562
rect 42476 18498 42532 18510
rect 42588 18564 42644 18574
rect 42476 17892 42532 17902
rect 42588 17892 42644 18508
rect 42476 17890 42644 17892
rect 42476 17838 42478 17890
rect 42530 17838 42644 17890
rect 42476 17836 42644 17838
rect 42476 17826 42532 17836
rect 42364 17054 42366 17106
rect 42418 17054 42420 17106
rect 42364 16212 42420 17054
rect 42924 17778 42980 19068
rect 43148 19012 43204 21196
rect 43148 18946 43204 18956
rect 43036 18340 43092 18350
rect 43036 18246 43092 18284
rect 43260 18228 43316 22540
rect 43372 22372 43428 22382
rect 43372 19460 43428 22316
rect 43708 22146 43764 22540
rect 43708 22094 43710 22146
rect 43762 22094 43764 22146
rect 43708 20804 43764 22094
rect 43596 20692 43652 20702
rect 43596 20598 43652 20636
rect 43596 20132 43652 20142
rect 43484 19906 43540 19918
rect 43484 19854 43486 19906
rect 43538 19854 43540 19906
rect 43484 19796 43540 19854
rect 43484 19730 43540 19740
rect 43372 19404 43540 19460
rect 43260 18162 43316 18172
rect 43372 18338 43428 18350
rect 43372 18286 43374 18338
rect 43426 18286 43428 18338
rect 42924 17726 42926 17778
rect 42978 17726 42980 17778
rect 42812 16884 42868 16894
rect 42700 16882 42868 16884
rect 42700 16830 42814 16882
rect 42866 16830 42868 16882
rect 42700 16828 42868 16830
rect 42364 16146 42420 16156
rect 42476 16772 42532 16782
rect 42252 16098 42308 16110
rect 42252 16046 42254 16098
rect 42306 16046 42308 16098
rect 42028 15988 42084 15998
rect 42084 15932 42196 15988
rect 42028 15894 42084 15932
rect 42140 15426 42196 15932
rect 42140 15374 42142 15426
rect 42194 15374 42196 15426
rect 42140 15362 42196 15374
rect 42252 15428 42308 16046
rect 42252 15362 42308 15372
rect 42364 15652 42420 15662
rect 42364 15426 42420 15596
rect 42364 15374 42366 15426
rect 42418 15374 42420 15426
rect 42364 15362 42420 15374
rect 41692 14028 41860 14084
rect 42028 15316 42084 15326
rect 42028 14420 42084 15260
rect 41244 9986 41300 9996
rect 41356 13636 41412 13646
rect 40460 9156 40516 9166
rect 40460 7698 40516 9100
rect 40460 7646 40462 7698
rect 40514 7646 40516 7698
rect 40460 7634 40516 7646
rect 40908 8484 40964 8494
rect 40908 7698 40964 8428
rect 41020 8146 41076 9548
rect 41020 8094 41022 8146
rect 41074 8094 41076 8146
rect 41020 8082 41076 8094
rect 41132 9492 41188 9502
rect 40908 7646 40910 7698
rect 40962 7646 40964 7698
rect 40908 7634 40964 7646
rect 40572 6468 40628 6478
rect 40348 6132 40404 6142
rect 40572 6132 40628 6412
rect 40348 6130 40628 6132
rect 40348 6078 40350 6130
rect 40402 6078 40628 6130
rect 40348 6076 40628 6078
rect 40348 6066 40404 6076
rect 40124 5852 40292 5908
rect 37996 5236 38052 5246
rect 37996 5122 38052 5180
rect 37996 5070 37998 5122
rect 38050 5070 38052 5122
rect 37996 5058 38052 5070
rect 40124 4564 40180 5852
rect 40124 4498 40180 4508
rect 40236 5684 40292 5694
rect 39564 4340 39620 4350
rect 39564 4246 39620 4284
rect 40236 4116 40292 5628
rect 40572 4898 40628 6076
rect 40572 4846 40574 4898
rect 40626 4846 40628 4898
rect 40572 4834 40628 4846
rect 40796 5908 40852 5918
rect 40796 5124 40852 5852
rect 40460 4564 40516 4574
rect 40460 4470 40516 4508
rect 40796 4562 40852 5068
rect 40796 4510 40798 4562
rect 40850 4510 40852 4562
rect 40796 4498 40852 4510
rect 40908 5682 40964 5694
rect 40908 5630 40910 5682
rect 40962 5630 40964 5682
rect 40236 4050 40292 4060
rect 38444 3892 38500 3902
rect 38444 3666 38500 3836
rect 38444 3614 38446 3666
rect 38498 3614 38500 3666
rect 38444 3444 38500 3614
rect 39228 3668 39284 3678
rect 39228 3554 39284 3612
rect 40908 3668 40964 5630
rect 41132 5346 41188 9436
rect 41356 9044 41412 13580
rect 41580 12740 41636 12750
rect 41468 12404 41524 12414
rect 41468 12310 41524 12348
rect 41468 12068 41524 12078
rect 41468 10836 41524 12012
rect 41580 11284 41636 12684
rect 41692 11508 41748 14028
rect 41804 13860 41860 13870
rect 41804 13858 41972 13860
rect 41804 13806 41806 13858
rect 41858 13806 41972 13858
rect 41804 13804 41972 13806
rect 41804 13794 41860 13804
rect 41916 13188 41972 13804
rect 42028 13746 42084 14364
rect 42476 14418 42532 16716
rect 42700 16548 42756 16828
rect 42812 16818 42868 16828
rect 42924 16660 42980 17726
rect 43372 17668 43428 18286
rect 43372 17602 43428 17612
rect 43372 17444 43428 17454
rect 43484 17444 43540 19404
rect 43596 19348 43652 20076
rect 43596 19282 43652 19292
rect 43372 17442 43540 17444
rect 43372 17390 43374 17442
rect 43426 17390 43540 17442
rect 43372 17388 43540 17390
rect 43596 18676 43652 18686
rect 43372 17378 43428 17388
rect 43372 17220 43428 17230
rect 43372 17106 43428 17164
rect 43372 17054 43374 17106
rect 43426 17054 43428 17106
rect 43372 17042 43428 17054
rect 43596 16884 43652 18620
rect 42700 16482 42756 16492
rect 42812 16604 42980 16660
rect 43372 16828 43652 16884
rect 42476 14366 42478 14418
rect 42530 14366 42532 14418
rect 42028 13694 42030 13746
rect 42082 13694 42084 13746
rect 42028 13682 42084 13694
rect 42252 13972 42308 13982
rect 42028 13188 42084 13198
rect 41916 13132 42028 13188
rect 41804 13074 41860 13086
rect 41804 13022 41806 13074
rect 41858 13022 41860 13074
rect 41804 12852 41860 13022
rect 42028 12962 42084 13132
rect 42028 12910 42030 12962
rect 42082 12910 42084 12962
rect 42028 12898 42084 12910
rect 41804 12786 41860 12796
rect 42252 12402 42308 13916
rect 42476 12516 42532 14366
rect 42700 15314 42756 15326
rect 42700 15262 42702 15314
rect 42754 15262 42756 15314
rect 42700 14306 42756 15262
rect 42700 14254 42702 14306
rect 42754 14254 42756 14306
rect 42700 14196 42756 14254
rect 42700 14130 42756 14140
rect 42812 13972 42868 16604
rect 43260 15874 43316 15886
rect 43260 15822 43262 15874
rect 43314 15822 43316 15874
rect 43260 15652 43316 15822
rect 42924 15316 42980 15326
rect 42924 14642 42980 15260
rect 43036 15204 43092 15242
rect 43036 15138 43092 15148
rect 42924 14590 42926 14642
rect 42978 14590 42980 14642
rect 42924 14578 42980 14590
rect 43148 14532 43204 14542
rect 43260 14532 43316 15596
rect 43148 14530 43316 14532
rect 43148 14478 43150 14530
rect 43202 14478 43316 14530
rect 43148 14476 43316 14478
rect 43148 14466 43204 14476
rect 42924 14420 42980 14430
rect 42924 14326 42980 14364
rect 43036 13972 43092 13982
rect 42812 13970 43092 13972
rect 42812 13918 43038 13970
rect 43090 13918 43092 13970
rect 42812 13916 43092 13918
rect 42700 13636 42756 13646
rect 42700 13542 42756 13580
rect 43036 13076 43092 13916
rect 43036 13010 43092 13020
rect 42588 12852 42644 12862
rect 43260 12852 43316 12862
rect 42588 12850 43316 12852
rect 42588 12798 42590 12850
rect 42642 12798 43262 12850
rect 43314 12798 43316 12850
rect 42588 12796 43316 12798
rect 42588 12786 42644 12796
rect 43260 12786 43316 12796
rect 42476 12460 42868 12516
rect 42252 12350 42254 12402
rect 42306 12350 42308 12402
rect 42252 12338 42308 12350
rect 42364 12292 42420 12302
rect 41804 11620 41860 11630
rect 41804 11526 41860 11564
rect 41692 11442 41748 11452
rect 42252 11508 42308 11518
rect 42252 11414 42308 11452
rect 41580 11228 41748 11284
rect 41580 10836 41636 10846
rect 41468 10834 41636 10836
rect 41468 10782 41582 10834
rect 41634 10782 41636 10834
rect 41468 10780 41636 10782
rect 41580 10770 41636 10780
rect 41692 10050 41748 11228
rect 41692 9998 41694 10050
rect 41746 9998 41748 10050
rect 41692 9986 41748 9998
rect 41916 10498 41972 10510
rect 41916 10446 41918 10498
rect 41970 10446 41972 10498
rect 41916 10052 41972 10446
rect 41916 9986 41972 9996
rect 42140 9604 42196 9614
rect 42140 9510 42196 9548
rect 41804 9380 41860 9390
rect 41804 9266 41860 9324
rect 41804 9214 41806 9266
rect 41858 9214 41860 9266
rect 41804 9202 41860 9214
rect 41356 8484 41412 8988
rect 41356 8418 41412 8428
rect 42252 8372 42308 8382
rect 42364 8372 42420 12236
rect 42700 12292 42756 12302
rect 42700 12198 42756 12236
rect 42588 11172 42644 11248
rect 42644 11116 42756 11172
rect 42588 11106 42644 11116
rect 42588 10948 42644 10958
rect 42588 10834 42644 10892
rect 42588 10782 42590 10834
rect 42642 10782 42644 10834
rect 42588 10770 42644 10782
rect 42476 9602 42532 9614
rect 42476 9550 42478 9602
rect 42530 9550 42532 9602
rect 42476 9156 42532 9550
rect 42588 9156 42644 9166
rect 42476 9100 42588 9156
rect 42588 9062 42644 9100
rect 42252 8370 42420 8372
rect 42252 8318 42254 8370
rect 42306 8318 42420 8370
rect 42252 8316 42420 8318
rect 42252 8306 42308 8316
rect 41804 8148 41860 8158
rect 41804 8054 41860 8092
rect 42700 8148 42756 11116
rect 42812 8370 42868 12460
rect 43372 12402 43428 16828
rect 43484 16436 43540 16446
rect 43484 15314 43540 16380
rect 43596 16100 43652 16110
rect 43708 16100 43764 20748
rect 43820 20356 43876 23100
rect 43932 25284 43988 25294
rect 44044 25286 44046 25338
rect 44098 25286 44100 25338
rect 44156 25330 44212 25340
rect 44044 25274 44100 25286
rect 43932 21476 43988 25228
rect 44156 24724 44212 24734
rect 44156 24630 44212 24668
rect 44492 24164 44548 24174
rect 44492 24050 44548 24108
rect 44492 23998 44494 24050
rect 44546 23998 44548 24050
rect 44492 23986 44548 23998
rect 44044 23940 44100 23950
rect 44044 23846 44100 23884
rect 44492 23266 44548 23278
rect 44492 23214 44494 23266
rect 44546 23214 44548 23266
rect 44380 23154 44436 23166
rect 44380 23102 44382 23154
rect 44434 23102 44436 23154
rect 44380 23044 44436 23102
rect 44380 22978 44436 22988
rect 44380 22484 44436 22494
rect 43932 20804 43988 21420
rect 44044 22258 44100 22270
rect 44044 22206 44046 22258
rect 44098 22206 44100 22258
rect 44044 21028 44100 22206
rect 44380 22148 44436 22428
rect 44492 22372 44548 23214
rect 44492 22306 44548 22316
rect 44492 22148 44548 22158
rect 44380 22146 44548 22148
rect 44380 22094 44494 22146
rect 44546 22094 44548 22146
rect 44380 22092 44548 22094
rect 44492 22082 44548 22092
rect 44156 21700 44212 21710
rect 44156 21586 44212 21644
rect 44156 21534 44158 21586
rect 44210 21534 44212 21586
rect 44156 21522 44212 21534
rect 44044 20962 44100 20972
rect 43932 20748 44100 20804
rect 43932 20580 43988 20590
rect 43932 20486 43988 20524
rect 43820 20300 43988 20356
rect 43820 19236 43876 19246
rect 43820 17332 43876 19180
rect 43820 17266 43876 17276
rect 43932 16212 43988 20300
rect 44044 19796 44100 20748
rect 44268 20692 44324 20702
rect 44268 20242 44324 20636
rect 44268 20190 44270 20242
rect 44322 20190 44324 20242
rect 44268 20178 44324 20190
rect 44380 20578 44436 20590
rect 44380 20526 44382 20578
rect 44434 20526 44436 20578
rect 44268 20020 44324 20030
rect 44268 19926 44324 19964
rect 44044 19730 44100 19740
rect 44380 19684 44436 20526
rect 44604 20356 44660 26460
rect 44828 26514 44884 27916
rect 45164 27972 45220 30156
rect 45164 27906 45220 27916
rect 44940 27858 44996 27870
rect 44940 27806 44942 27858
rect 44994 27806 44996 27858
rect 44940 27076 44996 27806
rect 44940 27010 44996 27020
rect 44828 26462 44830 26514
rect 44882 26462 44884 26514
rect 44828 26450 44884 26462
rect 45164 26740 45220 26750
rect 44716 26404 44772 26414
rect 44716 23378 44772 26348
rect 45052 26402 45108 26414
rect 45052 26350 45054 26402
rect 45106 26350 45108 26402
rect 45052 26180 45108 26350
rect 45164 26402 45220 26684
rect 45164 26350 45166 26402
rect 45218 26350 45220 26402
rect 45164 26338 45220 26350
rect 45052 26124 45220 26180
rect 45164 25844 45220 26124
rect 44716 23326 44718 23378
rect 44770 23326 44772 23378
rect 44716 23314 44772 23326
rect 44828 25788 45220 25844
rect 44828 23044 44884 25788
rect 44716 22260 44772 22270
rect 44716 21924 44772 22204
rect 44716 21858 44772 21868
rect 44604 20290 44660 20300
rect 44380 19618 44436 19628
rect 44604 19796 44660 19806
rect 44268 19572 44324 19582
rect 44156 19348 44212 19358
rect 44156 19254 44212 19292
rect 44044 19234 44100 19246
rect 44044 19182 44046 19234
rect 44098 19182 44100 19234
rect 44044 18564 44100 19182
rect 44156 18564 44212 18574
rect 44044 18562 44212 18564
rect 44044 18510 44158 18562
rect 44210 18510 44212 18562
rect 44044 18508 44212 18510
rect 44044 17892 44100 18508
rect 44156 18498 44212 18508
rect 44268 18564 44324 19516
rect 44268 18432 44324 18508
rect 44604 18452 44660 19740
rect 44716 19012 44772 19022
rect 44716 18918 44772 18956
rect 44828 18564 44884 22988
rect 44940 25508 44996 25518
rect 44940 21698 44996 25452
rect 45052 25396 45108 25406
rect 45052 24722 45108 25340
rect 45276 24946 45332 31948
rect 45388 31220 45444 32510
rect 45500 31892 45556 33182
rect 45612 33122 45668 33134
rect 45612 33070 45614 33122
rect 45666 33070 45668 33122
rect 45612 32564 45668 33070
rect 45612 32498 45668 32508
rect 45724 33122 45780 33134
rect 45724 33070 45726 33122
rect 45778 33070 45780 33122
rect 45724 32004 45780 33070
rect 45724 31938 45780 31948
rect 45948 32562 46004 32574
rect 45948 32510 45950 32562
rect 46002 32510 46004 32562
rect 45500 31826 45556 31836
rect 45948 31556 46004 32510
rect 46172 31780 46228 36988
rect 46284 35922 46340 37212
rect 46620 37156 46676 37774
rect 46844 37828 46900 37838
rect 46620 37090 46676 37100
rect 46732 37266 46788 37278
rect 46732 37214 46734 37266
rect 46786 37214 46788 37266
rect 46284 35870 46286 35922
rect 46338 35870 46340 35922
rect 46284 35858 46340 35870
rect 46732 36258 46788 37214
rect 46732 36206 46734 36258
rect 46786 36206 46788 36258
rect 46732 35924 46788 36206
rect 46732 35858 46788 35868
rect 46844 35698 46900 37772
rect 47180 37826 47236 37838
rect 47180 37774 47182 37826
rect 47234 37774 47236 37826
rect 47180 37044 47236 37774
rect 47180 36978 47236 36988
rect 47292 36708 47348 38892
rect 47404 37490 47460 40348
rect 47516 39058 47572 40796
rect 47516 39006 47518 39058
rect 47570 39006 47572 39058
rect 47516 38994 47572 39006
rect 47740 41076 47796 41086
rect 47740 40516 47796 41020
rect 47740 39618 47796 40460
rect 47740 39566 47742 39618
rect 47794 39566 47796 39618
rect 47628 38948 47684 38958
rect 47740 38948 47796 39566
rect 47628 38946 47796 38948
rect 47628 38894 47630 38946
rect 47682 38894 47796 38946
rect 47628 38892 47796 38894
rect 47628 38882 47684 38892
rect 47852 38668 47908 42028
rect 48076 41188 48132 42478
rect 48188 41970 48244 43372
rect 48412 42866 48468 43596
rect 48412 42814 48414 42866
rect 48466 42814 48468 42866
rect 48412 42802 48468 42814
rect 48524 43540 48580 43550
rect 48188 41918 48190 41970
rect 48242 41918 48244 41970
rect 48188 41906 48244 41918
rect 48524 42084 48580 43484
rect 49084 43540 49140 44270
rect 49084 43474 49140 43484
rect 49196 43652 49252 43662
rect 48972 42532 49028 42542
rect 48972 42530 49140 42532
rect 48972 42478 48974 42530
rect 49026 42478 49140 42530
rect 48972 42476 49140 42478
rect 48972 42466 49028 42476
rect 48524 41970 48580 42028
rect 48524 41918 48526 41970
rect 48578 41918 48580 41970
rect 48524 41906 48580 41918
rect 48524 41300 48580 41310
rect 48076 41132 48244 41188
rect 48076 40964 48132 40974
rect 48076 40870 48132 40908
rect 47964 40628 48020 40638
rect 47964 39508 48020 40572
rect 48188 40628 48244 41132
rect 48188 40562 48244 40572
rect 48524 40626 48580 41244
rect 48972 41076 49028 41086
rect 48524 40574 48526 40626
rect 48578 40574 48580 40626
rect 48300 40516 48356 40526
rect 48300 40514 48468 40516
rect 48300 40462 48302 40514
rect 48354 40462 48468 40514
rect 48300 40460 48468 40462
rect 48300 40450 48356 40460
rect 48076 39508 48132 39518
rect 47964 39506 48356 39508
rect 47964 39454 48078 39506
rect 48130 39454 48356 39506
rect 47964 39452 48356 39454
rect 48076 39442 48132 39452
rect 48300 39058 48356 39452
rect 48300 39006 48302 39058
rect 48354 39006 48356 39058
rect 48300 38994 48356 39006
rect 48412 39060 48468 40460
rect 48524 40404 48580 40574
rect 48636 41074 49028 41076
rect 48636 41022 48974 41074
rect 49026 41022 49028 41074
rect 48636 41020 49028 41022
rect 48636 40626 48692 41020
rect 48972 41010 49028 41020
rect 48636 40574 48638 40626
rect 48690 40574 48692 40626
rect 48636 40562 48692 40574
rect 48748 40628 48804 40638
rect 48748 40404 48804 40572
rect 48524 40338 48580 40348
rect 48636 40348 48804 40404
rect 48524 39396 48580 39406
rect 48524 39302 48580 39340
rect 48524 39060 48580 39070
rect 48412 39058 48580 39060
rect 48412 39006 48526 39058
rect 48578 39006 48580 39058
rect 48412 39004 48580 39006
rect 48524 38994 48580 39004
rect 48188 38834 48244 38846
rect 48188 38782 48190 38834
rect 48242 38782 48244 38834
rect 48188 38668 48244 38782
rect 48636 38668 48692 40348
rect 49084 40292 49140 42476
rect 49196 41074 49252 43596
rect 49308 43204 49364 46508
rect 49420 45444 49476 49534
rect 49532 49364 49588 49646
rect 49980 49698 50036 49710
rect 49980 49646 49982 49698
rect 50034 49646 50036 49698
rect 49980 49588 50036 49646
rect 49980 49522 50036 49532
rect 50316 49698 50372 49710
rect 50316 49646 50318 49698
rect 50370 49646 50372 49698
rect 50316 49586 50372 49646
rect 50316 49534 50318 49586
rect 50370 49534 50372 49586
rect 50316 49522 50372 49534
rect 49532 49298 49588 49308
rect 49980 49138 50036 49150
rect 49980 49086 49982 49138
rect 50034 49086 50036 49138
rect 49532 49028 49588 49038
rect 49532 48934 49588 48972
rect 49756 48468 49812 48478
rect 49644 48130 49700 48142
rect 49644 48078 49646 48130
rect 49698 48078 49700 48130
rect 49644 47458 49700 48078
rect 49644 47406 49646 47458
rect 49698 47406 49700 47458
rect 49644 47394 49700 47406
rect 49644 46676 49700 46686
rect 49644 46582 49700 46620
rect 49756 45890 49812 48412
rect 49868 48356 49924 48366
rect 49868 47124 49924 48300
rect 49868 46898 49924 47068
rect 49868 46846 49870 46898
rect 49922 46846 49924 46898
rect 49868 46834 49924 46846
rect 49980 48130 50036 49086
rect 50428 49026 50484 50372
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50988 49924 51044 49934
rect 50428 48974 50430 49026
rect 50482 48974 50484 49026
rect 50316 48244 50372 48254
rect 50428 48244 50484 48974
rect 50764 49698 50820 49710
rect 50764 49646 50766 49698
rect 50818 49646 50820 49698
rect 50764 48916 50820 49646
rect 50764 48850 50820 48860
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50316 48242 50484 48244
rect 50316 48190 50318 48242
rect 50370 48190 50484 48242
rect 50316 48188 50484 48190
rect 50316 48178 50372 48188
rect 49980 48078 49982 48130
rect 50034 48078 50036 48130
rect 49756 45838 49758 45890
rect 49810 45838 49812 45890
rect 49532 45780 49588 45790
rect 49532 45686 49588 45724
rect 49532 45444 49588 45454
rect 49420 45388 49532 45444
rect 49532 45106 49588 45388
rect 49532 45054 49534 45106
rect 49586 45054 49588 45106
rect 49532 45042 49588 45054
rect 49644 44546 49700 44558
rect 49644 44494 49646 44546
rect 49698 44494 49700 44546
rect 49644 44100 49700 44494
rect 49532 44098 49700 44100
rect 49532 44046 49646 44098
rect 49698 44046 49700 44098
rect 49532 44044 49700 44046
rect 49420 43428 49476 43438
rect 49420 43334 49476 43372
rect 49308 43148 49476 43204
rect 49308 42978 49364 42990
rect 49308 42926 49310 42978
rect 49362 42926 49364 42978
rect 49308 42866 49364 42926
rect 49308 42814 49310 42866
rect 49362 42814 49364 42866
rect 49308 42802 49364 42814
rect 49420 42084 49476 43148
rect 49532 43092 49588 44044
rect 49644 44034 49700 44044
rect 49756 43650 49812 45838
rect 49756 43598 49758 43650
rect 49810 43598 49812 43650
rect 49644 43538 49700 43550
rect 49644 43486 49646 43538
rect 49698 43486 49700 43538
rect 49644 43428 49700 43486
rect 49644 43362 49700 43372
rect 49756 43316 49812 43598
rect 49868 46676 49924 46686
rect 49868 43428 49924 46620
rect 49980 45220 50036 48078
rect 50428 47348 50484 48188
rect 50428 47282 50484 47292
rect 50204 47124 50260 47134
rect 50204 46004 50260 47068
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50316 46564 50372 46574
rect 50316 46470 50372 46508
rect 50764 46564 50820 46574
rect 50764 46228 50820 46508
rect 50316 46004 50372 46014
rect 50204 46002 50372 46004
rect 50204 45950 50318 46002
rect 50370 45950 50372 46002
rect 50204 45948 50372 45950
rect 49980 45154 50036 45164
rect 50092 45892 50148 45902
rect 50092 45106 50148 45836
rect 50092 45054 50094 45106
rect 50146 45054 50148 45106
rect 49980 44548 50036 44558
rect 50092 44548 50148 45054
rect 49980 44546 50148 44548
rect 49980 44494 49982 44546
rect 50034 44494 50148 44546
rect 49980 44492 50148 44494
rect 50204 44772 50260 44782
rect 49980 44482 50036 44492
rect 50204 44436 50260 44716
rect 50204 44322 50260 44380
rect 50204 44270 50206 44322
rect 50258 44270 50260 44322
rect 50204 44258 50260 44270
rect 50316 43988 50372 45948
rect 50764 46002 50820 46172
rect 50764 45950 50766 46002
rect 50818 45950 50820 46002
rect 50764 45938 50820 45950
rect 50876 46562 50932 46574
rect 50876 46510 50878 46562
rect 50930 46510 50932 46562
rect 50876 46452 50932 46510
rect 50876 45668 50932 46396
rect 50988 46116 51044 49868
rect 51324 49924 51380 50654
rect 52108 50482 52164 50494
rect 52108 50430 52110 50482
rect 52162 50430 52164 50482
rect 51324 49858 51380 49868
rect 51660 50036 51716 50046
rect 51324 49700 51380 49710
rect 51100 49698 51380 49700
rect 51100 49646 51326 49698
rect 51378 49646 51380 49698
rect 51100 49644 51380 49646
rect 51100 49138 51156 49644
rect 51324 49634 51380 49644
rect 51100 49086 51102 49138
rect 51154 49086 51156 49138
rect 51100 48468 51156 49086
rect 51548 48804 51604 48814
rect 51100 48402 51156 48412
rect 51436 48802 51604 48804
rect 51436 48750 51550 48802
rect 51602 48750 51604 48802
rect 51436 48748 51604 48750
rect 51324 48356 51380 48366
rect 51324 48262 51380 48300
rect 50988 46050 51044 46060
rect 51100 47348 51156 47358
rect 50876 45602 50932 45612
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50428 45332 50484 45342
rect 50428 44098 50484 45276
rect 50428 44046 50430 44098
rect 50482 44046 50484 44098
rect 50428 44034 50484 44046
rect 50876 44210 50932 44222
rect 50876 44158 50878 44210
rect 50930 44158 50932 44210
rect 50204 43932 50372 43988
rect 50556 43932 50820 43942
rect 50204 43652 50260 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50204 43586 50260 43596
rect 50316 43764 50372 43774
rect 50316 43650 50372 43708
rect 50316 43598 50318 43650
rect 50370 43598 50372 43650
rect 49868 43372 50260 43428
rect 49756 43250 49812 43260
rect 49532 43036 50036 43092
rect 49420 42018 49476 42028
rect 49868 41860 49924 41870
rect 49308 41858 49924 41860
rect 49308 41806 49870 41858
rect 49922 41806 49924 41858
rect 49308 41804 49924 41806
rect 49308 41410 49364 41804
rect 49868 41794 49924 41804
rect 49308 41358 49310 41410
rect 49362 41358 49364 41410
rect 49308 41346 49364 41358
rect 49196 41022 49198 41074
rect 49250 41022 49252 41074
rect 49196 41010 49252 41022
rect 49756 40962 49812 40974
rect 49756 40910 49758 40962
rect 49810 40910 49812 40962
rect 49756 40628 49812 40910
rect 49756 40562 49812 40572
rect 49868 40964 49924 40974
rect 49980 40964 50036 43036
rect 50092 42868 50148 42878
rect 50092 42774 50148 42812
rect 50204 42644 50260 43372
rect 50316 43204 50372 43598
rect 50876 43652 50932 44158
rect 50876 43586 50932 43596
rect 50988 43764 51044 43774
rect 50316 43138 50372 43148
rect 50428 43540 50484 43550
rect 50428 42868 50484 43484
rect 50316 42812 50484 42868
rect 50316 42754 50372 42812
rect 50316 42702 50318 42754
rect 50370 42702 50372 42754
rect 50316 42690 50372 42702
rect 50876 42756 50932 42766
rect 50988 42756 51044 43708
rect 51100 43540 51156 47292
rect 51436 47348 51492 48748
rect 51548 48738 51604 48748
rect 51660 48466 51716 49980
rect 51996 49700 52052 49710
rect 51884 49644 51996 49700
rect 51884 48916 51940 49644
rect 51996 49568 52052 49644
rect 51996 49364 52052 49374
rect 51996 49138 52052 49308
rect 51996 49086 51998 49138
rect 52050 49086 52052 49138
rect 51996 49074 52052 49086
rect 51884 48860 52052 48916
rect 51660 48414 51662 48466
rect 51714 48414 51716 48466
rect 51660 48402 51716 48414
rect 51548 48244 51604 48254
rect 51548 47460 51604 48188
rect 51772 48244 51828 48254
rect 51772 48242 51940 48244
rect 51772 48190 51774 48242
rect 51826 48190 51940 48242
rect 51772 48188 51940 48190
rect 51772 48178 51828 48188
rect 51548 47328 51604 47404
rect 51660 47796 51716 47806
rect 51660 47570 51716 47740
rect 51660 47518 51662 47570
rect 51714 47518 51716 47570
rect 51436 47282 51492 47292
rect 51324 47234 51380 47246
rect 51324 47182 51326 47234
rect 51378 47182 51380 47234
rect 51212 46564 51268 46574
rect 51212 46470 51268 46508
rect 51212 46116 51268 46126
rect 51212 46002 51268 46060
rect 51212 45950 51214 46002
rect 51266 45950 51268 46002
rect 51212 45938 51268 45950
rect 51100 43474 51156 43484
rect 51212 44660 51268 44670
rect 51100 43314 51156 43326
rect 51100 43262 51102 43314
rect 51154 43262 51156 43314
rect 51100 43092 51156 43262
rect 51100 43026 51156 43036
rect 50876 42754 51044 42756
rect 50876 42702 50878 42754
rect 50930 42702 51044 42754
rect 50876 42700 51044 42702
rect 50876 42690 50932 42700
rect 49924 40908 50036 40964
rect 50092 42588 50260 42644
rect 50428 42644 50484 42654
rect 49532 40516 49588 40526
rect 49532 40422 49588 40460
rect 49868 40514 49924 40908
rect 50092 40852 50148 42588
rect 50428 42196 50484 42588
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 51212 42196 51268 44604
rect 51324 44322 51380 47182
rect 51324 44270 51326 44322
rect 51378 44270 51380 44322
rect 51324 43764 51380 44270
rect 51324 43698 51380 43708
rect 51436 46340 51492 46350
rect 51436 45444 51492 46284
rect 51324 43540 51380 43550
rect 51324 43446 51380 43484
rect 50316 42140 50484 42196
rect 50988 42140 51268 42196
rect 50204 42084 50260 42094
rect 50204 41970 50260 42028
rect 50204 41918 50206 41970
rect 50258 41918 50260 41970
rect 50204 41906 50260 41918
rect 50204 40962 50260 40974
rect 50204 40910 50206 40962
rect 50258 40910 50260 40962
rect 50204 40852 50260 40910
rect 49868 40462 49870 40514
rect 49922 40462 49924 40514
rect 49868 40450 49924 40462
rect 49980 40796 50260 40852
rect 49084 40236 49700 40292
rect 49084 39620 49140 39630
rect 49084 39526 49140 39564
rect 49644 39620 49700 40236
rect 49644 39618 49812 39620
rect 49644 39566 49646 39618
rect 49698 39566 49812 39618
rect 49644 39564 49812 39566
rect 49644 39554 49700 39564
rect 47852 38612 48132 38668
rect 47964 37828 48020 37838
rect 47404 37438 47406 37490
rect 47458 37438 47460 37490
rect 47404 37426 47460 37438
rect 47628 37826 48020 37828
rect 47628 37774 47966 37826
rect 48018 37774 48020 37826
rect 47628 37772 48020 37774
rect 47180 36652 47292 36708
rect 47180 36036 47236 36652
rect 47292 36642 47348 36652
rect 47516 37380 47572 37390
rect 47292 36372 47348 36382
rect 47292 36278 47348 36316
rect 47180 35970 47236 35980
rect 46844 35646 46846 35698
rect 46898 35646 46900 35698
rect 46844 35634 46900 35646
rect 46620 35474 46676 35486
rect 46620 35422 46622 35474
rect 46674 35422 46676 35474
rect 46396 34802 46452 34814
rect 46396 34750 46398 34802
rect 46450 34750 46452 34802
rect 46396 34356 46452 34750
rect 46396 34224 46452 34300
rect 46284 34132 46340 34142
rect 46284 32788 46340 34076
rect 46620 33460 46676 35422
rect 46844 35252 46900 35262
rect 46844 34690 46900 35196
rect 46844 34638 46846 34690
rect 46898 34638 46900 34690
rect 46844 34580 46900 34638
rect 46844 34514 46900 34524
rect 47292 34690 47348 34702
rect 47292 34638 47294 34690
rect 47346 34638 47348 34690
rect 47292 34468 47348 34638
rect 47292 34402 47348 34412
rect 47292 34242 47348 34254
rect 47292 34190 47294 34242
rect 47346 34190 47348 34242
rect 46732 34132 46788 34142
rect 46844 34132 46900 34142
rect 46732 34130 46844 34132
rect 46732 34078 46734 34130
rect 46786 34078 46844 34130
rect 46732 34076 46844 34078
rect 46732 34066 46788 34076
rect 46620 33394 46676 33404
rect 46396 33124 46452 33134
rect 46732 33124 46788 33134
rect 46396 33122 46788 33124
rect 46396 33070 46398 33122
rect 46450 33070 46734 33122
rect 46786 33070 46788 33122
rect 46396 33068 46788 33070
rect 46396 33058 46452 33068
rect 46508 32900 46564 33068
rect 46732 33058 46788 33068
rect 46508 32834 46564 32844
rect 46396 32788 46452 32798
rect 46284 32786 46452 32788
rect 46284 32734 46398 32786
rect 46450 32734 46452 32786
rect 46284 32732 46452 32734
rect 46396 32722 46452 32732
rect 46284 32562 46340 32574
rect 46284 32510 46286 32562
rect 46338 32510 46340 32562
rect 46284 32116 46340 32510
rect 46508 32564 46564 32574
rect 46508 32562 46676 32564
rect 46508 32510 46510 32562
rect 46562 32510 46676 32562
rect 46508 32508 46676 32510
rect 46508 32498 46564 32508
rect 46284 32050 46340 32060
rect 46508 32004 46564 32014
rect 45948 31490 46004 31500
rect 46060 31778 46228 31780
rect 46060 31726 46174 31778
rect 46226 31726 46228 31778
rect 46060 31724 46228 31726
rect 45388 31154 45444 31164
rect 45836 31220 45892 31230
rect 45500 30996 45556 31006
rect 45836 30996 45892 31164
rect 45500 30994 45892 30996
rect 45500 30942 45502 30994
rect 45554 30942 45892 30994
rect 45500 30940 45892 30942
rect 45500 30930 45556 30940
rect 45724 30324 45780 30334
rect 45724 30210 45780 30268
rect 45724 30158 45726 30210
rect 45778 30158 45780 30210
rect 45724 30146 45780 30158
rect 45500 30100 45556 30110
rect 45388 29988 45444 29998
rect 45388 29894 45444 29932
rect 45388 28868 45444 28878
rect 45388 28754 45444 28812
rect 45388 28702 45390 28754
rect 45442 28702 45444 28754
rect 45388 27524 45444 28702
rect 45388 27458 45444 27468
rect 45500 27300 45556 30044
rect 45388 27244 45556 27300
rect 45612 29986 45668 29998
rect 45612 29934 45614 29986
rect 45666 29934 45668 29986
rect 45388 26180 45444 27244
rect 45500 26850 45556 26862
rect 45500 26798 45502 26850
rect 45554 26798 45556 26850
rect 45500 26740 45556 26798
rect 45500 26674 45556 26684
rect 45612 26404 45668 29934
rect 46060 29204 46116 31724
rect 46172 31714 46228 31724
rect 46284 31892 46340 31902
rect 46284 31332 46340 31836
rect 46508 31778 46564 31948
rect 46620 31892 46676 32508
rect 46732 31892 46788 31902
rect 46620 31890 46788 31892
rect 46620 31838 46734 31890
rect 46786 31838 46788 31890
rect 46620 31836 46788 31838
rect 46508 31726 46510 31778
rect 46562 31726 46564 31778
rect 46508 31714 46564 31726
rect 46732 31556 46788 31836
rect 46732 31490 46788 31500
rect 46340 31276 46452 31332
rect 46284 31266 46340 31276
rect 46284 30884 46340 30894
rect 46284 30790 46340 30828
rect 46396 30660 46452 31276
rect 46284 30604 46452 30660
rect 46172 30212 46228 30222
rect 46172 30118 46228 30156
rect 45836 29148 46116 29204
rect 45724 27972 45780 27982
rect 45724 27858 45780 27916
rect 45724 27806 45726 27858
rect 45778 27806 45780 27858
rect 45724 27794 45780 27806
rect 45836 27636 45892 29148
rect 46060 28530 46116 28542
rect 46060 28478 46062 28530
rect 46114 28478 46116 28530
rect 45948 27748 46004 27758
rect 45948 27654 46004 27692
rect 45612 26338 45668 26348
rect 45724 27580 45892 27636
rect 45612 26180 45668 26190
rect 45388 26178 45668 26180
rect 45388 26126 45614 26178
rect 45666 26126 45668 26178
rect 45388 26124 45668 26126
rect 45612 26068 45668 26124
rect 45612 26002 45668 26012
rect 45612 25620 45668 25630
rect 45612 25526 45668 25564
rect 45724 25506 45780 27580
rect 45948 27524 46004 27534
rect 45724 25454 45726 25506
rect 45778 25454 45780 25506
rect 45276 24894 45278 24946
rect 45330 24894 45332 24946
rect 45276 24882 45332 24894
rect 45500 25394 45556 25406
rect 45500 25342 45502 25394
rect 45554 25342 45556 25394
rect 45052 24670 45054 24722
rect 45106 24670 45108 24722
rect 45052 24658 45108 24670
rect 45164 24834 45220 24846
rect 45164 24782 45166 24834
rect 45218 24782 45220 24834
rect 45164 24612 45220 24782
rect 45052 23156 45108 23166
rect 45052 23062 45108 23100
rect 44940 21646 44942 21698
rect 44994 21646 44996 21698
rect 44940 21634 44996 21646
rect 45164 21252 45220 24556
rect 45500 24052 45556 25342
rect 45500 23986 45556 23996
rect 45612 24722 45668 24734
rect 45612 24670 45614 24722
rect 45666 24670 45668 24722
rect 45612 24050 45668 24670
rect 45612 23998 45614 24050
rect 45666 23998 45668 24050
rect 45612 23986 45668 23998
rect 45724 23938 45780 25454
rect 45836 26962 45892 26974
rect 45836 26910 45838 26962
rect 45890 26910 45892 26962
rect 45836 25508 45892 26910
rect 45836 25442 45892 25452
rect 45836 24836 45892 24846
rect 45948 24836 46004 27468
rect 46060 26404 46116 28478
rect 46060 26338 46116 26348
rect 46172 26740 46228 26750
rect 46060 26180 46116 26190
rect 46172 26180 46228 26684
rect 46060 26178 46228 26180
rect 46060 26126 46062 26178
rect 46114 26126 46228 26178
rect 46060 26124 46228 26126
rect 46060 26114 46116 26124
rect 46172 25956 46228 26124
rect 46060 25394 46116 25406
rect 46060 25342 46062 25394
rect 46114 25342 46116 25394
rect 46060 25284 46116 25342
rect 46060 25218 46116 25228
rect 46172 25060 46228 25900
rect 45836 24834 46004 24836
rect 45836 24782 45838 24834
rect 45890 24782 46004 24834
rect 45836 24780 46004 24782
rect 45836 24770 45892 24780
rect 45724 23886 45726 23938
rect 45778 23886 45780 23938
rect 45500 23716 45556 23726
rect 45500 23622 45556 23660
rect 45276 23266 45332 23278
rect 45276 23214 45278 23266
rect 45330 23214 45332 23266
rect 45276 22260 45332 23214
rect 45388 23156 45444 23166
rect 45388 23154 45556 23156
rect 45388 23102 45390 23154
rect 45442 23102 45556 23154
rect 45388 23100 45556 23102
rect 45388 23090 45444 23100
rect 45276 22036 45332 22204
rect 45276 21970 45332 21980
rect 45500 22372 45556 23100
rect 44940 21196 45220 21252
rect 44940 20132 44996 21196
rect 45388 20916 45444 20926
rect 45388 20822 45444 20860
rect 44940 19236 44996 20076
rect 45276 20804 45332 20814
rect 45276 20130 45332 20748
rect 45276 20078 45278 20130
rect 45330 20078 45332 20130
rect 45276 20066 45332 20078
rect 45164 20018 45220 20030
rect 45164 19966 45166 20018
rect 45218 19966 45220 20018
rect 45164 19684 45220 19966
rect 45164 19618 45220 19628
rect 45388 19348 45444 19358
rect 44940 19170 44996 19180
rect 45164 19236 45220 19246
rect 44828 18508 44996 18564
rect 44716 18452 44772 18462
rect 44604 18450 44884 18452
rect 44604 18398 44718 18450
rect 44770 18398 44884 18450
rect 44604 18396 44884 18398
rect 44716 18386 44772 18396
rect 44156 18228 44212 18266
rect 44156 18162 44212 18172
rect 44604 18116 44660 18126
rect 44044 17826 44100 17836
rect 44156 18004 44212 18014
rect 44156 17108 44212 17948
rect 44380 18004 44436 18014
rect 44268 17666 44324 17678
rect 44268 17614 44270 17666
rect 44322 17614 44324 17666
rect 44268 17444 44324 17614
rect 44268 17378 44324 17388
rect 44268 17108 44324 17118
rect 44156 17106 44324 17108
rect 44156 17054 44270 17106
rect 44322 17054 44324 17106
rect 44156 17052 44324 17054
rect 44156 16996 44212 17052
rect 44268 17042 44324 17052
rect 44156 16930 44212 16940
rect 44380 16884 44436 17948
rect 44604 17108 44660 18060
rect 44716 17668 44772 17678
rect 44716 17574 44772 17612
rect 44604 17052 44772 17108
rect 44716 16996 44772 17052
rect 44716 16930 44772 16940
rect 44268 16828 44436 16884
rect 44604 16882 44660 16894
rect 44604 16830 44606 16882
rect 44658 16830 44660 16882
rect 44156 16212 44212 16222
rect 43932 16210 44212 16212
rect 43932 16158 44158 16210
rect 44210 16158 44212 16210
rect 43932 16156 44212 16158
rect 44156 16146 44212 16156
rect 43708 16044 44100 16100
rect 43596 16006 43652 16044
rect 43484 15262 43486 15314
rect 43538 15262 43540 15314
rect 43484 15092 43540 15262
rect 43708 15316 43764 15326
rect 43708 15222 43764 15260
rect 43932 15204 43988 15242
rect 43932 15138 43988 15148
rect 43484 15026 43540 15036
rect 43484 14868 43540 14878
rect 43484 13972 43540 14812
rect 43932 14868 43988 14878
rect 43708 14420 43764 14430
rect 43708 14326 43764 14364
rect 43484 13840 43540 13916
rect 43820 14196 43876 14206
rect 43372 12350 43374 12402
rect 43426 12350 43428 12402
rect 43372 12338 43428 12350
rect 43484 13412 43540 13422
rect 43036 11508 43092 11518
rect 43036 11414 43092 11452
rect 43484 11506 43540 13356
rect 43596 12740 43652 12750
rect 43596 12738 43764 12740
rect 43596 12686 43598 12738
rect 43650 12686 43764 12738
rect 43596 12684 43764 12686
rect 43596 12674 43652 12684
rect 43484 11454 43486 11506
rect 43538 11454 43540 11506
rect 43148 10836 43204 10846
rect 43484 10836 43540 11454
rect 43148 10834 43540 10836
rect 43148 10782 43150 10834
rect 43202 10782 43540 10834
rect 43148 10780 43540 10782
rect 43596 12516 43652 12526
rect 43148 10770 43204 10780
rect 43596 10724 43652 12460
rect 43708 12404 43764 12684
rect 43708 12338 43764 12348
rect 43708 12066 43764 12078
rect 43708 12014 43710 12066
rect 43762 12014 43764 12066
rect 43708 11956 43764 12014
rect 43708 11890 43764 11900
rect 43372 10668 43652 10724
rect 43036 10500 43092 10510
rect 43036 9938 43092 10444
rect 43036 9886 43038 9938
rect 43090 9886 43092 9938
rect 43036 9874 43092 9886
rect 43372 9938 43428 10668
rect 43596 10500 43652 10510
rect 43372 9886 43374 9938
rect 43426 9886 43428 9938
rect 42812 8318 42814 8370
rect 42866 8318 42868 8370
rect 42812 8306 42868 8318
rect 43260 8372 43316 8382
rect 43260 8278 43316 8316
rect 42700 8082 42756 8092
rect 42140 7362 42196 7374
rect 42140 7310 42142 7362
rect 42194 7310 42196 7362
rect 41356 6468 41412 6478
rect 41356 6374 41412 6412
rect 41916 6466 41972 6478
rect 41916 6414 41918 6466
rect 41970 6414 41972 6466
rect 41468 5908 41524 5918
rect 41468 5814 41524 5852
rect 41132 5294 41134 5346
rect 41186 5294 41188 5346
rect 41132 5282 41188 5294
rect 41356 5796 41412 5806
rect 40908 3602 40964 3612
rect 41356 3666 41412 5740
rect 41916 5348 41972 6414
rect 42028 5906 42084 5918
rect 42028 5854 42030 5906
rect 42082 5854 42084 5906
rect 42028 5796 42084 5854
rect 42028 5730 42084 5740
rect 41916 5282 41972 5292
rect 41916 5010 41972 5022
rect 41916 4958 41918 5010
rect 41970 4958 41972 5010
rect 41916 4788 41972 4958
rect 41916 4722 41972 4732
rect 42140 4340 42196 7310
rect 42588 7364 42644 7374
rect 42588 6578 42644 7308
rect 43372 6916 43428 9886
rect 43484 10498 43652 10500
rect 43484 10446 43598 10498
rect 43650 10446 43652 10498
rect 43484 10444 43652 10446
rect 43484 9940 43540 10444
rect 43596 10434 43652 10444
rect 43484 9874 43540 9884
rect 43596 10052 43652 10062
rect 43596 8370 43652 9996
rect 43596 8318 43598 8370
rect 43650 8318 43652 8370
rect 43596 8306 43652 8318
rect 43820 8372 43876 14140
rect 43932 11508 43988 14812
rect 44044 14644 44100 16044
rect 44268 15148 44324 16828
rect 44604 16660 44660 16830
rect 44604 16594 44660 16604
rect 44492 16212 44548 16222
rect 44380 15540 44436 15550
rect 44380 15446 44436 15484
rect 44268 15092 44436 15148
rect 44380 14868 44436 15092
rect 44380 14802 44436 14812
rect 44044 14588 44212 14644
rect 44044 14418 44100 14430
rect 44044 14366 44046 14418
rect 44098 14366 44100 14418
rect 44044 14308 44100 14366
rect 44044 13748 44100 14252
rect 44044 13682 44100 13692
rect 44156 13074 44212 14588
rect 44492 14532 44548 16156
rect 44828 15092 44884 18396
rect 44940 18116 44996 18508
rect 44940 18050 44996 18060
rect 45164 18004 45220 19180
rect 45388 18450 45444 19292
rect 45500 18676 45556 22316
rect 45612 19460 45668 19470
rect 45612 19366 45668 19404
rect 45612 18676 45668 18686
rect 45500 18674 45668 18676
rect 45500 18622 45614 18674
rect 45666 18622 45668 18674
rect 45500 18620 45668 18622
rect 45612 18610 45668 18620
rect 45388 18398 45390 18450
rect 45442 18398 45444 18450
rect 45388 18386 45444 18398
rect 45612 18452 45668 18462
rect 45164 17938 45220 17948
rect 45500 17892 45556 17902
rect 44828 15026 44884 15036
rect 44940 17444 44996 17454
rect 44380 14476 44548 14532
rect 44268 13972 44324 13982
rect 44268 13878 44324 13916
rect 44156 13022 44158 13074
rect 44210 13022 44212 13074
rect 44156 13010 44212 13022
rect 44268 12404 44324 12414
rect 44044 11508 44100 11518
rect 43932 11506 44100 11508
rect 43932 11454 44046 11506
rect 44098 11454 44100 11506
rect 43932 11452 44100 11454
rect 44044 11442 44100 11452
rect 44044 10498 44100 10510
rect 44044 10446 44046 10498
rect 44098 10446 44100 10498
rect 43820 8306 43876 8316
rect 43932 10386 43988 10398
rect 43932 10334 43934 10386
rect 43986 10334 43988 10386
rect 43932 9602 43988 10334
rect 43932 9550 43934 9602
rect 43986 9550 43988 9602
rect 43932 8036 43988 9550
rect 44044 9604 44100 10446
rect 44044 9538 44100 9548
rect 44156 8372 44212 8382
rect 44156 8278 44212 8316
rect 43932 7970 43988 7980
rect 43372 6850 43428 6860
rect 42588 6526 42590 6578
rect 42642 6526 42644 6578
rect 42588 6514 42644 6526
rect 43708 6804 43764 6814
rect 43708 4788 43764 6748
rect 43932 5234 43988 5246
rect 43932 5182 43934 5234
rect 43986 5182 43988 5234
rect 43708 4722 43764 4732
rect 43820 5012 43876 5022
rect 42140 4208 42196 4284
rect 41356 3614 41358 3666
rect 41410 3614 41412 3666
rect 41356 3602 41412 3614
rect 41692 3668 41748 3678
rect 41692 3574 41748 3612
rect 43820 3666 43876 4956
rect 43820 3614 43822 3666
rect 43874 3614 43876 3666
rect 43820 3602 43876 3614
rect 39228 3502 39230 3554
rect 39282 3502 39284 3554
rect 39228 3490 39284 3502
rect 38444 3378 38500 3388
rect 40124 3442 40180 3454
rect 40124 3390 40126 3442
rect 40178 3390 40180 3442
rect 40124 3388 40180 3390
rect 42476 3444 42532 3482
rect 38108 3330 38164 3342
rect 40124 3332 40404 3388
rect 42476 3378 42532 3388
rect 43932 3444 43988 5182
rect 44268 4340 44324 12348
rect 44380 11508 44436 14476
rect 44492 14308 44548 14318
rect 44492 14214 44548 14252
rect 44380 11442 44436 11452
rect 44492 13860 44548 13870
rect 44492 13412 44548 13804
rect 44716 13634 44772 13646
rect 44716 13582 44718 13634
rect 44770 13582 44772 13634
rect 44492 11172 44548 13356
rect 44604 13524 44660 13534
rect 44604 13074 44660 13468
rect 44716 13412 44772 13582
rect 44716 13346 44772 13356
rect 44604 13022 44606 13074
rect 44658 13022 44660 13074
rect 44604 13010 44660 13022
rect 44828 12740 44884 12750
rect 44828 12402 44884 12684
rect 44828 12350 44830 12402
rect 44882 12350 44884 12402
rect 44828 12338 44884 12350
rect 44604 12180 44660 12190
rect 44604 12086 44660 12124
rect 44716 11172 44772 11182
rect 44380 10498 44436 10510
rect 44380 10446 44382 10498
rect 44434 10446 44436 10498
rect 44380 10386 44436 10446
rect 44380 10334 44382 10386
rect 44434 10334 44436 10386
rect 44380 10322 44436 10334
rect 44380 9940 44436 9950
rect 44492 9940 44548 11116
rect 44380 9938 44548 9940
rect 44380 9886 44382 9938
rect 44434 9886 44548 9938
rect 44380 9884 44548 9886
rect 44604 11170 44772 11172
rect 44604 11118 44718 11170
rect 44770 11118 44772 11170
rect 44604 11116 44772 11118
rect 44380 9874 44436 9884
rect 44604 8372 44660 11116
rect 44716 11106 44772 11116
rect 44716 10388 44772 10398
rect 44940 10388 44996 17388
rect 45500 17444 45556 17836
rect 45500 17350 45556 17388
rect 45052 16996 45108 17006
rect 45052 15538 45108 16940
rect 45388 16996 45444 17006
rect 45388 16902 45444 16940
rect 45500 16772 45556 16782
rect 45500 16322 45556 16716
rect 45500 16270 45502 16322
rect 45554 16270 45556 16322
rect 45500 16258 45556 16270
rect 45052 15486 45054 15538
rect 45106 15486 45108 15538
rect 45052 15474 45108 15486
rect 45388 16212 45444 16222
rect 45388 15426 45444 16156
rect 45388 15374 45390 15426
rect 45442 15374 45444 15426
rect 45388 15362 45444 15374
rect 45276 15092 45332 15102
rect 45276 14196 45332 15036
rect 45612 14644 45668 18396
rect 45724 18450 45780 23886
rect 45836 24164 45892 24174
rect 45836 23604 45892 24108
rect 45836 23378 45892 23548
rect 45836 23326 45838 23378
rect 45890 23326 45892 23378
rect 45836 23314 45892 23326
rect 45836 22260 45892 22270
rect 45836 22166 45892 22204
rect 45948 22148 46004 24780
rect 46060 25004 46228 25060
rect 46060 22820 46116 25004
rect 46172 23940 46228 23950
rect 46172 23846 46228 23884
rect 46060 22754 46116 22764
rect 46172 22258 46228 22270
rect 46172 22206 46174 22258
rect 46226 22206 46228 22258
rect 46060 22148 46116 22158
rect 45948 22146 46116 22148
rect 45948 22094 46062 22146
rect 46114 22094 46116 22146
rect 45948 22092 46116 22094
rect 45948 21924 46004 21934
rect 45836 21700 45892 21710
rect 45948 21700 46004 21868
rect 45836 21698 46004 21700
rect 45836 21646 45838 21698
rect 45890 21646 46004 21698
rect 45836 21644 46004 21646
rect 45836 21028 45892 21644
rect 45836 20962 45892 20972
rect 46060 21028 46116 22092
rect 46172 21588 46228 22206
rect 46172 21522 46228 21532
rect 46060 20962 46116 20972
rect 45836 20580 45892 20590
rect 45836 20578 46116 20580
rect 45836 20526 45838 20578
rect 45890 20526 46116 20578
rect 45836 20524 46116 20526
rect 45836 20514 45892 20524
rect 45836 20244 45892 20254
rect 45836 20150 45892 20188
rect 45948 19348 46004 19358
rect 45948 19254 46004 19292
rect 45836 19124 45892 19134
rect 45836 19030 45892 19068
rect 46060 19012 46116 20524
rect 46284 20244 46340 30604
rect 46396 29988 46452 29998
rect 46396 29538 46452 29932
rect 46396 29486 46398 29538
rect 46450 29486 46452 29538
rect 46396 29474 46452 29486
rect 46620 29986 46676 29998
rect 46620 29934 46622 29986
rect 46674 29934 46676 29986
rect 46620 28980 46676 29934
rect 46396 28924 46676 28980
rect 46396 27412 46452 28924
rect 46844 28868 46900 34076
rect 47292 33348 47348 34190
rect 47348 33292 47460 33348
rect 47292 33282 47348 33292
rect 47180 33236 47236 33246
rect 46956 33234 47236 33236
rect 46956 33182 47182 33234
rect 47234 33182 47236 33234
rect 46956 33180 47236 33182
rect 46956 31892 47012 33180
rect 47180 33170 47236 33180
rect 47068 33012 47124 33022
rect 47068 32340 47124 32956
rect 47180 32900 47236 32910
rect 47180 32786 47236 32844
rect 47180 32734 47182 32786
rect 47234 32734 47236 32786
rect 47180 32722 47236 32734
rect 47292 32564 47348 32574
rect 47292 32470 47348 32508
rect 47180 32340 47236 32350
rect 47068 32338 47236 32340
rect 47068 32286 47182 32338
rect 47234 32286 47236 32338
rect 47068 32284 47236 32286
rect 47180 32274 47236 32284
rect 46956 31826 47012 31836
rect 47404 31892 47460 33292
rect 47516 32340 47572 37324
rect 47628 34356 47684 37772
rect 47964 37762 48020 37772
rect 48076 37492 48132 38612
rect 47964 37436 48132 37492
rect 48188 38612 48692 38668
rect 49532 39172 49588 39182
rect 47740 37042 47796 37054
rect 47740 36990 47742 37042
rect 47794 36990 47796 37042
rect 47740 36372 47796 36990
rect 47964 36594 48020 37436
rect 48188 36932 48244 38612
rect 49532 38500 49588 39116
rect 49756 38668 49812 39564
rect 49532 38434 49588 38444
rect 49644 38612 49812 38668
rect 49868 38836 49924 38846
rect 49980 38836 50036 40796
rect 49868 38834 50036 38836
rect 49868 38782 49870 38834
rect 49922 38782 50036 38834
rect 49868 38780 50036 38782
rect 50092 40404 50148 40414
rect 48748 37940 48804 37950
rect 48748 37846 48804 37884
rect 48300 37828 48356 37838
rect 49420 37828 49476 37838
rect 48356 37772 48580 37828
rect 48300 37734 48356 37772
rect 48188 36866 48244 36876
rect 48300 37378 48356 37390
rect 48300 37326 48302 37378
rect 48354 37326 48356 37378
rect 47964 36542 47966 36594
rect 48018 36542 48020 36594
rect 47964 36530 48020 36542
rect 48076 36482 48132 36494
rect 48076 36430 48078 36482
rect 48130 36430 48132 36482
rect 48076 36372 48132 36430
rect 47740 36316 48132 36372
rect 47740 35588 47796 35598
rect 47740 35586 47908 35588
rect 47740 35534 47742 35586
rect 47794 35534 47908 35586
rect 47740 35532 47908 35534
rect 47740 35522 47796 35532
rect 47628 33796 47684 34300
rect 47740 34690 47796 34702
rect 47740 34638 47742 34690
rect 47794 34638 47796 34690
rect 47740 33908 47796 34638
rect 47740 33842 47796 33852
rect 47628 33730 47684 33740
rect 47852 33012 47908 35532
rect 47964 33796 48020 33806
rect 47964 33346 48020 33740
rect 47964 33294 47966 33346
rect 48018 33294 48020 33346
rect 47964 33282 48020 33294
rect 47852 32946 47908 32956
rect 47964 32562 48020 32574
rect 47964 32510 47966 32562
rect 48018 32510 48020 32562
rect 47964 32340 48020 32510
rect 47516 32284 47908 32340
rect 47404 31826 47460 31836
rect 47740 31780 47796 31790
rect 47740 31686 47796 31724
rect 47068 31556 47124 31566
rect 47068 31106 47124 31500
rect 47068 31054 47070 31106
rect 47122 31054 47124 31106
rect 46956 30884 47012 30894
rect 46956 29426 47012 30828
rect 47068 30324 47124 31054
rect 47516 31556 47572 31566
rect 47516 31108 47572 31500
rect 47516 30994 47572 31052
rect 47516 30942 47518 30994
rect 47570 30942 47572 30994
rect 47404 30770 47460 30782
rect 47404 30718 47406 30770
rect 47458 30718 47460 30770
rect 47292 30436 47348 30446
rect 47292 30342 47348 30380
rect 47068 30258 47124 30268
rect 47404 30210 47460 30718
rect 47404 30158 47406 30210
rect 47458 30158 47460 30210
rect 47404 30146 47460 30158
rect 47516 29876 47572 30942
rect 47516 29810 47572 29820
rect 47628 30996 47684 31006
rect 46956 29374 46958 29426
rect 47010 29374 47012 29426
rect 46956 29362 47012 29374
rect 46508 28812 46900 28868
rect 47180 29316 47236 29326
rect 46508 28642 46564 28812
rect 47068 28756 47124 28766
rect 46508 28590 46510 28642
rect 46562 28590 46564 28642
rect 46508 28578 46564 28590
rect 46620 28754 47124 28756
rect 46620 28702 47070 28754
rect 47122 28702 47124 28754
rect 46620 28700 47124 28702
rect 46396 27186 46452 27356
rect 46396 27134 46398 27186
rect 46450 27134 46452 27186
rect 46396 27122 46452 27134
rect 46620 26740 46676 28700
rect 47068 28690 47124 28700
rect 47180 28084 47236 29260
rect 47516 29316 47572 29326
rect 47404 28868 47460 28878
rect 47404 28774 47460 28812
rect 47516 28642 47572 29260
rect 47516 28590 47518 28642
rect 47570 28590 47572 28642
rect 47516 28578 47572 28590
rect 47068 28028 47236 28084
rect 46732 27972 46788 27982
rect 46732 27412 46788 27916
rect 46844 27858 46900 27870
rect 46844 27806 46846 27858
rect 46898 27806 46900 27858
rect 46844 27636 46900 27806
rect 46956 27748 47012 27758
rect 46956 27654 47012 27692
rect 46844 27570 46900 27580
rect 46732 27356 46900 27412
rect 46620 26674 46676 26684
rect 46732 26964 46788 26974
rect 46620 26516 46676 26526
rect 46620 26422 46676 26460
rect 46620 26180 46676 26190
rect 46732 26180 46788 26908
rect 46844 26290 46900 27356
rect 46844 26238 46846 26290
rect 46898 26238 46900 26290
rect 46844 26226 46900 26238
rect 46956 26962 47012 26974
rect 46956 26910 46958 26962
rect 47010 26910 47012 26962
rect 46956 26852 47012 26910
rect 46676 26124 46788 26180
rect 46620 25730 46676 26124
rect 46620 25678 46622 25730
rect 46674 25678 46676 25730
rect 46620 25666 46676 25678
rect 46956 25620 47012 26796
rect 46844 25564 47012 25620
rect 46620 25508 46676 25518
rect 46620 25414 46676 25452
rect 46620 24948 46676 24958
rect 46396 23604 46452 23614
rect 46396 22708 46452 23548
rect 46620 23378 46676 24892
rect 46732 24836 46788 24846
rect 46732 24722 46788 24780
rect 46732 24670 46734 24722
rect 46786 24670 46788 24722
rect 46732 24658 46788 24670
rect 46844 23714 46900 25564
rect 46956 25394 47012 25406
rect 46956 25342 46958 25394
rect 47010 25342 47012 25394
rect 46956 25172 47012 25342
rect 46956 25106 47012 25116
rect 47068 24834 47124 28028
rect 47292 27860 47348 27870
rect 47292 27186 47348 27804
rect 47292 27134 47294 27186
rect 47346 27134 47348 27186
rect 47292 27122 47348 27134
rect 47628 26908 47684 30940
rect 47852 28082 47908 32284
rect 47964 32274 48020 32284
rect 48076 32002 48132 36316
rect 48188 36372 48244 36382
rect 48188 36278 48244 36316
rect 48300 35922 48356 37326
rect 48300 35870 48302 35922
rect 48354 35870 48356 35922
rect 48300 35858 48356 35870
rect 48412 37268 48468 37278
rect 48188 35698 48244 35710
rect 48188 35646 48190 35698
rect 48242 35646 48244 35698
rect 48188 34916 48244 35646
rect 48412 35252 48468 37212
rect 48524 37044 48580 37772
rect 48524 36978 48580 36988
rect 49308 37826 49476 37828
rect 49308 37774 49422 37826
rect 49474 37774 49476 37826
rect 49308 37772 49476 37774
rect 48524 36708 48580 36718
rect 48524 35700 48580 36652
rect 48524 35698 48692 35700
rect 48524 35646 48526 35698
rect 48578 35646 48692 35698
rect 48524 35644 48692 35646
rect 48524 35634 48580 35644
rect 48412 35186 48468 35196
rect 48524 34916 48580 34926
rect 48188 34914 48580 34916
rect 48188 34862 48526 34914
rect 48578 34862 48580 34914
rect 48188 34860 48580 34862
rect 48188 34020 48244 34030
rect 48188 34018 48356 34020
rect 48188 33966 48190 34018
rect 48242 33966 48356 34018
rect 48188 33964 48356 33966
rect 48188 33954 48244 33964
rect 48076 31950 48078 32002
rect 48130 31950 48132 32002
rect 48076 31938 48132 31950
rect 48188 33684 48244 33694
rect 47964 31892 48020 31902
rect 47964 30884 48020 31836
rect 47964 30818 48020 30828
rect 48188 31890 48244 33628
rect 48188 31838 48190 31890
rect 48242 31838 48244 31890
rect 48188 30772 48244 31838
rect 48300 31444 48356 33964
rect 48412 33458 48468 34860
rect 48524 34850 48580 34860
rect 48636 34804 48692 35644
rect 48748 35698 48804 35710
rect 48748 35646 48750 35698
rect 48802 35646 48804 35698
rect 48748 34916 48804 35646
rect 48748 34850 48804 34860
rect 48636 34710 48692 34748
rect 48636 34356 48692 34366
rect 48524 34020 48580 34030
rect 48524 33926 48580 33964
rect 48412 33406 48414 33458
rect 48466 33406 48468 33458
rect 48412 33394 48468 33406
rect 48524 33346 48580 33358
rect 48524 33294 48526 33346
rect 48578 33294 48580 33346
rect 48524 33012 48580 33294
rect 48524 32946 48580 32956
rect 48412 32452 48468 32462
rect 48412 32450 48580 32452
rect 48412 32398 48414 32450
rect 48466 32398 48580 32450
rect 48412 32396 48580 32398
rect 48412 32386 48468 32396
rect 48412 31892 48468 31902
rect 48412 31778 48468 31836
rect 48412 31726 48414 31778
rect 48466 31726 48468 31778
rect 48412 31714 48468 31726
rect 48524 31556 48580 32396
rect 48524 31490 48580 31500
rect 48300 31378 48356 31388
rect 48636 31332 48692 34300
rect 49308 34244 49364 37772
rect 49420 37762 49476 37772
rect 49532 37156 49588 37166
rect 49308 34178 49364 34188
rect 49420 37154 49588 37156
rect 49420 37102 49534 37154
rect 49586 37102 49588 37154
rect 49420 37100 49588 37102
rect 49420 34020 49476 37100
rect 49532 37090 49588 37100
rect 49644 36708 49700 38612
rect 49868 38276 49924 38780
rect 50092 38722 50148 40348
rect 50092 38670 50094 38722
rect 50146 38670 50148 38722
rect 50092 38658 50148 38670
rect 49868 38210 49924 38220
rect 50204 38388 50260 38398
rect 50204 38162 50260 38332
rect 50204 38110 50206 38162
rect 50258 38110 50260 38162
rect 50204 38098 50260 38110
rect 49644 36642 49700 36652
rect 49756 37826 49812 37838
rect 49756 37774 49758 37826
rect 49810 37774 49812 37826
rect 49644 36482 49700 36494
rect 49644 36430 49646 36482
rect 49698 36430 49700 36482
rect 49532 35588 49588 35598
rect 49532 35494 49588 35532
rect 49644 35026 49700 36430
rect 49756 36372 49812 37774
rect 49756 36306 49812 36316
rect 50204 37378 50260 37390
rect 50204 37326 50206 37378
rect 50258 37326 50260 37378
rect 49644 34974 49646 35026
rect 49698 34974 49700 35026
rect 49644 34962 49700 34974
rect 49756 35700 49812 35710
rect 49756 34354 49812 35644
rect 50204 35700 50260 37326
rect 50316 37154 50372 42140
rect 50428 41972 50484 41982
rect 50428 41878 50484 41916
rect 50652 40964 50708 40974
rect 50652 40962 50932 40964
rect 50652 40910 50654 40962
rect 50706 40910 50932 40962
rect 50652 40908 50932 40910
rect 50652 40898 50708 40908
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50764 40404 50820 40414
rect 50764 40310 50820 40348
rect 50428 40290 50484 40302
rect 50428 40238 50430 40290
rect 50482 40238 50484 40290
rect 50428 37492 50484 40238
rect 50876 39620 50932 40908
rect 50988 40628 51044 42140
rect 51100 41972 51156 41982
rect 51100 41878 51156 41916
rect 51324 41410 51380 41422
rect 51324 41358 51326 41410
rect 51378 41358 51380 41410
rect 51324 41298 51380 41358
rect 51324 41246 51326 41298
rect 51378 41246 51380 41298
rect 51212 40628 51268 40638
rect 50988 40626 51268 40628
rect 50988 40574 51214 40626
rect 51266 40574 51268 40626
rect 50988 40572 51268 40574
rect 50876 39554 50932 39564
rect 51100 40404 51156 40414
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50988 39060 51044 39070
rect 50988 38966 51044 39004
rect 50540 38836 50596 38846
rect 50540 38742 50596 38780
rect 50652 37828 50708 37838
rect 50652 37826 50932 37828
rect 50652 37774 50654 37826
rect 50706 37774 50932 37826
rect 50652 37772 50932 37774
rect 50652 37762 50708 37772
rect 50876 37716 50932 37772
rect 50556 37660 50820 37670
rect 50876 37660 51044 37716
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50428 37436 50596 37492
rect 50316 37102 50318 37154
rect 50370 37102 50372 37154
rect 50316 37090 50372 37102
rect 50428 37266 50484 37278
rect 50428 37214 50430 37266
rect 50482 37214 50484 37266
rect 50428 35924 50484 37214
rect 50540 37268 50596 37436
rect 50540 37202 50596 37212
rect 50764 37268 50820 37278
rect 50764 37266 50932 37268
rect 50764 37214 50766 37266
rect 50818 37214 50932 37266
rect 50764 37212 50932 37214
rect 50764 37202 50820 37212
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50428 35868 50596 35924
rect 50540 35812 50596 35868
rect 50540 35718 50596 35756
rect 50204 35634 50260 35644
rect 50428 35700 50484 35710
rect 50428 35606 50484 35644
rect 50652 35700 50708 35710
rect 50876 35700 50932 37212
rect 50652 35698 50932 35700
rect 50652 35646 50654 35698
rect 50706 35646 50932 35698
rect 50652 35644 50932 35646
rect 49756 34302 49758 34354
rect 49810 34302 49812 34354
rect 49756 34290 49812 34302
rect 49980 35588 50036 35598
rect 49644 34244 49700 34254
rect 49644 34150 49700 34188
rect 48412 31276 48692 31332
rect 49084 33234 49140 33246
rect 49084 33182 49086 33234
rect 49138 33182 49140 33234
rect 48188 30324 48244 30716
rect 48188 30258 48244 30268
rect 48300 31108 48356 31118
rect 48300 30994 48356 31052
rect 48300 30942 48302 30994
rect 48354 30942 48356 30994
rect 47964 29652 48020 29662
rect 47964 29558 48020 29596
rect 48076 29540 48132 29550
rect 48076 29446 48132 29484
rect 47964 29204 48020 29214
rect 47964 29202 48132 29204
rect 47964 29150 47966 29202
rect 48018 29150 48132 29202
rect 47964 29148 48132 29150
rect 47964 29138 48020 29148
rect 47852 28030 47854 28082
rect 47906 28030 47908 28082
rect 47852 28018 47908 28030
rect 48076 28084 48132 29148
rect 48300 28644 48356 30942
rect 48300 28578 48356 28588
rect 47740 27860 47796 27870
rect 47740 27766 47796 27804
rect 47964 27858 48020 27870
rect 47964 27806 47966 27858
rect 48018 27806 48020 27858
rect 47852 27300 47908 27310
rect 47852 27186 47908 27244
rect 47852 27134 47854 27186
rect 47906 27134 47908 27186
rect 47852 27122 47908 27134
rect 47068 24782 47070 24834
rect 47122 24782 47124 24834
rect 47068 24770 47124 24782
rect 47180 26850 47236 26862
rect 47180 26798 47182 26850
rect 47234 26798 47236 26850
rect 46844 23662 46846 23714
rect 46898 23662 46900 23714
rect 46844 23604 46900 23662
rect 46844 23538 46900 23548
rect 46956 24610 47012 24622
rect 46956 24558 46958 24610
rect 47010 24558 47012 24610
rect 46620 23326 46622 23378
rect 46674 23326 46676 23378
rect 46620 23314 46676 23326
rect 46844 23154 46900 23166
rect 46844 23102 46846 23154
rect 46898 23102 46900 23154
rect 46508 22932 46564 22942
rect 46508 22838 46564 22876
rect 46396 22652 46564 22708
rect 46396 22258 46452 22270
rect 46396 22206 46398 22258
rect 46450 22206 46452 22258
rect 46396 21924 46452 22206
rect 46396 21858 46452 21868
rect 46284 20178 46340 20188
rect 46396 21588 46452 21598
rect 46508 21588 46564 22652
rect 46844 22148 46900 23102
rect 46956 22594 47012 24558
rect 47180 24388 47236 26798
rect 47404 26850 47460 26862
rect 47404 26798 47406 26850
rect 47458 26798 47460 26850
rect 47404 26740 47460 26798
rect 47404 26674 47460 26684
rect 47516 26852 47684 26908
rect 47404 25284 47460 25294
rect 47516 25284 47572 26852
rect 47740 26404 47796 26414
rect 47740 26310 47796 26348
rect 47852 26292 47908 26302
rect 47404 25282 47572 25284
rect 47404 25230 47406 25282
rect 47458 25230 47572 25282
rect 47404 25228 47572 25230
rect 47628 25284 47684 25294
rect 47404 25060 47460 25228
rect 47404 24994 47460 25004
rect 47516 24724 47572 24734
rect 47180 24322 47236 24332
rect 47292 24722 47572 24724
rect 47292 24670 47518 24722
rect 47570 24670 47572 24722
rect 47292 24668 47572 24670
rect 47180 24052 47236 24062
rect 47292 24052 47348 24668
rect 47516 24658 47572 24668
rect 47180 24050 47348 24052
rect 47180 23998 47182 24050
rect 47234 23998 47348 24050
rect 47180 23996 47348 23998
rect 47180 23986 47236 23996
rect 47292 23828 47348 23838
rect 47292 23734 47348 23772
rect 47068 23716 47124 23726
rect 47516 23716 47572 23726
rect 47068 23714 47236 23716
rect 47068 23662 47070 23714
rect 47122 23662 47236 23714
rect 47068 23660 47236 23662
rect 47068 23650 47124 23660
rect 46956 22542 46958 22594
rect 47010 22542 47012 22594
rect 46956 22530 47012 22542
rect 47180 23492 47236 23660
rect 47068 22370 47124 22382
rect 47068 22318 47070 22370
rect 47122 22318 47124 22370
rect 47068 22260 47124 22318
rect 47068 22194 47124 22204
rect 46844 22092 47012 22148
rect 46396 21586 46564 21588
rect 46396 21534 46398 21586
rect 46450 21534 46564 21586
rect 46396 21532 46564 21534
rect 46172 20018 46228 20030
rect 46396 20020 46452 21532
rect 46620 21252 46676 21262
rect 46620 21026 46676 21196
rect 46620 20974 46622 21026
rect 46674 20974 46676 21026
rect 46620 20962 46676 20974
rect 46620 20804 46676 20814
rect 46620 20690 46676 20748
rect 46620 20638 46622 20690
rect 46674 20638 46676 20690
rect 46620 20626 46676 20638
rect 46732 20690 46788 20702
rect 46732 20638 46734 20690
rect 46786 20638 46788 20690
rect 46172 19966 46174 20018
rect 46226 19966 46228 20018
rect 46172 19684 46228 19966
rect 46172 19618 46228 19628
rect 46284 19964 46452 20020
rect 46620 20356 46676 20366
rect 46620 20020 46676 20300
rect 46732 20244 46788 20638
rect 46732 20178 46788 20188
rect 46732 20020 46788 20030
rect 46620 20018 46788 20020
rect 46620 19966 46734 20018
rect 46786 19966 46788 20018
rect 46620 19964 46788 19966
rect 46172 19460 46228 19470
rect 46172 19366 46228 19404
rect 46172 19012 46228 19022
rect 46060 18956 46172 19012
rect 46060 18676 46116 18686
rect 46060 18562 46116 18620
rect 46060 18510 46062 18562
rect 46114 18510 46116 18562
rect 46060 18498 46116 18510
rect 45724 18398 45726 18450
rect 45778 18398 45780 18450
rect 45724 17892 45780 18398
rect 46172 18004 46228 18956
rect 46172 17938 46228 17948
rect 46060 17892 46116 17902
rect 45724 17890 46116 17892
rect 45724 17838 46062 17890
rect 46114 17838 46116 17890
rect 45724 17836 46116 17838
rect 45724 17106 45780 17836
rect 46060 17826 46116 17836
rect 46284 17668 46340 19964
rect 46732 19954 46788 19964
rect 46508 19908 46564 19918
rect 46396 19234 46452 19246
rect 46396 19182 46398 19234
rect 46450 19182 46452 19234
rect 46396 18900 46452 19182
rect 46396 18834 46452 18844
rect 46060 17612 46340 17668
rect 45724 17054 45726 17106
rect 45778 17054 45780 17106
rect 45724 15204 45780 17054
rect 45836 17442 45892 17454
rect 45836 17390 45838 17442
rect 45890 17390 45892 17442
rect 45836 16996 45892 17390
rect 45892 16940 46004 16996
rect 45836 16930 45892 16940
rect 45836 16660 45892 16670
rect 45836 16098 45892 16604
rect 45836 16046 45838 16098
rect 45890 16046 45892 16098
rect 45836 15876 45892 16046
rect 45836 15810 45892 15820
rect 45948 15538 46004 16940
rect 46060 16660 46116 17612
rect 46284 17444 46340 17454
rect 46284 17442 46452 17444
rect 46284 17390 46286 17442
rect 46338 17390 46452 17442
rect 46284 17388 46452 17390
rect 46284 17378 46340 17388
rect 46172 16884 46228 16894
rect 46172 16790 46228 16828
rect 46060 16604 46228 16660
rect 46060 16098 46116 16110
rect 46060 16046 46062 16098
rect 46114 16046 46116 16098
rect 46060 15652 46116 16046
rect 46060 15586 46116 15596
rect 45948 15486 45950 15538
rect 46002 15486 46004 15538
rect 45948 15474 46004 15486
rect 45724 15148 46004 15204
rect 45948 14754 46004 15148
rect 45948 14702 45950 14754
rect 46002 14702 46004 14754
rect 45948 14690 46004 14702
rect 45612 14588 45780 14644
rect 45276 14130 45332 14140
rect 45500 14418 45556 14430
rect 45500 14366 45502 14418
rect 45554 14366 45556 14418
rect 45276 13972 45332 13982
rect 44716 10386 44996 10388
rect 44716 10334 44718 10386
rect 44770 10334 44996 10386
rect 44716 10332 44996 10334
rect 45052 10610 45108 10622
rect 45052 10558 45054 10610
rect 45106 10558 45108 10610
rect 44716 10322 44772 10332
rect 45052 10052 45108 10558
rect 45052 9986 45108 9996
rect 44716 9604 44772 9614
rect 44716 8708 44772 9548
rect 45276 9604 45332 13916
rect 45388 13858 45444 13870
rect 45388 13806 45390 13858
rect 45442 13806 45444 13858
rect 45388 12404 45444 13806
rect 45500 13748 45556 14366
rect 45612 14420 45668 14430
rect 45612 14326 45668 14364
rect 45612 13748 45668 13758
rect 45500 13746 45668 13748
rect 45500 13694 45614 13746
rect 45666 13694 45668 13746
rect 45500 13692 45668 13694
rect 45500 13074 45556 13692
rect 45612 13682 45668 13692
rect 45724 13524 45780 14588
rect 46172 14532 46228 16604
rect 46396 15652 46452 17388
rect 46396 15586 46452 15596
rect 46508 16212 46564 19852
rect 46620 19348 46676 19358
rect 46620 19124 46676 19292
rect 46956 19348 47012 22092
rect 47180 22036 47236 23436
rect 47292 23380 47348 23390
rect 47292 23286 47348 23324
rect 47516 22930 47572 23660
rect 47516 22878 47518 22930
rect 47570 22878 47572 22930
rect 47516 22866 47572 22878
rect 47292 22482 47348 22494
rect 47292 22430 47294 22482
rect 47346 22430 47348 22482
rect 47292 22372 47348 22430
rect 47292 22306 47348 22316
rect 47516 22370 47572 22382
rect 47516 22318 47518 22370
rect 47570 22318 47572 22370
rect 47180 21970 47236 21980
rect 47404 21812 47460 21822
rect 47404 21586 47460 21756
rect 47516 21810 47572 22318
rect 47628 22372 47684 25228
rect 47740 24388 47796 24398
rect 47740 23268 47796 24332
rect 47852 23492 47908 26236
rect 47964 24948 48020 27806
rect 48076 26740 48132 28028
rect 48300 28196 48356 28206
rect 48300 27748 48356 28140
rect 48412 28084 48468 31276
rect 49084 31220 49140 33182
rect 49420 32340 49476 33964
rect 49868 34130 49924 34142
rect 49868 34078 49870 34130
rect 49922 34078 49924 34130
rect 49868 33460 49924 34078
rect 49868 33394 49924 33404
rect 49980 33236 50036 35532
rect 50652 35364 50708 35644
rect 50428 35308 50708 35364
rect 50204 34132 50260 34142
rect 50204 34038 50260 34076
rect 50428 33458 50484 35308
rect 50876 35140 50932 35150
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50652 34244 50708 34254
rect 50652 34150 50708 34188
rect 50428 33406 50430 33458
rect 50482 33406 50484 33458
rect 50428 33394 50484 33406
rect 49868 33180 50036 33236
rect 49532 33122 49588 33134
rect 49532 33070 49534 33122
rect 49586 33070 49588 33122
rect 49532 32788 49588 33070
rect 49868 33124 49924 33180
rect 50316 33124 50372 33134
rect 50540 33124 50596 33134
rect 49532 32732 49812 32788
rect 49644 32562 49700 32574
rect 49644 32510 49646 32562
rect 49698 32510 49700 32562
rect 49532 32340 49588 32350
rect 49420 32284 49532 32340
rect 49308 31780 49364 31790
rect 49308 31686 49364 31724
rect 49420 31220 49476 31230
rect 49084 31218 49476 31220
rect 49084 31166 49422 31218
rect 49474 31166 49476 31218
rect 49084 31164 49476 31166
rect 49420 31154 49476 31164
rect 48636 31108 48692 31118
rect 48524 31106 48692 31108
rect 48524 31054 48638 31106
rect 48690 31054 48692 31106
rect 48524 31052 48692 31054
rect 48524 28980 48580 31052
rect 48636 31042 48692 31052
rect 49532 31106 49588 32284
rect 49644 32116 49700 32510
rect 49644 32050 49700 32060
rect 49756 31892 49812 32732
rect 49756 31826 49812 31836
rect 49532 31054 49534 31106
rect 49586 31054 49588 31106
rect 49532 30996 49588 31054
rect 49196 30940 49588 30996
rect 49644 31666 49700 31678
rect 49644 31614 49646 31666
rect 49698 31614 49700 31666
rect 49644 30996 49700 31614
rect 49756 31556 49812 31566
rect 49756 31218 49812 31500
rect 49868 31554 49924 33068
rect 50092 33122 50372 33124
rect 50092 33070 50318 33122
rect 50370 33070 50372 33122
rect 50092 33068 50372 33070
rect 50092 32786 50148 33068
rect 50316 33058 50372 33068
rect 50428 33122 50596 33124
rect 50428 33070 50542 33122
rect 50594 33070 50596 33122
rect 50428 33068 50596 33070
rect 50092 32734 50094 32786
rect 50146 32734 50148 32786
rect 50092 32722 50148 32734
rect 50428 32676 50484 33068
rect 50540 33058 50596 33068
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50428 32610 50484 32620
rect 50764 32788 50820 32798
rect 49980 32562 50036 32574
rect 49980 32510 49982 32562
rect 50034 32510 50036 32562
rect 49980 32340 50036 32510
rect 50204 32564 50260 32574
rect 50204 32470 50260 32508
rect 49980 32004 50036 32284
rect 50764 32340 50820 32732
rect 50764 32274 50820 32284
rect 49980 31938 50036 31948
rect 49868 31502 49870 31554
rect 49922 31502 49924 31554
rect 49868 31490 49924 31502
rect 50204 31668 50260 31678
rect 49756 31166 49758 31218
rect 49810 31166 49812 31218
rect 49756 31154 49812 31166
rect 49980 30996 50036 31006
rect 49644 30994 50036 30996
rect 49644 30942 49982 30994
rect 50034 30942 50036 30994
rect 49644 30940 50036 30942
rect 48860 30098 48916 30110
rect 48860 30046 48862 30098
rect 48914 30046 48916 30098
rect 48748 29428 48804 29438
rect 48748 29334 48804 29372
rect 48636 29314 48692 29326
rect 48636 29262 48638 29314
rect 48690 29262 48692 29314
rect 48636 29204 48692 29262
rect 48636 29138 48692 29148
rect 48524 28914 48580 28924
rect 48860 28868 48916 30046
rect 48860 28802 48916 28812
rect 48972 28754 49028 28766
rect 48972 28702 48974 28754
rect 49026 28702 49028 28754
rect 48636 28642 48692 28654
rect 48636 28590 48638 28642
rect 48690 28590 48692 28642
rect 48636 28532 48692 28590
rect 48636 28466 48692 28476
rect 48972 28196 49028 28702
rect 48972 28130 49028 28140
rect 48412 28018 48468 28028
rect 48300 27692 48468 27748
rect 48300 27298 48356 27310
rect 48300 27246 48302 27298
rect 48354 27246 48356 27298
rect 48300 27186 48356 27246
rect 48300 27134 48302 27186
rect 48354 27134 48356 27186
rect 48300 27122 48356 27134
rect 48076 26674 48132 26684
rect 48076 26292 48132 26302
rect 48076 26198 48132 26236
rect 48300 26068 48356 26078
rect 48076 25508 48132 25518
rect 48076 25414 48132 25452
rect 48188 25284 48244 25294
rect 48188 25190 48244 25228
rect 47964 24882 48020 24892
rect 48076 24836 48132 24846
rect 47964 24722 48020 24734
rect 47964 24670 47966 24722
rect 48018 24670 48020 24722
rect 47964 24164 48020 24670
rect 48076 24500 48132 24780
rect 48076 24434 48132 24444
rect 48300 24500 48356 26012
rect 48412 25284 48468 27692
rect 48860 27524 48916 27534
rect 48524 26180 48580 26190
rect 48524 26178 48692 26180
rect 48524 26126 48526 26178
rect 48578 26126 48692 26178
rect 48524 26124 48692 26126
rect 48524 26114 48580 26124
rect 48412 25190 48468 25228
rect 48524 25172 48580 25182
rect 48300 24434 48356 24444
rect 48412 24498 48468 24510
rect 48412 24446 48414 24498
rect 48466 24446 48468 24498
rect 48412 24164 48468 24446
rect 47964 24098 48020 24108
rect 48076 24108 48468 24164
rect 47852 23426 47908 23436
rect 47740 23212 47908 23268
rect 47740 23042 47796 23054
rect 47740 22990 47742 23042
rect 47794 22990 47796 23042
rect 47740 22820 47796 22990
rect 47740 22754 47796 22764
rect 47628 22306 47684 22316
rect 47516 21758 47518 21810
rect 47570 21758 47572 21810
rect 47516 21746 47572 21758
rect 47740 21700 47796 21710
rect 47740 21606 47796 21644
rect 47404 21534 47406 21586
rect 47458 21534 47460 21586
rect 47404 20916 47460 21534
rect 47516 21588 47572 21598
rect 47516 21494 47572 21532
rect 47740 21028 47796 21038
rect 47852 21028 47908 23212
rect 47964 21700 48020 21710
rect 48076 21700 48132 24108
rect 48524 24050 48580 25116
rect 48636 24836 48692 26124
rect 48636 24770 48692 24780
rect 48636 24610 48692 24622
rect 48636 24558 48638 24610
rect 48690 24558 48692 24610
rect 48636 24498 48692 24558
rect 48636 24446 48638 24498
rect 48690 24446 48692 24498
rect 48636 24434 48692 24446
rect 48524 23998 48526 24050
rect 48578 23998 48580 24050
rect 48524 23986 48580 23998
rect 48748 24052 48804 24062
rect 48188 23940 48244 23950
rect 48188 23846 48244 23884
rect 48748 23938 48804 23996
rect 48748 23886 48750 23938
rect 48802 23886 48804 23938
rect 48412 23828 48468 23838
rect 48412 23716 48468 23772
rect 48636 23716 48692 23726
rect 48412 23714 48580 23716
rect 48412 23662 48414 23714
rect 48466 23662 48580 23714
rect 48412 23660 48580 23662
rect 48412 23650 48468 23660
rect 48188 23268 48244 23278
rect 48188 22708 48244 23212
rect 48188 22642 48244 22652
rect 48412 22260 48468 22270
rect 48412 22166 48468 22204
rect 47964 21698 48132 21700
rect 47964 21646 47966 21698
rect 48018 21646 48132 21698
rect 47964 21644 48132 21646
rect 48188 22036 48244 22046
rect 47964 21364 48020 21644
rect 47964 21298 48020 21308
rect 47740 21026 47908 21028
rect 47740 20974 47742 21026
rect 47794 20974 47908 21026
rect 47740 20972 47908 20974
rect 47964 21026 48020 21038
rect 47964 20974 47966 21026
rect 48018 20974 48020 21026
rect 47404 20860 47572 20916
rect 47404 20692 47460 20702
rect 47404 20598 47460 20636
rect 47516 20244 47572 20860
rect 47628 20578 47684 20590
rect 47628 20526 47630 20578
rect 47682 20526 47684 20578
rect 47628 20468 47684 20526
rect 47628 20402 47684 20412
rect 47516 20188 47684 20244
rect 47404 20132 47460 20142
rect 47460 20076 47572 20132
rect 47404 20066 47460 20076
rect 47180 20018 47236 20030
rect 47180 19966 47182 20018
rect 47234 19966 47236 20018
rect 47180 19908 47236 19966
rect 47180 19842 47236 19852
rect 47404 19906 47460 19918
rect 47404 19854 47406 19906
rect 47458 19854 47460 19906
rect 47404 19460 47460 19854
rect 47516 19794 47572 20076
rect 47516 19742 47518 19794
rect 47570 19742 47572 19794
rect 47516 19572 47572 19742
rect 47516 19506 47572 19516
rect 47404 19394 47460 19404
rect 46956 19282 47012 19292
rect 46620 18674 46676 19068
rect 47628 19124 47684 20188
rect 47628 19030 47684 19068
rect 46956 19012 47012 19022
rect 46956 18918 47012 18956
rect 47516 18900 47572 18910
rect 46620 18622 46622 18674
rect 46674 18622 46676 18674
rect 46620 18610 46676 18622
rect 46956 18676 47012 18686
rect 46956 18562 47012 18620
rect 46956 18510 46958 18562
rect 47010 18510 47012 18562
rect 46956 18498 47012 18510
rect 47180 18452 47236 18462
rect 46732 17890 46788 17902
rect 46732 17838 46734 17890
rect 46786 17838 46788 17890
rect 46732 17778 46788 17838
rect 46732 17726 46734 17778
rect 46786 17726 46788 17778
rect 46732 17714 46788 17726
rect 47180 17780 47236 18396
rect 47180 17648 47236 17724
rect 46844 17556 46900 17566
rect 46844 17106 46900 17500
rect 46844 17054 46846 17106
rect 46898 17054 46900 17106
rect 46844 17042 46900 17054
rect 47068 17220 47124 17230
rect 46732 16996 46788 17006
rect 46284 15538 46340 15550
rect 46284 15486 46286 15538
rect 46338 15486 46340 15538
rect 46284 15428 46340 15486
rect 46508 15428 46564 16156
rect 46620 16324 46676 16334
rect 46620 15988 46676 16268
rect 46620 15894 46676 15932
rect 46732 15540 46788 16940
rect 46956 15986 47012 15998
rect 46956 15934 46958 15986
rect 47010 15934 47012 15986
rect 46844 15540 46900 15550
rect 46732 15538 46900 15540
rect 46732 15486 46846 15538
rect 46898 15486 46900 15538
rect 46732 15484 46900 15486
rect 46844 15474 46900 15484
rect 46284 15372 46564 15428
rect 46508 15204 46564 15372
rect 46956 15428 47012 15934
rect 46396 15148 46564 15204
rect 46844 15316 46900 15326
rect 46956 15296 47012 15372
rect 46172 14466 46228 14476
rect 46284 14754 46340 14766
rect 46284 14702 46286 14754
rect 46338 14702 46340 14754
rect 45836 14306 45892 14318
rect 45836 14254 45838 14306
rect 45890 14254 45892 14306
rect 45836 14196 45892 14254
rect 45836 14130 45892 14140
rect 46284 14306 46340 14702
rect 46284 14254 46286 14306
rect 46338 14254 46340 14306
rect 45500 13022 45502 13074
rect 45554 13022 45556 13074
rect 45500 13010 45556 13022
rect 45612 13468 45780 13524
rect 45388 12338 45444 12348
rect 45388 12180 45444 12190
rect 45388 11060 45444 12124
rect 45500 11172 45556 11182
rect 45612 11172 45668 13468
rect 46060 13076 46116 13086
rect 45724 12404 45780 12414
rect 45724 12310 45780 12348
rect 45500 11170 45668 11172
rect 45500 11118 45502 11170
rect 45554 11118 45668 11170
rect 45500 11116 45668 11118
rect 45500 11106 45556 11116
rect 45388 10994 45444 11004
rect 45276 9538 45332 9548
rect 45388 10612 45444 10622
rect 45276 9156 45332 9166
rect 44828 9044 44884 9054
rect 44828 8950 44884 8988
rect 44716 8642 44772 8652
rect 44828 8372 44884 8382
rect 44604 8316 44828 8372
rect 44828 8278 44884 8316
rect 45164 7924 45220 7934
rect 44492 6580 44548 6590
rect 44492 6486 44548 6524
rect 44604 6468 44660 6478
rect 44604 6132 44660 6412
rect 44604 6130 44996 6132
rect 44604 6078 44606 6130
rect 44658 6078 44996 6130
rect 44604 6076 44996 6078
rect 44604 6066 44660 6076
rect 44716 5460 44772 5470
rect 44716 5234 44772 5404
rect 44716 5182 44718 5234
rect 44770 5182 44772 5234
rect 44716 5170 44772 5182
rect 44268 4274 44324 4284
rect 43932 3378 43988 3388
rect 44940 3442 44996 6076
rect 45164 6130 45220 7868
rect 45164 6078 45166 6130
rect 45218 6078 45220 6130
rect 45164 6066 45220 6078
rect 45276 3892 45332 9100
rect 45388 5460 45444 10556
rect 45388 5394 45444 5404
rect 45500 10052 45556 10062
rect 45500 9826 45556 9996
rect 45500 9774 45502 9826
rect 45554 9774 45556 9826
rect 45500 9042 45556 9774
rect 45500 8990 45502 9042
rect 45554 8990 45556 9042
rect 45500 8258 45556 8990
rect 45612 9940 45668 11116
rect 45612 8820 45668 9884
rect 45948 9826 46004 9838
rect 45948 9774 45950 9826
rect 46002 9774 46004 9826
rect 45948 9716 46004 9774
rect 45612 8754 45668 8764
rect 45836 9660 45948 9716
rect 45500 8206 45502 8258
rect 45554 8206 45556 8258
rect 45500 6690 45556 8206
rect 45500 6638 45502 6690
rect 45554 6638 45556 6690
rect 45500 5124 45556 6638
rect 45724 7474 45780 7486
rect 45724 7422 45726 7474
rect 45778 7422 45780 7474
rect 45612 5906 45668 5918
rect 45612 5854 45614 5906
rect 45666 5854 45668 5906
rect 45612 5348 45668 5854
rect 45612 5282 45668 5292
rect 45612 5124 45668 5134
rect 45500 5122 45668 5124
rect 45500 5070 45614 5122
rect 45666 5070 45668 5122
rect 45500 5068 45668 5070
rect 45612 5012 45668 5068
rect 45612 4946 45668 4956
rect 45724 5124 45780 7422
rect 45276 3554 45332 3836
rect 45276 3502 45278 3554
rect 45330 3502 45332 3554
rect 45276 3490 45332 3502
rect 44940 3390 44942 3442
rect 44994 3390 44996 3442
rect 44940 3378 44996 3390
rect 38108 3278 38110 3330
rect 38162 3278 38164 3330
rect 38108 2772 38164 3278
rect 38108 2706 38164 2716
rect 37884 1474 37940 1484
rect 40348 800 40404 3332
rect 45724 800 45780 5068
rect 45836 3666 45892 9660
rect 45948 9650 46004 9660
rect 46060 9266 46116 13020
rect 46172 12962 46228 12974
rect 46172 12910 46174 12962
rect 46226 12910 46228 12962
rect 46172 12740 46228 12910
rect 46172 12674 46228 12684
rect 46172 12516 46228 12526
rect 46172 12402 46228 12460
rect 46172 12350 46174 12402
rect 46226 12350 46228 12402
rect 46172 12068 46228 12350
rect 46284 12292 46340 14254
rect 46396 13188 46452 15148
rect 46732 14306 46788 14318
rect 46732 14254 46734 14306
rect 46786 14254 46788 14306
rect 46732 14196 46788 14254
rect 46508 13972 46564 13982
rect 46508 13878 46564 13916
rect 46396 13132 46564 13188
rect 46396 12964 46452 12974
rect 46396 12870 46452 12908
rect 46508 12516 46564 13132
rect 46508 12450 46564 12460
rect 46732 12402 46788 14140
rect 46732 12350 46734 12402
rect 46786 12350 46788 12402
rect 46732 12338 46788 12350
rect 46620 12292 46676 12302
rect 46284 12236 46564 12292
rect 46172 12002 46228 12012
rect 46284 11618 46340 11630
rect 46284 11566 46286 11618
rect 46338 11566 46340 11618
rect 46284 11506 46340 11566
rect 46284 11454 46286 11506
rect 46338 11454 46340 11506
rect 46284 11442 46340 11454
rect 46060 9214 46062 9266
rect 46114 9214 46116 9266
rect 46060 9202 46116 9214
rect 46396 8930 46452 8942
rect 46396 8878 46398 8930
rect 46450 8878 46452 8930
rect 46396 8820 46452 8878
rect 46396 8754 46452 8764
rect 45948 8260 46004 8270
rect 45948 8166 46004 8204
rect 46508 7700 46564 12236
rect 46620 11506 46676 12236
rect 46844 11618 46900 15260
rect 46956 15092 47012 15102
rect 46956 13524 47012 15036
rect 47068 14308 47124 17164
rect 47180 16884 47236 16894
rect 47180 16790 47236 16828
rect 47180 16660 47236 16670
rect 47180 14642 47236 16604
rect 47404 15202 47460 15214
rect 47404 15150 47406 15202
rect 47458 15150 47460 15202
rect 47404 14868 47460 15150
rect 47404 14802 47460 14812
rect 47180 14590 47182 14642
rect 47234 14590 47236 14642
rect 47180 14578 47236 14590
rect 47068 13970 47124 14252
rect 47516 13972 47572 18844
rect 47628 18452 47684 18462
rect 47740 18452 47796 20972
rect 47852 19460 47908 19470
rect 47852 19346 47908 19404
rect 47852 19294 47854 19346
rect 47906 19294 47908 19346
rect 47852 19282 47908 19294
rect 47628 18450 47796 18452
rect 47628 18398 47630 18450
rect 47682 18398 47796 18450
rect 47628 18396 47796 18398
rect 47852 19124 47908 19134
rect 47628 18340 47684 18396
rect 47628 18274 47684 18284
rect 47740 17780 47796 17790
rect 47740 17220 47796 17724
rect 47852 17220 47908 19068
rect 47964 17444 48020 20974
rect 48188 20916 48244 21980
rect 48412 21476 48468 21486
rect 47964 17350 48020 17388
rect 48076 20914 48244 20916
rect 48076 20862 48190 20914
rect 48242 20862 48244 20914
rect 48076 20860 48244 20862
rect 47852 17164 48020 17220
rect 47740 16996 47796 17164
rect 47852 16996 47908 17006
rect 47740 16994 47908 16996
rect 47740 16942 47854 16994
rect 47906 16942 47908 16994
rect 47740 16940 47908 16942
rect 47852 16930 47908 16940
rect 47628 16660 47684 16670
rect 47628 16100 47684 16604
rect 47628 15968 47684 16044
rect 47852 16436 47908 16446
rect 47852 15986 47908 16380
rect 47852 15934 47854 15986
rect 47906 15934 47908 15986
rect 47852 15922 47908 15934
rect 47740 15428 47796 15438
rect 47628 14308 47684 14318
rect 47628 14214 47684 14252
rect 47068 13918 47070 13970
rect 47122 13918 47124 13970
rect 47068 13906 47124 13918
rect 47404 13916 47572 13972
rect 46956 13458 47012 13468
rect 47068 13636 47124 13646
rect 47068 12740 47124 13580
rect 47292 13076 47348 13086
rect 47068 12738 47236 12740
rect 47068 12686 47070 12738
rect 47122 12686 47236 12738
rect 47068 12684 47236 12686
rect 47068 12674 47124 12684
rect 46844 11566 46846 11618
rect 46898 11566 46900 11618
rect 46844 11554 46900 11566
rect 46956 12516 47012 12526
rect 46620 11454 46622 11506
rect 46674 11454 46676 11506
rect 46620 11442 46676 11454
rect 46844 9268 46900 9278
rect 46956 9268 47012 12460
rect 47068 11732 47124 11742
rect 47068 11506 47124 11676
rect 47068 11454 47070 11506
rect 47122 11454 47124 11506
rect 47068 11442 47124 11454
rect 47180 9604 47236 12684
rect 47292 12402 47348 13020
rect 47292 12350 47294 12402
rect 47346 12350 47348 12402
rect 47292 12338 47348 12350
rect 47180 9538 47236 9548
rect 46508 7634 46564 7644
rect 46620 9266 47012 9268
rect 46620 9214 46846 9266
rect 46898 9214 47012 9266
rect 46620 9212 47012 9214
rect 47404 9266 47460 13916
rect 47628 13746 47684 13758
rect 47628 13694 47630 13746
rect 47682 13694 47684 13746
rect 47628 12964 47684 13694
rect 47628 12898 47684 12908
rect 47740 12962 47796 15372
rect 47852 14754 47908 14766
rect 47852 14702 47854 14754
rect 47906 14702 47908 14754
rect 47852 13970 47908 14702
rect 47852 13918 47854 13970
rect 47906 13918 47908 13970
rect 47852 13906 47908 13918
rect 47740 12910 47742 12962
rect 47794 12910 47796 12962
rect 47740 12404 47796 12910
rect 47852 13412 47908 13422
rect 47852 12516 47908 13356
rect 47964 13188 48020 17164
rect 48076 16772 48132 20860
rect 48188 20850 48244 20860
rect 48300 21474 48468 21476
rect 48300 21422 48414 21474
rect 48466 21422 48468 21474
rect 48300 21420 48468 21422
rect 48300 20356 48356 21420
rect 48412 21410 48468 21420
rect 48300 20290 48356 20300
rect 48412 20804 48468 20814
rect 48412 20130 48468 20748
rect 48524 20242 48580 23660
rect 48636 23622 48692 23660
rect 48636 23380 48692 23390
rect 48636 23286 48692 23324
rect 48636 22930 48692 22942
rect 48636 22878 48638 22930
rect 48690 22878 48692 22930
rect 48636 22258 48692 22878
rect 48636 22206 48638 22258
rect 48690 22206 48692 22258
rect 48636 21026 48692 22206
rect 48636 20974 48638 21026
rect 48690 20974 48692 21026
rect 48636 20962 48692 20974
rect 48636 20580 48692 20590
rect 48636 20486 48692 20524
rect 48524 20190 48526 20242
rect 48578 20190 48580 20242
rect 48524 20178 48580 20190
rect 48636 20244 48692 20254
rect 48412 20078 48414 20130
rect 48466 20078 48468 20130
rect 48412 20066 48468 20078
rect 48300 20020 48356 20030
rect 48300 19460 48356 19964
rect 48300 19394 48356 19404
rect 48636 19348 48692 20188
rect 48748 19460 48804 23886
rect 48860 22482 48916 27468
rect 49084 26850 49140 26862
rect 49084 26798 49086 26850
rect 49138 26798 49140 26850
rect 49084 26180 49140 26798
rect 49196 26404 49252 30940
rect 49980 30548 50036 30940
rect 49532 30324 49588 30334
rect 49420 30210 49476 30222
rect 49420 30158 49422 30210
rect 49474 30158 49476 30210
rect 49420 28866 49476 30158
rect 49420 28814 49422 28866
rect 49474 28814 49476 28866
rect 49420 28802 49476 28814
rect 49532 28642 49588 30268
rect 49980 29540 50036 30492
rect 50204 30436 50260 31612
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50876 31332 50932 35084
rect 50988 34244 51044 37660
rect 51100 35922 51156 40348
rect 51212 39620 51268 40572
rect 51212 39554 51268 39564
rect 51212 37828 51268 37838
rect 51212 37734 51268 37772
rect 51324 37716 51380 41246
rect 51436 40404 51492 45388
rect 51548 44098 51604 44110
rect 51548 44046 51550 44098
rect 51602 44046 51604 44098
rect 51548 43652 51604 44046
rect 51660 43876 51716 47518
rect 51884 47572 51940 48188
rect 51996 48132 52052 48860
rect 52108 48356 52164 50430
rect 52108 48290 52164 48300
rect 52220 49588 52276 49598
rect 51996 48076 52164 48132
rect 51884 47458 51940 47516
rect 51884 47406 51886 47458
rect 51938 47406 51940 47458
rect 51884 47394 51940 47406
rect 51996 46900 52052 46910
rect 51996 46786 52052 46844
rect 51996 46734 51998 46786
rect 52050 46734 52052 46786
rect 51996 46722 52052 46734
rect 52108 46676 52164 48076
rect 52220 46676 52276 49532
rect 52332 48466 52388 55468
rect 56588 55412 56756 55468
rect 54348 55300 54404 55310
rect 54348 55206 54404 55244
rect 55132 55300 55188 55310
rect 55132 55206 55188 55244
rect 56028 55186 56084 55198
rect 56028 55134 56030 55186
rect 56082 55134 56084 55186
rect 56028 54516 56084 55134
rect 56028 54450 56084 54460
rect 56588 55074 56644 55412
rect 56588 55022 56590 55074
rect 56642 55022 56644 55074
rect 56588 53844 56644 55022
rect 56588 53778 56644 53788
rect 56924 55300 56980 55310
rect 55356 50708 55412 50718
rect 55356 50428 55412 50652
rect 55356 50372 55524 50428
rect 53228 49924 53284 49934
rect 52444 49700 52500 49710
rect 52444 49606 52500 49644
rect 52892 49700 52948 49710
rect 52892 49606 52948 49644
rect 53228 49698 53284 49868
rect 53228 49646 53230 49698
rect 53282 49646 53284 49698
rect 52668 49476 52724 49486
rect 52332 48414 52334 48466
rect 52386 48414 52388 48466
rect 52332 47124 52388 48414
rect 52332 47058 52388 47068
rect 52444 48468 52500 48478
rect 52444 46900 52500 48412
rect 52668 48356 52724 49420
rect 52780 48804 52836 48814
rect 52780 48802 52948 48804
rect 52780 48750 52782 48802
rect 52834 48750 52948 48802
rect 52780 48748 52948 48750
rect 52780 48738 52836 48748
rect 52780 48356 52836 48366
rect 52668 48354 52836 48356
rect 52668 48302 52782 48354
rect 52834 48302 52836 48354
rect 52668 48300 52836 48302
rect 52780 48290 52836 48300
rect 52668 47348 52724 47358
rect 52556 47236 52612 47246
rect 52556 47142 52612 47180
rect 52444 46844 52612 46900
rect 52444 46676 52500 46686
rect 52220 46620 52388 46676
rect 52108 45892 52164 46620
rect 51996 45836 52164 45892
rect 52220 46452 52276 46462
rect 51996 44546 52052 45836
rect 51996 44494 51998 44546
rect 52050 44494 52052 44546
rect 51996 44482 52052 44494
rect 52108 45668 52164 45678
rect 51884 44100 51940 44110
rect 51660 43810 51716 43820
rect 51772 44098 51940 44100
rect 51772 44046 51886 44098
rect 51938 44046 51940 44098
rect 51772 44044 51940 44046
rect 51548 42754 51604 43596
rect 51548 42702 51550 42754
rect 51602 42702 51604 42754
rect 51548 42084 51604 42702
rect 51660 43650 51716 43662
rect 51660 43598 51662 43650
rect 51714 43598 51716 43650
rect 51660 42644 51716 43598
rect 51660 42578 51716 42588
rect 51548 42018 51604 42028
rect 51548 41860 51604 41870
rect 51548 41766 51604 41804
rect 51548 41412 51604 41422
rect 51772 41412 51828 44044
rect 51884 44034 51940 44044
rect 51548 41410 51828 41412
rect 51548 41358 51550 41410
rect 51602 41358 51828 41410
rect 51548 41356 51828 41358
rect 51884 43876 51940 43886
rect 51548 41346 51604 41356
rect 51884 41300 51940 43820
rect 51996 43764 52052 43774
rect 51996 43650 52052 43708
rect 51996 43598 51998 43650
rect 52050 43598 52052 43650
rect 51996 43586 52052 43598
rect 52108 43652 52164 45612
rect 52220 44434 52276 46396
rect 52332 45332 52388 46620
rect 52444 46582 52500 46620
rect 52556 46116 52612 46844
rect 52444 46060 52612 46116
rect 52668 46114 52724 47292
rect 52892 46900 52948 48748
rect 53228 47796 53284 49646
rect 53788 49698 53844 49710
rect 53788 49646 53790 49698
rect 53842 49646 53844 49698
rect 53452 48804 53508 48814
rect 53452 48710 53508 48748
rect 53228 47730 53284 47740
rect 53340 48356 53396 48366
rect 52668 46062 52670 46114
rect 52722 46062 52724 46114
rect 52444 45556 52500 46060
rect 52668 46050 52724 46062
rect 52780 46844 52892 46900
rect 52556 45780 52612 45790
rect 52556 45686 52612 45724
rect 52444 45500 52612 45556
rect 52444 45332 52500 45342
rect 52332 45330 52500 45332
rect 52332 45278 52446 45330
rect 52498 45278 52500 45330
rect 52332 45276 52500 45278
rect 52332 44996 52388 45276
rect 52444 45266 52500 45276
rect 52332 44930 52388 44940
rect 52220 44382 52222 44434
rect 52274 44382 52276 44434
rect 52220 44370 52276 44382
rect 52108 43596 52388 43652
rect 52108 43428 52164 43438
rect 51996 43426 52164 43428
rect 51996 43374 52110 43426
rect 52162 43374 52164 43426
rect 51996 43372 52164 43374
rect 51996 42084 52052 43372
rect 52108 43362 52164 43372
rect 52220 43428 52276 43438
rect 52108 43204 52164 43214
rect 52108 42194 52164 43148
rect 52220 42642 52276 43372
rect 52220 42590 52222 42642
rect 52274 42590 52276 42642
rect 52220 42578 52276 42590
rect 52108 42142 52110 42194
rect 52162 42142 52164 42194
rect 52108 42130 52164 42142
rect 51996 42018 52052 42028
rect 51660 41244 51940 41300
rect 52220 41860 52276 41870
rect 51436 40338 51492 40348
rect 51548 40964 51604 40974
rect 51436 39396 51492 39406
rect 51436 39058 51492 39340
rect 51436 39006 51438 39058
rect 51490 39006 51492 39058
rect 51436 38948 51492 39006
rect 51436 38882 51492 38892
rect 51548 38668 51604 40908
rect 51324 37650 51380 37660
rect 51436 38612 51604 38668
rect 51660 38668 51716 41244
rect 52108 41076 52164 41086
rect 51772 40964 51828 40974
rect 51772 40870 51828 40908
rect 51884 40628 51940 40638
rect 51884 40534 51940 40572
rect 52108 40404 52164 41020
rect 52220 40962 52276 41804
rect 52220 40910 52222 40962
rect 52274 40910 52276 40962
rect 52220 40516 52276 40910
rect 52332 40740 52388 43596
rect 52444 43314 52500 43326
rect 52444 43262 52446 43314
rect 52498 43262 52500 43314
rect 52444 42194 52500 43262
rect 52444 42142 52446 42194
rect 52498 42142 52500 42194
rect 52444 41076 52500 42142
rect 52444 41010 52500 41020
rect 52556 42754 52612 45500
rect 52668 44100 52724 44110
rect 52668 44006 52724 44044
rect 52780 43652 52836 46844
rect 52892 46834 52948 46844
rect 53340 47684 53396 48300
rect 53452 48244 53508 48254
rect 53452 48150 53508 48188
rect 52892 46676 52948 46686
rect 53340 46676 53396 47628
rect 53676 48130 53732 48142
rect 53676 48078 53678 48130
rect 53730 48078 53732 48130
rect 53676 47572 53732 48078
rect 53788 47684 53844 49646
rect 54236 49700 54292 49710
rect 54236 49698 54516 49700
rect 54236 49646 54238 49698
rect 54290 49646 54516 49698
rect 54236 49644 54516 49646
rect 54236 49634 54292 49644
rect 53900 48802 53956 48814
rect 53900 48750 53902 48802
rect 53954 48750 53956 48802
rect 53900 48468 53956 48750
rect 54348 48804 54404 48814
rect 54348 48710 54404 48748
rect 54236 48468 54292 48478
rect 53956 48466 54292 48468
rect 53956 48414 54238 48466
rect 54290 48414 54292 48466
rect 53956 48412 54292 48414
rect 53900 48336 53956 48412
rect 54236 48402 54292 48412
rect 54460 48020 54516 49644
rect 54572 49698 54628 49710
rect 55132 49700 55188 49710
rect 54572 49646 54574 49698
rect 54626 49646 54628 49698
rect 54572 48244 54628 49646
rect 54572 48178 54628 48188
rect 55020 49698 55188 49700
rect 55020 49646 55134 49698
rect 55186 49646 55188 49698
rect 55020 49644 55188 49646
rect 55020 48244 55076 49644
rect 55132 49634 55188 49644
rect 55468 49698 55524 50372
rect 55468 49646 55470 49698
rect 55522 49646 55524 49698
rect 55132 49028 55188 49038
rect 55468 49028 55524 49646
rect 55132 49026 55524 49028
rect 55132 48974 55134 49026
rect 55186 48974 55524 49026
rect 55132 48972 55524 48974
rect 55132 48962 55188 48972
rect 56028 48914 56084 48926
rect 56028 48862 56030 48914
rect 56082 48862 56084 48914
rect 55020 48178 55076 48188
rect 55468 48804 55524 48814
rect 54348 47964 54516 48020
rect 54684 48132 54740 48142
rect 54236 47796 54292 47806
rect 53788 47628 54180 47684
rect 53732 47516 54068 47572
rect 53564 47460 53620 47470
rect 53676 47440 53732 47516
rect 54012 47460 54068 47516
rect 53452 47348 53508 47358
rect 53452 47254 53508 47292
rect 53564 46898 53620 47404
rect 54012 47366 54068 47404
rect 53564 46846 53566 46898
rect 53618 46846 53620 46898
rect 53564 46834 53620 46846
rect 53788 47346 53844 47358
rect 53788 47294 53790 47346
rect 53842 47294 53844 47346
rect 53788 46676 53844 47294
rect 54124 47236 54180 47628
rect 54236 47682 54292 47740
rect 54236 47630 54238 47682
rect 54290 47630 54292 47682
rect 54236 47618 54292 47630
rect 54012 47180 54180 47236
rect 53340 46620 53732 46676
rect 52892 46582 52948 46620
rect 53228 45780 53284 45790
rect 53228 45330 53284 45724
rect 53452 45780 53508 45818
rect 53452 45714 53508 45724
rect 53228 45278 53230 45330
rect 53282 45278 53284 45330
rect 53228 45266 53284 45278
rect 53452 45556 53508 45566
rect 52668 43596 52836 43652
rect 53116 44660 53172 44670
rect 52668 43314 52724 43596
rect 52780 43428 52836 43438
rect 52780 43426 53060 43428
rect 52780 43374 52782 43426
rect 52834 43374 53060 43426
rect 52780 43372 53060 43374
rect 52780 43362 52836 43372
rect 52668 43262 52670 43314
rect 52722 43262 52724 43314
rect 52668 43250 52724 43262
rect 52556 42702 52558 42754
rect 52610 42702 52612 42754
rect 52556 40852 52612 42702
rect 53004 41076 53060 43372
rect 53116 42196 53172 44604
rect 53452 44322 53508 45500
rect 53676 44882 53732 46620
rect 53788 46610 53844 46620
rect 53900 47012 53956 47022
rect 53900 46674 53956 46956
rect 53900 46622 53902 46674
rect 53954 46622 53956 46674
rect 53788 45666 53844 45678
rect 53788 45614 53790 45666
rect 53842 45614 53844 45666
rect 53788 45332 53844 45614
rect 53900 45556 53956 46622
rect 53900 45490 53956 45500
rect 54012 45444 54068 47180
rect 54348 47012 54404 47964
rect 54348 46946 54404 46956
rect 54460 47460 54516 47470
rect 54460 46898 54516 47404
rect 54460 46846 54462 46898
rect 54514 46846 54516 46898
rect 54460 46834 54516 46846
rect 54572 47236 54628 47246
rect 54236 45668 54292 45678
rect 54012 45378 54068 45388
rect 54124 45666 54292 45668
rect 54124 45614 54238 45666
rect 54290 45614 54292 45666
rect 54124 45612 54292 45614
rect 53788 45266 53844 45276
rect 54012 45220 54068 45230
rect 54012 45126 54068 45164
rect 53676 44830 53678 44882
rect 53730 44830 53732 44882
rect 53676 44548 53732 44830
rect 53676 44482 53732 44492
rect 53788 45106 53844 45118
rect 53788 45054 53790 45106
rect 53842 45054 53844 45106
rect 53452 44270 53454 44322
rect 53506 44270 53508 44322
rect 53340 43540 53396 43550
rect 53228 43428 53284 43438
rect 53228 43334 53284 43372
rect 53340 42866 53396 43484
rect 53340 42814 53342 42866
rect 53394 42814 53396 42866
rect 53340 42802 53396 42814
rect 53116 42064 53172 42140
rect 53004 41020 53396 41076
rect 52332 40674 52388 40684
rect 52444 40796 52612 40852
rect 52668 40964 52724 40974
rect 52220 40450 52276 40460
rect 52332 40516 52388 40526
rect 52444 40516 52500 40796
rect 52332 40514 52500 40516
rect 52332 40462 52334 40514
rect 52386 40462 52500 40514
rect 52332 40460 52500 40462
rect 52556 40628 52612 40638
rect 52556 40514 52612 40572
rect 52556 40462 52558 40514
rect 52610 40462 52612 40514
rect 52108 40338 52164 40348
rect 52332 40292 52388 40460
rect 52556 40450 52612 40462
rect 52220 40236 52388 40292
rect 52444 40346 52500 40358
rect 52444 40294 52446 40346
rect 52498 40294 52500 40346
rect 52444 40292 52500 40294
rect 52108 39620 52164 39630
rect 52108 39394 52164 39564
rect 52108 39342 52110 39394
rect 52162 39342 52164 39394
rect 52108 39330 52164 39342
rect 52108 39060 52164 39070
rect 51996 38948 52052 38958
rect 51996 38854 52052 38892
rect 52108 38668 52164 39004
rect 51660 38612 51828 38668
rect 51436 37268 51492 38612
rect 51324 37212 51492 37268
rect 51212 37156 51268 37166
rect 51212 37062 51268 37100
rect 51212 36484 51268 36494
rect 51324 36484 51380 37212
rect 51212 36482 51380 36484
rect 51212 36430 51214 36482
rect 51266 36430 51380 36482
rect 51212 36428 51380 36430
rect 51212 36418 51268 36428
rect 51100 35870 51102 35922
rect 51154 35870 51156 35922
rect 51100 35858 51156 35870
rect 51660 35924 51716 35934
rect 51548 35812 51604 35822
rect 51548 35718 51604 35756
rect 51660 34914 51716 35868
rect 51660 34862 51662 34914
rect 51714 34862 51716 34914
rect 51660 34850 51716 34862
rect 51324 34804 51380 34814
rect 51324 34354 51380 34748
rect 51324 34302 51326 34354
rect 51378 34302 51380 34354
rect 51324 34290 51380 34302
rect 50988 34178 51044 34188
rect 51772 33796 51828 38612
rect 51996 38612 52164 38668
rect 51884 38050 51940 38062
rect 51884 37998 51886 38050
rect 51938 37998 51940 38050
rect 51884 37716 51940 37998
rect 51884 37650 51940 37660
rect 51884 35812 51940 35822
rect 51884 35718 51940 35756
rect 51996 35140 52052 38612
rect 52108 38050 52164 38062
rect 52108 37998 52110 38050
rect 52162 37998 52164 38050
rect 52108 37268 52164 37998
rect 52108 37202 52164 37212
rect 52220 36820 52276 40236
rect 52444 40226 52500 40236
rect 52556 40180 52612 40190
rect 52444 40068 52500 40078
rect 52332 39172 52388 39182
rect 52332 39058 52388 39116
rect 52332 39006 52334 39058
rect 52386 39006 52388 39058
rect 52332 38994 52388 39006
rect 52332 38052 52388 38062
rect 52332 37380 52388 37996
rect 52332 37314 52388 37324
rect 52220 36764 52388 36820
rect 52220 36596 52276 36606
rect 52220 36502 52276 36540
rect 52108 36484 52164 36494
rect 52108 36390 52164 36428
rect 52220 35698 52276 35710
rect 52220 35646 52222 35698
rect 52274 35646 52276 35698
rect 52220 35588 52276 35646
rect 52220 35522 52276 35532
rect 51996 35074 52052 35084
rect 52108 35364 52164 35374
rect 51996 34916 52052 34926
rect 51996 34468 52052 34860
rect 51996 34402 52052 34412
rect 51884 34244 51940 34254
rect 51884 34130 51940 34188
rect 51884 34078 51886 34130
rect 51938 34078 51940 34130
rect 51884 34066 51940 34078
rect 51772 33740 51940 33796
rect 51436 33572 51492 33582
rect 51436 33478 51492 33516
rect 51548 33460 51604 33470
rect 51548 33366 51604 33404
rect 50988 33348 51044 33358
rect 50988 33124 51044 33292
rect 50988 33058 51044 33068
rect 51660 33122 51716 33134
rect 51660 33070 51662 33122
rect 51714 33070 51716 33122
rect 51660 32788 51716 33070
rect 51660 32722 51716 32732
rect 51772 32676 51828 32686
rect 51100 32562 51156 32574
rect 51100 32510 51102 32562
rect 51154 32510 51156 32562
rect 50988 32004 51044 32014
rect 50988 31666 51044 31948
rect 51100 31780 51156 32510
rect 51548 32450 51604 32462
rect 51548 32398 51550 32450
rect 51602 32398 51604 32450
rect 51436 31892 51492 31902
rect 51324 31780 51380 31790
rect 51436 31780 51492 31836
rect 51100 31778 51492 31780
rect 51100 31726 51326 31778
rect 51378 31726 51492 31778
rect 51100 31724 51492 31726
rect 51324 31714 51380 31724
rect 50988 31614 50990 31666
rect 51042 31614 51044 31666
rect 50988 31602 51044 31614
rect 50876 31276 51044 31332
rect 50204 30370 50260 30380
rect 50428 31220 50484 31230
rect 50428 30324 50484 31164
rect 50428 30258 50484 30268
rect 50540 31108 50596 31118
rect 50204 29986 50260 29998
rect 50540 29988 50596 31052
rect 50876 31106 50932 31118
rect 50876 31054 50878 31106
rect 50930 31054 50932 31106
rect 50876 30996 50932 31054
rect 50876 30930 50932 30940
rect 50988 31106 51044 31276
rect 51548 31220 51604 32398
rect 51548 31154 51604 31164
rect 50988 31054 50990 31106
rect 51042 31054 51044 31106
rect 50876 30772 50932 30782
rect 50876 30678 50932 30716
rect 50988 30436 51044 31054
rect 51660 30994 51716 31006
rect 51660 30942 51662 30994
rect 51714 30942 51716 30994
rect 51660 30772 51716 30942
rect 51660 30706 51716 30716
rect 50988 30380 51156 30436
rect 50204 29934 50206 29986
rect 50258 29934 50260 29986
rect 50204 29764 50260 29934
rect 50204 29698 50260 29708
rect 50428 29932 50596 29988
rect 50988 30098 51044 30110
rect 50988 30046 50990 30098
rect 51042 30046 51044 30098
rect 49980 29474 50036 29484
rect 49756 29428 49812 29438
rect 49532 28590 49534 28642
rect 49586 28590 49588 28642
rect 49420 26964 49476 27002
rect 49420 26898 49476 26908
rect 49196 26338 49252 26348
rect 49532 26180 49588 28590
rect 49644 29372 49756 29428
rect 49644 27860 49700 29372
rect 49756 29334 49812 29372
rect 50204 29428 50260 29438
rect 49980 29314 50036 29326
rect 49980 29262 49982 29314
rect 50034 29262 50036 29314
rect 49980 28644 50036 29262
rect 50092 29202 50148 29214
rect 50092 29150 50094 29202
rect 50146 29150 50148 29202
rect 50092 28756 50148 29150
rect 50092 28690 50148 28700
rect 49980 28578 50036 28588
rect 49868 28530 49924 28542
rect 49868 28478 49870 28530
rect 49922 28478 49924 28530
rect 49868 28308 49924 28478
rect 50204 28420 50260 29372
rect 49868 28242 49924 28252
rect 49980 28364 50260 28420
rect 49868 28084 49924 28094
rect 49868 27990 49924 28028
rect 49644 27728 49700 27804
rect 49980 27748 50036 28364
rect 50428 28308 50484 29932
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50876 29540 50932 29550
rect 50876 29446 50932 29484
rect 50988 29204 51044 30046
rect 51100 30100 51156 30380
rect 51324 30434 51380 30446
rect 51324 30382 51326 30434
rect 51378 30382 51380 30434
rect 51100 30034 51156 30044
rect 51212 30322 51268 30334
rect 51212 30270 51214 30322
rect 51266 30270 51268 30322
rect 51212 29204 51268 30270
rect 50988 29202 51156 29204
rect 50988 29150 50990 29202
rect 51042 29150 51156 29202
rect 50988 29148 51156 29150
rect 50988 29138 51044 29148
rect 50988 28980 51044 28990
rect 50652 28644 50708 28654
rect 50652 28530 50708 28588
rect 50652 28478 50654 28530
rect 50706 28478 50708 28530
rect 50652 28466 50708 28478
rect 50988 28530 51044 28924
rect 50988 28478 50990 28530
rect 51042 28478 51044 28530
rect 50876 28420 50932 28430
rect 50876 28326 50932 28364
rect 50204 28252 50484 28308
rect 50556 28252 50820 28262
rect 49868 27692 50036 27748
rect 50092 28084 50148 28094
rect 49868 26514 49924 27692
rect 49868 26462 49870 26514
rect 49922 26462 49924 26514
rect 49868 26450 49924 26462
rect 49980 27076 50036 27086
rect 50092 27076 50148 28028
rect 50204 27972 50260 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50988 28084 51044 28478
rect 51100 28532 51156 29148
rect 51212 29110 51268 29148
rect 51324 29316 51380 30382
rect 51772 29540 51828 32620
rect 51772 29474 51828 29484
rect 51324 29202 51380 29260
rect 51324 29150 51326 29202
rect 51378 29150 51380 29202
rect 51100 28466 51156 28476
rect 51212 28530 51268 28542
rect 51212 28478 51214 28530
rect 51266 28478 51268 28530
rect 51212 28196 51268 28478
rect 51212 28130 51268 28140
rect 50988 28028 51156 28084
rect 50428 27972 50484 27982
rect 50204 27906 50260 27916
rect 50316 27970 50484 27972
rect 50316 27918 50430 27970
rect 50482 27918 50484 27970
rect 50316 27916 50484 27918
rect 50316 27860 50372 27916
rect 50428 27906 50484 27916
rect 50652 27970 50708 27982
rect 50652 27918 50654 27970
rect 50706 27918 50708 27970
rect 50316 27794 50372 27804
rect 49980 27074 50148 27076
rect 49980 27022 49982 27074
rect 50034 27022 50148 27074
rect 49980 27020 50148 27022
rect 50540 27746 50596 27758
rect 50540 27694 50542 27746
rect 50594 27694 50596 27746
rect 49084 26124 49588 26180
rect 49196 25844 49252 25854
rect 49196 25730 49252 25788
rect 49196 25678 49198 25730
rect 49250 25678 49252 25730
rect 49196 25666 49252 25678
rect 48972 25620 49028 25630
rect 48972 25394 49028 25564
rect 48972 25342 48974 25394
rect 49026 25342 49028 25394
rect 48972 25330 49028 25342
rect 49084 25396 49140 25406
rect 49084 25302 49140 25340
rect 48972 25060 49028 25070
rect 48972 23492 49028 25004
rect 49532 24948 49588 26124
rect 49756 26290 49812 26302
rect 49756 26238 49758 26290
rect 49810 26238 49812 26290
rect 49756 25956 49812 26238
rect 49756 25890 49812 25900
rect 49868 26292 49924 26302
rect 49868 25508 49924 26236
rect 49980 25732 50036 27020
rect 50428 26964 50484 26974
rect 50540 26908 50596 27694
rect 50092 26852 50148 26862
rect 50316 26852 50372 26862
rect 50092 26758 50148 26796
rect 50204 26850 50372 26852
rect 50204 26798 50318 26850
rect 50370 26798 50372 26850
rect 50204 26796 50372 26798
rect 50092 26404 50148 26414
rect 50092 26310 50148 26348
rect 50204 26292 50260 26796
rect 50316 26786 50372 26796
rect 50428 26852 50596 26908
rect 50652 27524 50708 27918
rect 50652 26852 50708 27468
rect 50764 27972 50820 27982
rect 50764 27186 50820 27916
rect 50764 27134 50766 27186
rect 50818 27134 50820 27186
rect 50764 27122 50820 27134
rect 50204 26226 50260 26236
rect 50316 26290 50372 26302
rect 50316 26238 50318 26290
rect 50370 26238 50372 26290
rect 50204 25844 50260 25854
rect 49980 25676 50148 25732
rect 49980 25508 50036 25518
rect 49868 25506 50036 25508
rect 49868 25454 49982 25506
rect 50034 25454 50036 25506
rect 49868 25452 50036 25454
rect 49980 25442 50036 25452
rect 49756 25394 49812 25406
rect 49756 25342 49758 25394
rect 49810 25342 49812 25394
rect 49756 25172 49812 25342
rect 49756 25106 49812 25116
rect 49868 25284 49924 25294
rect 49532 24892 49812 24948
rect 49532 24724 49588 24734
rect 49196 24722 49588 24724
rect 49196 24670 49534 24722
rect 49586 24670 49588 24722
rect 49196 24668 49588 24670
rect 49196 23548 49252 24668
rect 49532 24658 49588 24668
rect 49644 24724 49700 24734
rect 49308 24164 49364 24174
rect 49308 24070 49364 24108
rect 49644 23940 49700 24668
rect 49532 23884 49700 23940
rect 49420 23828 49476 23838
rect 49420 23734 49476 23772
rect 49532 23548 49588 23884
rect 49196 23492 49364 23548
rect 48972 23436 49140 23492
rect 49084 22820 49140 23436
rect 49532 23482 49588 23492
rect 49644 23716 49700 23726
rect 49756 23716 49812 24892
rect 49868 24722 49924 25228
rect 49868 24670 49870 24722
rect 49922 24670 49924 24722
rect 49868 24658 49924 24670
rect 50092 24164 50148 25676
rect 49644 23714 49812 23716
rect 49644 23662 49646 23714
rect 49698 23662 49812 23714
rect 49644 23660 49812 23662
rect 49868 24108 50148 24164
rect 49308 23426 49364 23436
rect 49644 23380 49700 23660
rect 49868 23548 49924 24108
rect 49980 23940 50036 23950
rect 49980 23938 50148 23940
rect 49980 23886 49982 23938
rect 50034 23886 50148 23938
rect 49980 23884 50148 23886
rect 49980 23874 50036 23884
rect 50092 23548 50148 23884
rect 49868 23492 50036 23548
rect 49532 23324 49700 23380
rect 49980 23380 50036 23492
rect 50092 23482 50148 23492
rect 50092 23380 50148 23390
rect 49980 23324 50092 23380
rect 49532 23266 49588 23324
rect 50092 23314 50148 23324
rect 49532 23214 49534 23266
rect 49586 23214 49588 23266
rect 49532 23202 49588 23214
rect 49756 23268 49812 23278
rect 49756 23174 49812 23212
rect 49084 22754 49140 22764
rect 49308 23154 49364 23166
rect 49308 23102 49310 23154
rect 49362 23102 49364 23154
rect 48860 22430 48862 22482
rect 48914 22430 48916 22482
rect 48860 22418 48916 22430
rect 48972 22372 49028 22382
rect 48972 21026 49028 22316
rect 48972 20974 48974 21026
rect 49026 20974 49028 21026
rect 48972 20962 49028 20974
rect 49084 20578 49140 20590
rect 49084 20526 49086 20578
rect 49138 20526 49140 20578
rect 49084 20468 49140 20526
rect 49084 20402 49140 20412
rect 49084 20132 49140 20142
rect 48860 20020 48916 20030
rect 48860 19926 48916 19964
rect 48748 19404 48916 19460
rect 48412 19292 48692 19348
rect 48300 18452 48356 18462
rect 48412 18452 48468 19292
rect 48748 19236 48804 19246
rect 48524 19180 48748 19236
rect 48524 18674 48580 19180
rect 48748 19104 48804 19180
rect 48524 18622 48526 18674
rect 48578 18622 48580 18674
rect 48524 18610 48580 18622
rect 48636 18788 48692 18798
rect 48636 18562 48692 18732
rect 48636 18510 48638 18562
rect 48690 18510 48692 18562
rect 48412 18396 48580 18452
rect 48300 17668 48356 18396
rect 48412 18228 48468 18238
rect 48412 18134 48468 18172
rect 48300 17602 48356 17612
rect 48412 17556 48468 17566
rect 48300 17444 48356 17454
rect 48412 17444 48468 17500
rect 48300 17442 48468 17444
rect 48300 17390 48302 17442
rect 48354 17390 48468 17442
rect 48300 17388 48468 17390
rect 48300 17378 48356 17388
rect 48188 16884 48244 16894
rect 48188 16790 48244 16828
rect 48412 16882 48468 17388
rect 48412 16830 48414 16882
rect 48466 16830 48468 16882
rect 48076 16706 48132 16716
rect 48300 16212 48356 16222
rect 48300 16118 48356 16156
rect 48412 15652 48468 16830
rect 48076 15596 48468 15652
rect 48524 15652 48580 18396
rect 48636 16996 48692 18510
rect 48748 17780 48804 17790
rect 48860 17780 48916 19404
rect 48972 19348 49028 19358
rect 48972 19254 49028 19292
rect 48804 17724 48916 17780
rect 49084 19234 49140 20076
rect 49084 19182 49086 19234
rect 49138 19182 49140 19234
rect 48748 17648 48804 17724
rect 49084 17108 49140 19182
rect 49196 18004 49252 18014
rect 49196 17778 49252 17948
rect 49196 17726 49198 17778
rect 49250 17726 49252 17778
rect 49196 17714 49252 17726
rect 49308 17444 49364 23102
rect 50092 23044 50148 23054
rect 49644 22932 49700 22942
rect 49644 22838 49700 22876
rect 49980 22930 50036 22942
rect 49980 22878 49982 22930
rect 50034 22878 50036 22930
rect 49980 22820 50036 22878
rect 49756 22372 49812 22382
rect 49644 22370 49812 22372
rect 49644 22318 49758 22370
rect 49810 22318 49812 22370
rect 49644 22316 49812 22318
rect 49420 21924 49476 21934
rect 49420 21810 49476 21868
rect 49420 21758 49422 21810
rect 49474 21758 49476 21810
rect 49420 21746 49476 21758
rect 49644 21812 49700 22316
rect 49756 22306 49812 22316
rect 49644 21746 49700 21756
rect 49756 22148 49812 22158
rect 49644 21364 49700 21374
rect 49420 21026 49476 21038
rect 49420 20974 49422 21026
rect 49474 20974 49476 21026
rect 49420 20580 49476 20974
rect 49532 20580 49588 20590
rect 49420 20578 49588 20580
rect 49420 20526 49534 20578
rect 49586 20526 49588 20578
rect 49420 20524 49588 20526
rect 49532 19796 49588 20524
rect 49532 19730 49588 19740
rect 49532 19124 49588 19134
rect 49532 18674 49588 19068
rect 49532 18622 49534 18674
rect 49586 18622 49588 18674
rect 49532 18610 49588 18622
rect 49532 18452 49588 18462
rect 49308 17378 49364 17388
rect 49420 18340 49476 18350
rect 49084 17042 49140 17052
rect 48636 16940 48804 16996
rect 48524 15596 48692 15652
rect 48076 14754 48132 15596
rect 48188 15428 48244 15438
rect 48188 15334 48244 15372
rect 48524 15426 48580 15438
rect 48524 15374 48526 15426
rect 48578 15374 48580 15426
rect 48524 15204 48580 15374
rect 48524 15138 48580 15148
rect 48076 14702 48078 14754
rect 48130 14702 48132 14754
rect 48076 13300 48132 14702
rect 48412 14756 48468 14766
rect 48188 14644 48244 14654
rect 48188 14550 48244 14588
rect 48188 14308 48244 14318
rect 48188 13524 48244 14252
rect 48412 13970 48468 14700
rect 48636 14308 48692 15596
rect 48748 15204 48804 16940
rect 49308 16212 49364 16222
rect 49308 16098 49364 16156
rect 49308 16046 49310 16098
rect 49362 16046 49364 16098
rect 49308 16034 49364 16046
rect 48972 15876 49028 15886
rect 48972 15782 49028 15820
rect 49084 15874 49140 15886
rect 49084 15822 49086 15874
rect 49138 15822 49140 15874
rect 48748 15138 48804 15148
rect 48748 14756 48804 14766
rect 48748 14642 48804 14700
rect 48748 14590 48750 14642
rect 48802 14590 48804 14642
rect 48748 14578 48804 14590
rect 48636 14242 48692 14252
rect 48972 14532 49028 14542
rect 48412 13918 48414 13970
rect 48466 13918 48468 13970
rect 48412 13906 48468 13918
rect 48188 13458 48244 13468
rect 48748 13746 48804 13758
rect 48748 13694 48750 13746
rect 48802 13694 48804 13746
rect 48076 13244 48244 13300
rect 47964 13132 48132 13188
rect 47964 12964 48020 12974
rect 47964 12870 48020 12908
rect 47852 12460 48020 12516
rect 47740 12338 47796 12348
rect 47852 12292 47908 12302
rect 47740 12068 47796 12078
rect 47740 11974 47796 12012
rect 47628 11508 47684 11518
rect 47628 11414 47684 11452
rect 47740 11060 47796 11070
rect 47404 9214 47406 9266
rect 47458 9214 47460 9266
rect 46620 7476 46676 9212
rect 46844 9202 46900 9212
rect 47404 9202 47460 9214
rect 47628 10948 47684 10958
rect 47292 7700 47348 7710
rect 47292 7606 47348 7644
rect 45948 6692 46004 6702
rect 45948 6598 46004 6636
rect 46508 6132 46564 6142
rect 46620 6132 46676 7420
rect 46508 6130 46676 6132
rect 46508 6078 46510 6130
rect 46562 6078 46676 6130
rect 46508 6076 46676 6078
rect 46956 7588 47012 7598
rect 46956 6130 47012 7532
rect 46956 6078 46958 6130
rect 47010 6078 47012 6130
rect 46508 6066 46564 6076
rect 46956 6066 47012 6078
rect 47068 6692 47124 6702
rect 45948 6020 46004 6030
rect 45948 6018 46116 6020
rect 45948 5966 45950 6018
rect 46002 5966 46116 6018
rect 45948 5964 46116 5966
rect 45948 5954 46004 5964
rect 45948 5122 46004 5134
rect 45948 5070 45950 5122
rect 46002 5070 46004 5122
rect 45948 4564 46004 5070
rect 45948 4498 46004 4508
rect 46060 3892 46116 5964
rect 46732 5012 46788 5022
rect 46732 4226 46788 4956
rect 46732 4174 46734 4226
rect 46786 4174 46788 4226
rect 46172 3892 46228 3902
rect 46060 3836 46172 3892
rect 45836 3614 45838 3666
rect 45890 3614 45892 3666
rect 45836 3602 45892 3614
rect 46172 3666 46228 3836
rect 46172 3614 46174 3666
rect 46226 3614 46228 3666
rect 46172 3602 46228 3614
rect 46732 3668 46788 4174
rect 46732 3574 46788 3612
rect 47068 3666 47124 6636
rect 47628 6132 47684 10892
rect 47740 7700 47796 11004
rect 47852 9266 47908 12236
rect 47964 11508 48020 12460
rect 48076 11732 48132 13132
rect 48076 11666 48132 11676
rect 47964 11506 48132 11508
rect 47964 11454 47966 11506
rect 48018 11454 48132 11506
rect 47964 11452 48132 11454
rect 47964 11442 48020 11452
rect 47964 10834 48020 10846
rect 47964 10782 47966 10834
rect 48018 10782 48020 10834
rect 47964 9940 48020 10782
rect 47964 9874 48020 9884
rect 48076 9716 48132 11452
rect 48076 9650 48132 9660
rect 47852 9214 47854 9266
rect 47906 9214 47908 9266
rect 47852 9202 47908 9214
rect 48188 9044 48244 13244
rect 48300 13188 48356 13198
rect 48748 13188 48804 13694
rect 48300 13186 48804 13188
rect 48300 13134 48302 13186
rect 48354 13134 48804 13186
rect 48300 13132 48804 13134
rect 48300 13122 48356 13132
rect 48636 12964 48692 12974
rect 48636 12292 48692 12908
rect 48748 12852 48804 13132
rect 48860 13300 48916 13310
rect 48972 13300 49028 14476
rect 49084 13860 49140 15822
rect 49308 15652 49364 15662
rect 49308 15428 49364 15596
rect 49308 15362 49364 15372
rect 49420 15202 49476 18284
rect 49532 16436 49588 18396
rect 49644 18004 49700 21308
rect 49756 21252 49812 22092
rect 49756 21186 49812 21196
rect 49980 20804 50036 22764
rect 49868 20748 50036 20804
rect 49868 20356 49924 20748
rect 49980 20580 50036 20590
rect 49980 20486 50036 20524
rect 49868 20300 50036 20356
rect 49756 20132 49812 20142
rect 49756 20018 49812 20076
rect 49756 19966 49758 20018
rect 49810 19966 49812 20018
rect 49756 18676 49812 19966
rect 49868 19236 49924 19246
rect 49868 19142 49924 19180
rect 49868 18676 49924 18686
rect 49756 18674 49924 18676
rect 49756 18622 49870 18674
rect 49922 18622 49924 18674
rect 49756 18620 49924 18622
rect 49644 17948 49812 18004
rect 49644 17780 49700 17790
rect 49644 17686 49700 17724
rect 49644 16996 49700 17006
rect 49644 16902 49700 16940
rect 49756 16772 49812 17948
rect 49868 17668 49924 18620
rect 49980 18340 50036 20300
rect 49980 18274 50036 18284
rect 49868 17602 49924 17612
rect 49980 17556 50036 17566
rect 49980 16882 50036 17500
rect 49980 16830 49982 16882
rect 50034 16830 50036 16882
rect 49980 16818 50036 16830
rect 49756 16770 49924 16772
rect 49756 16718 49758 16770
rect 49810 16718 49924 16770
rect 49756 16716 49924 16718
rect 49756 16706 49812 16716
rect 49532 16370 49588 16380
rect 49644 16100 49700 16110
rect 49644 16006 49700 16044
rect 49420 15150 49422 15202
rect 49474 15150 49476 15202
rect 49420 15148 49476 15150
rect 49420 15092 49812 15148
rect 49420 14418 49476 14430
rect 49420 14366 49422 14418
rect 49474 14366 49476 14418
rect 49420 14196 49476 14366
rect 49532 14308 49588 14318
rect 49532 14214 49588 14252
rect 49644 14306 49700 14318
rect 49644 14254 49646 14306
rect 49698 14254 49700 14306
rect 49420 14130 49476 14140
rect 49084 13794 49140 13804
rect 49644 13860 49700 14254
rect 49644 13794 49700 13804
rect 49644 13634 49700 13646
rect 49644 13582 49646 13634
rect 49698 13582 49700 13634
rect 48972 13244 49140 13300
rect 48860 13076 48916 13244
rect 48972 13076 49028 13086
rect 48860 13020 48972 13076
rect 48972 12982 49028 13020
rect 48748 12786 48804 12796
rect 48748 12516 48804 12526
rect 48748 12402 48804 12460
rect 48748 12350 48750 12402
rect 48802 12350 48804 12402
rect 48748 12338 48804 12350
rect 48524 12290 48692 12292
rect 48524 12238 48638 12290
rect 48690 12238 48692 12290
rect 48524 12236 48692 12238
rect 48524 11282 48580 12236
rect 48636 12226 48692 12236
rect 48524 11230 48526 11282
rect 48578 11230 48580 11282
rect 48524 11218 48580 11230
rect 48636 11732 48692 11742
rect 48524 10388 48580 10398
rect 48524 10294 48580 10332
rect 48636 10164 48692 11676
rect 48860 11284 48916 11294
rect 49084 11284 49140 13244
rect 49532 13076 49588 13086
rect 49644 13076 49700 13582
rect 49756 13412 49812 15092
rect 49868 13636 49924 16716
rect 50092 16212 50148 22988
rect 50204 22370 50260 25788
rect 50316 24724 50372 26238
rect 50316 24658 50372 24668
rect 50428 24722 50484 26852
rect 50652 26786 50708 26796
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 51100 26628 51156 28028
rect 51212 27746 51268 27758
rect 51212 27694 51214 27746
rect 51266 27694 51268 27746
rect 51212 27076 51268 27694
rect 51212 27010 51268 27020
rect 51324 26964 51380 29150
rect 51660 28644 51716 28654
rect 51324 26898 51380 26908
rect 51548 27074 51604 27086
rect 51548 27022 51550 27074
rect 51602 27022 51604 27074
rect 50764 26516 50820 26526
rect 50764 26422 50820 26460
rect 51100 26292 51156 26572
rect 51100 26226 51156 26236
rect 51324 26740 51380 26750
rect 51212 26178 51268 26190
rect 51212 26126 51214 26178
rect 51266 26126 51268 26178
rect 51100 26066 51156 26078
rect 51100 26014 51102 26066
rect 51154 26014 51156 26066
rect 51100 25618 51156 26014
rect 51212 26068 51268 26126
rect 51212 26002 51268 26012
rect 51100 25566 51102 25618
rect 51154 25566 51156 25618
rect 51100 25554 51156 25566
rect 51212 25508 51268 25518
rect 51212 25414 51268 25452
rect 50764 25396 50820 25406
rect 50764 25394 50932 25396
rect 50764 25342 50766 25394
rect 50818 25342 50932 25394
rect 50764 25340 50932 25342
rect 50764 25330 50820 25340
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50876 24834 50932 25340
rect 51324 25284 51380 26684
rect 51548 25732 51604 27022
rect 51660 26404 51716 28588
rect 51772 28530 51828 28542
rect 51772 28478 51774 28530
rect 51826 28478 51828 28530
rect 51772 28420 51828 28478
rect 51772 28354 51828 28364
rect 51884 28196 51940 33740
rect 52108 31892 52164 35308
rect 52332 34804 52388 36764
rect 52444 36708 52500 40012
rect 52556 39732 52612 40124
rect 52668 39844 52724 40908
rect 52780 40964 52836 40974
rect 52780 40962 53060 40964
rect 52780 40910 52782 40962
rect 52834 40910 53060 40962
rect 52780 40908 53060 40910
rect 52780 40898 52836 40908
rect 52892 40740 52948 40750
rect 52780 39844 52836 39854
rect 52668 39842 52836 39844
rect 52668 39790 52782 39842
rect 52834 39790 52836 39842
rect 52668 39788 52836 39790
rect 52780 39778 52836 39788
rect 52556 39676 52724 39732
rect 52444 36642 52500 36652
rect 52556 38724 52612 38734
rect 52444 36372 52500 36382
rect 52444 36278 52500 36316
rect 52556 35476 52612 38668
rect 52668 37490 52724 39676
rect 52780 38276 52836 38286
rect 52780 38182 52836 38220
rect 52892 38052 52948 40684
rect 52892 37986 52948 37996
rect 52668 37438 52670 37490
rect 52722 37438 52724 37490
rect 52668 37426 52724 37438
rect 52780 37716 52836 37726
rect 52780 37266 52836 37660
rect 53004 37492 53060 40908
rect 52780 37214 52782 37266
rect 52834 37214 52836 37266
rect 52780 37202 52836 37214
rect 52892 37436 53060 37492
rect 53116 40516 53172 40526
rect 52668 36596 52724 36606
rect 52668 36482 52724 36540
rect 52668 36430 52670 36482
rect 52722 36430 52724 36482
rect 52668 36418 52724 36430
rect 52668 35924 52724 35934
rect 52668 35830 52724 35868
rect 52892 35698 52948 37436
rect 53004 37268 53060 37278
rect 53116 37268 53172 40460
rect 53228 40404 53284 40414
rect 53228 40310 53284 40348
rect 53340 38668 53396 41020
rect 53452 40068 53508 44270
rect 53676 44322 53732 44334
rect 53676 44270 53678 44322
rect 53730 44270 53732 44322
rect 53676 44212 53732 44270
rect 53676 44146 53732 44156
rect 53452 40002 53508 40012
rect 53564 43540 53620 43550
rect 53452 39394 53508 39406
rect 53452 39342 53454 39394
rect 53506 39342 53508 39394
rect 53452 39060 53508 39342
rect 53452 38994 53508 39004
rect 53564 38668 53620 43484
rect 53676 43204 53732 43214
rect 53676 42644 53732 43148
rect 53788 42756 53844 45054
rect 53900 44322 53956 44334
rect 53900 44270 53902 44322
rect 53954 44270 53956 44322
rect 53900 43876 53956 44270
rect 53900 43810 53956 43820
rect 54012 44324 54068 44334
rect 53900 43538 53956 43550
rect 53900 43486 53902 43538
rect 53954 43486 53956 43538
rect 53900 43316 53956 43486
rect 53900 43250 53956 43260
rect 54012 42978 54068 44268
rect 54124 43764 54180 45612
rect 54236 45602 54292 45612
rect 54460 45444 54516 45454
rect 54460 45106 54516 45388
rect 54460 45054 54462 45106
rect 54514 45054 54516 45106
rect 54460 45042 54516 45054
rect 54236 44882 54292 44894
rect 54236 44830 54238 44882
rect 54290 44830 54292 44882
rect 54236 44548 54292 44830
rect 54460 44884 54516 44894
rect 54572 44884 54628 47180
rect 54516 44828 54628 44884
rect 54684 46674 54740 48076
rect 54796 48130 54852 48142
rect 54796 48078 54798 48130
rect 54850 48078 54852 48130
rect 54796 48020 54852 48078
rect 55244 48132 55300 48142
rect 55244 48130 55412 48132
rect 55244 48078 55246 48130
rect 55298 48078 55412 48130
rect 55244 48076 55412 48078
rect 55244 48066 55300 48076
rect 54796 47964 55076 48020
rect 54908 47348 54964 47358
rect 54908 47254 54964 47292
rect 54684 46622 54686 46674
rect 54738 46622 54740 46674
rect 54348 44548 54404 44558
rect 54236 44546 54404 44548
rect 54236 44494 54350 44546
rect 54402 44494 54404 44546
rect 54236 44492 54404 44494
rect 54348 44482 54404 44492
rect 54124 43708 54292 43764
rect 54012 42926 54014 42978
rect 54066 42926 54068 42978
rect 54012 42914 54068 42926
rect 54124 43538 54180 43550
rect 54124 43486 54126 43538
rect 54178 43486 54180 43538
rect 54012 42756 54068 42766
rect 53788 42700 53956 42756
rect 53676 42588 53844 42644
rect 53676 41858 53732 41870
rect 53676 41806 53678 41858
rect 53730 41806 53732 41858
rect 53676 39172 53732 41806
rect 53788 41074 53844 42588
rect 53900 41860 53956 42700
rect 54012 42642 54068 42700
rect 54012 42590 54014 42642
rect 54066 42590 54068 42642
rect 54012 42578 54068 42590
rect 54124 42644 54180 43486
rect 54236 42756 54292 43708
rect 54348 43652 54404 43662
rect 54460 43652 54516 44828
rect 54684 44212 54740 46622
rect 54796 45668 54852 45678
rect 54796 45574 54852 45612
rect 54684 44146 54740 44156
rect 54908 45332 54964 45342
rect 55020 45332 55076 47964
rect 55244 47684 55300 47694
rect 55244 47346 55300 47628
rect 55244 47294 55246 47346
rect 55298 47294 55300 47346
rect 55244 47282 55300 47294
rect 55356 47236 55412 48076
rect 55356 47170 55412 47180
rect 55468 46788 55524 48748
rect 56028 48468 56084 48862
rect 56028 48402 56084 48412
rect 55356 46564 55412 46574
rect 55356 46470 55412 46508
rect 55244 45668 55300 45678
rect 55244 45666 55412 45668
rect 55244 45614 55246 45666
rect 55298 45614 55412 45666
rect 55244 45612 55412 45614
rect 55244 45602 55300 45612
rect 54964 45276 55076 45332
rect 54908 44436 54964 45276
rect 54348 43650 54516 43652
rect 54348 43598 54350 43650
rect 54402 43598 54516 43650
rect 54348 43596 54516 43598
rect 54348 43092 54404 43596
rect 54348 43026 54404 43036
rect 54460 43314 54516 43326
rect 54460 43262 54462 43314
rect 54514 43262 54516 43314
rect 54460 42756 54516 43262
rect 54572 42756 54628 42766
rect 54236 42700 54404 42756
rect 54460 42754 54628 42756
rect 54460 42702 54574 42754
rect 54626 42702 54628 42754
rect 54460 42700 54628 42702
rect 54124 42642 54292 42644
rect 54124 42590 54126 42642
rect 54178 42590 54292 42642
rect 54124 42588 54292 42590
rect 54124 42578 54180 42588
rect 53900 41804 54068 41860
rect 53788 41022 53790 41074
rect 53842 41022 53844 41074
rect 53788 40068 53844 41022
rect 53788 40002 53844 40012
rect 53900 39956 53956 39966
rect 53788 39396 53844 39406
rect 53788 39302 53844 39340
rect 53676 39106 53732 39116
rect 53676 38836 53732 38846
rect 53676 38742 53732 38780
rect 53340 38612 53508 38668
rect 53564 38612 53732 38668
rect 53340 38388 53396 38398
rect 53340 38162 53396 38332
rect 53340 38110 53342 38162
rect 53394 38110 53396 38162
rect 53340 38098 53396 38110
rect 53060 37212 53172 37268
rect 53228 37380 53284 37390
rect 53004 37174 53060 37212
rect 52892 35646 52894 35698
rect 52946 35646 52948 35698
rect 52556 35420 52724 35476
rect 52220 34748 52388 34804
rect 52556 35252 52612 35262
rect 52220 32228 52276 34748
rect 52444 34692 52500 34702
rect 52332 34690 52500 34692
rect 52332 34638 52446 34690
rect 52498 34638 52500 34690
rect 52332 34636 52500 34638
rect 52332 34356 52388 34636
rect 52444 34626 52500 34636
rect 52332 34290 52388 34300
rect 52444 34356 52500 34366
rect 52556 34356 52612 35196
rect 52444 34354 52612 34356
rect 52444 34302 52446 34354
rect 52498 34302 52612 34354
rect 52444 34300 52612 34302
rect 52444 34290 52500 34300
rect 52668 33348 52724 35420
rect 52892 34692 52948 35646
rect 52892 34626 52948 34636
rect 53004 36932 53060 36942
rect 52780 34244 52836 34254
rect 52780 34150 52836 34188
rect 52556 33292 52724 33348
rect 52892 33572 52948 33582
rect 52332 33124 52388 33134
rect 52332 33030 52388 33068
rect 52332 32900 52388 32910
rect 52332 32452 52388 32844
rect 52332 32386 52388 32396
rect 52444 32450 52500 32462
rect 52444 32398 52446 32450
rect 52498 32398 52500 32450
rect 52220 32172 52388 32228
rect 52108 31836 52276 31892
rect 51996 31778 52052 31790
rect 51996 31726 51998 31778
rect 52050 31726 52052 31778
rect 51996 31332 52052 31726
rect 52220 31780 52276 31836
rect 52220 31714 52276 31724
rect 52220 31554 52276 31566
rect 52220 31502 52222 31554
rect 52274 31502 52276 31554
rect 52220 31444 52276 31502
rect 51996 31266 52052 31276
rect 52108 31388 52276 31444
rect 52108 30436 52164 31388
rect 52332 31332 52388 32172
rect 52444 32004 52500 32398
rect 52444 31938 52500 31948
rect 52444 31780 52500 31790
rect 52556 31780 52612 33292
rect 52668 33124 52724 33134
rect 52668 33030 52724 33068
rect 52892 32786 52948 33516
rect 52892 32734 52894 32786
rect 52946 32734 52948 32786
rect 52892 32722 52948 32734
rect 52444 31778 52612 31780
rect 52444 31726 52446 31778
rect 52498 31726 52612 31778
rect 52444 31724 52612 31726
rect 52444 31714 52500 31724
rect 51996 30380 52164 30436
rect 52220 31276 52388 31332
rect 51996 30212 52052 30380
rect 52220 30324 52276 31276
rect 51996 30146 52052 30156
rect 52108 30268 52276 30324
rect 52332 31108 52388 31118
rect 51996 28644 52052 28654
rect 51996 28530 52052 28588
rect 51996 28478 51998 28530
rect 52050 28478 52052 28530
rect 51996 28466 52052 28478
rect 52108 28530 52164 30268
rect 52332 29764 52388 31052
rect 52556 30660 52612 31724
rect 52668 31780 52724 31790
rect 52668 31686 52724 31724
rect 53004 31332 53060 36876
rect 53116 34132 53172 34142
rect 53116 33124 53172 34076
rect 53116 33058 53172 33068
rect 53004 31266 53060 31276
rect 53116 31220 53172 31230
rect 53116 31126 53172 31164
rect 52556 30604 52836 30660
rect 52556 30436 52612 30446
rect 52556 30342 52612 30380
rect 52444 30210 52500 30222
rect 52444 30158 52446 30210
rect 52498 30158 52500 30210
rect 52444 30100 52500 30158
rect 52500 30044 52612 30100
rect 52444 30034 52500 30044
rect 52332 29314 52388 29708
rect 52332 29262 52334 29314
rect 52386 29262 52388 29314
rect 52332 29250 52388 29262
rect 52444 29316 52500 29326
rect 52556 29316 52612 30044
rect 52556 29260 52724 29316
rect 52332 28644 52388 28654
rect 52108 28478 52110 28530
rect 52162 28478 52164 28530
rect 52108 28466 52164 28478
rect 52220 28642 52388 28644
rect 52220 28590 52334 28642
rect 52386 28590 52388 28642
rect 52220 28588 52388 28590
rect 51660 26338 51716 26348
rect 51772 28140 51940 28196
rect 51996 28308 52052 28318
rect 51660 26180 51716 26190
rect 51660 26086 51716 26124
rect 51772 26066 51828 28140
rect 51884 27972 51940 27982
rect 51884 27878 51940 27916
rect 51884 27300 51940 27338
rect 51884 27234 51940 27244
rect 51772 26014 51774 26066
rect 51826 26014 51828 26066
rect 51772 26002 51828 26014
rect 51884 27074 51940 27086
rect 51884 27022 51886 27074
rect 51938 27022 51940 27074
rect 51660 25732 51716 25742
rect 51548 25730 51716 25732
rect 51548 25678 51662 25730
rect 51714 25678 51716 25730
rect 51548 25676 51716 25678
rect 51660 25666 51716 25676
rect 51884 25620 51940 27022
rect 51996 26180 52052 28252
rect 52108 27970 52164 27982
rect 52108 27918 52110 27970
rect 52162 27918 52164 27970
rect 52108 27636 52164 27918
rect 52220 27746 52276 28588
rect 52332 28578 52388 28588
rect 52220 27694 52222 27746
rect 52274 27694 52276 27746
rect 52220 27682 52276 27694
rect 52108 27076 52164 27580
rect 52444 27412 52500 29260
rect 52108 26514 52164 27020
rect 52108 26462 52110 26514
rect 52162 26462 52164 26514
rect 52108 26450 52164 26462
rect 52220 27356 52500 27412
rect 52556 28642 52612 28654
rect 52556 28590 52558 28642
rect 52610 28590 52612 28642
rect 51996 26114 52052 26124
rect 51772 25564 51884 25620
rect 51324 25218 51380 25228
rect 51660 25284 51716 25294
rect 50876 24782 50878 24834
rect 50930 24782 50932 24834
rect 50876 24770 50932 24782
rect 50428 24670 50430 24722
rect 50482 24670 50484 24722
rect 50428 24658 50484 24670
rect 51100 24724 51156 24734
rect 51100 24630 51156 24668
rect 51212 24722 51268 24734
rect 51212 24670 51214 24722
rect 51266 24670 51268 24722
rect 50764 24612 50820 24622
rect 50204 22318 50206 22370
rect 50258 22318 50260 22370
rect 50204 21812 50260 22318
rect 50316 24388 50372 24398
rect 50316 22372 50372 24332
rect 50764 24162 50820 24556
rect 50764 24110 50766 24162
rect 50818 24110 50820 24162
rect 50764 24098 50820 24110
rect 50876 24052 50932 24062
rect 50540 23828 50596 23838
rect 50540 23734 50596 23772
rect 50316 22306 50372 22316
rect 50428 23716 50484 23726
rect 50428 22148 50484 23660
rect 50652 23716 50708 23754
rect 50652 23650 50708 23660
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50652 23266 50708 23278
rect 50652 23214 50654 23266
rect 50706 23214 50708 23266
rect 50540 23044 50596 23054
rect 50540 22260 50596 22988
rect 50652 22484 50708 23214
rect 50652 22418 50708 22428
rect 50540 22194 50596 22204
rect 50764 22260 50820 22270
rect 50764 22166 50820 22204
rect 50428 22082 50484 22092
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50540 21812 50596 21850
rect 50876 21812 50932 23996
rect 51100 23380 51156 23390
rect 50204 21756 50484 21812
rect 50316 21586 50372 21598
rect 50316 21534 50318 21586
rect 50370 21534 50372 21586
rect 50316 20916 50372 21534
rect 50428 21026 50484 21756
rect 50540 21746 50596 21756
rect 50764 21756 50932 21812
rect 50988 23154 51044 23166
rect 50988 23102 50990 23154
rect 51042 23102 51044 23154
rect 50988 22036 51044 23102
rect 50988 21812 51044 21980
rect 50540 21588 50596 21598
rect 50540 21494 50596 21532
rect 50428 20974 50430 21026
rect 50482 20974 50484 21026
rect 50428 20962 50484 20974
rect 50764 21028 50820 21756
rect 50988 21746 51044 21756
rect 50876 21588 50932 21598
rect 50876 21494 50932 21532
rect 51100 21476 51156 23324
rect 51212 22596 51268 24670
rect 51548 24052 51604 24062
rect 51548 23938 51604 23996
rect 51548 23886 51550 23938
rect 51602 23886 51604 23938
rect 51548 23874 51604 23886
rect 51548 23492 51604 23502
rect 51548 23378 51604 23436
rect 51548 23326 51550 23378
rect 51602 23326 51604 23378
rect 51548 23314 51604 23326
rect 51212 22530 51268 22540
rect 51324 23156 51380 23166
rect 51324 22594 51380 23100
rect 51324 22542 51326 22594
rect 51378 22542 51380 22594
rect 51324 22530 51380 22542
rect 51548 22596 51604 22606
rect 51100 21410 51156 21420
rect 51212 22372 51268 22382
rect 50204 20860 50372 20916
rect 50764 20916 50820 20972
rect 50988 21252 51044 21262
rect 50876 20916 50932 20926
rect 50764 20914 50932 20916
rect 50764 20862 50878 20914
rect 50930 20862 50932 20914
rect 50764 20860 50932 20862
rect 50204 20020 50260 20860
rect 50876 20850 50932 20860
rect 50316 20690 50372 20702
rect 50316 20638 50318 20690
rect 50370 20638 50372 20690
rect 50316 20244 50372 20638
rect 50428 20580 50484 20590
rect 50988 20580 51044 21196
rect 50428 20578 51044 20580
rect 50428 20526 50430 20578
rect 50482 20526 51044 20578
rect 50428 20524 51044 20526
rect 50428 20514 50484 20524
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50316 20188 50596 20244
rect 50316 20020 50372 20030
rect 50204 19964 50316 20020
rect 50316 19926 50372 19964
rect 50540 19906 50596 20188
rect 50540 19854 50542 19906
rect 50594 19854 50596 19906
rect 50540 19236 50596 19854
rect 50764 20020 50820 20030
rect 50652 19796 50708 19806
rect 50652 19702 50708 19740
rect 50540 19170 50596 19180
rect 50652 19348 50708 19358
rect 50764 19348 50820 19964
rect 50652 19346 50820 19348
rect 50652 19294 50654 19346
rect 50706 19294 50820 19346
rect 50652 19292 50820 19294
rect 50204 19124 50260 19134
rect 50204 19010 50260 19068
rect 50652 19124 50708 19292
rect 50652 19058 50708 19068
rect 50988 19236 51044 19246
rect 50204 18958 50206 19010
rect 50258 18958 50260 19010
rect 50204 18900 50260 18958
rect 50204 18834 50260 18844
rect 50556 18844 50820 18854
rect 50316 18788 50372 18798
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50316 18674 50372 18732
rect 50316 18622 50318 18674
rect 50370 18622 50372 18674
rect 50316 18610 50372 18622
rect 50876 18564 50932 18574
rect 50764 18340 50820 18350
rect 50764 18246 50820 18284
rect 50316 17892 50372 17902
rect 50204 17890 50372 17892
rect 50204 17838 50318 17890
rect 50370 17838 50372 17890
rect 50204 17836 50372 17838
rect 50204 17332 50260 17836
rect 50316 17826 50372 17836
rect 50876 17780 50932 18508
rect 50988 17892 51044 19180
rect 51212 19012 51268 22316
rect 51436 22370 51492 22382
rect 51436 22318 51438 22370
rect 51490 22318 51492 22370
rect 51436 22036 51492 22318
rect 51436 21970 51492 21980
rect 51548 21812 51604 22540
rect 51660 22036 51716 25228
rect 51772 23828 51828 25564
rect 51884 25554 51940 25564
rect 51996 25730 52052 25742
rect 51996 25678 51998 25730
rect 52050 25678 52052 25730
rect 51884 25284 51940 25294
rect 51996 25284 52052 25678
rect 51884 25282 52052 25284
rect 51884 25230 51886 25282
rect 51938 25230 52052 25282
rect 51884 25228 52052 25230
rect 51884 25218 51940 25228
rect 51884 23828 51940 23838
rect 51772 23826 51940 23828
rect 51772 23774 51886 23826
rect 51938 23774 51940 23826
rect 51772 23772 51940 23774
rect 51772 22372 51828 23772
rect 51884 23762 51940 23772
rect 51884 23044 51940 23054
rect 51884 22950 51940 22988
rect 51996 22484 52052 25228
rect 52220 23548 52276 27356
rect 52332 27188 52388 27198
rect 52332 27094 52388 27132
rect 52332 25620 52388 25630
rect 52332 25526 52388 25564
rect 52444 25284 52500 25294
rect 52332 25060 52388 25070
rect 52332 24388 52388 25004
rect 52332 24050 52388 24332
rect 52332 23998 52334 24050
rect 52386 23998 52388 24050
rect 52332 23986 52388 23998
rect 52444 24834 52500 25228
rect 52556 24946 52612 28590
rect 52556 24894 52558 24946
rect 52610 24894 52612 24946
rect 52556 24882 52612 24894
rect 52444 24782 52446 24834
rect 52498 24782 52500 24834
rect 52220 23492 52388 23548
rect 51996 22418 52052 22428
rect 52108 22708 52164 22718
rect 51772 22316 51940 22372
rect 51660 21970 51716 21980
rect 51772 22146 51828 22158
rect 51772 22094 51774 22146
rect 51826 22094 51828 22146
rect 51324 21756 51604 21812
rect 51772 21812 51828 22094
rect 51884 21812 51940 22316
rect 52108 22370 52164 22652
rect 52108 22318 52110 22370
rect 52162 22318 52164 22370
rect 52108 22306 52164 22318
rect 52332 22372 52388 23492
rect 52444 23492 52500 24782
rect 52444 23436 52612 23492
rect 52444 23268 52500 23278
rect 52444 23174 52500 23212
rect 52332 22278 52388 22316
rect 51996 22258 52052 22270
rect 51996 22206 51998 22258
rect 52050 22206 52052 22258
rect 51996 22036 52052 22206
rect 51996 21970 52052 21980
rect 52444 22260 52500 22270
rect 51884 21756 52052 21812
rect 51324 19908 51380 21756
rect 51772 21746 51828 21756
rect 51660 21698 51716 21710
rect 51660 21646 51662 21698
rect 51714 21646 51716 21698
rect 51660 21476 51716 21646
rect 51884 21586 51940 21598
rect 51884 21534 51886 21586
rect 51938 21534 51940 21586
rect 51548 21420 51716 21476
rect 51772 21474 51828 21486
rect 51772 21422 51774 21474
rect 51826 21422 51828 21474
rect 51436 21028 51492 21038
rect 51436 20692 51492 20972
rect 51548 20916 51604 21420
rect 51772 21364 51828 21422
rect 51772 21298 51828 21308
rect 51884 20916 51940 21534
rect 51548 20850 51604 20860
rect 51660 20860 51940 20916
rect 51660 20804 51716 20860
rect 51548 20692 51604 20702
rect 51436 20690 51604 20692
rect 51436 20638 51550 20690
rect 51602 20638 51604 20690
rect 51436 20636 51604 20638
rect 51548 20626 51604 20636
rect 51548 20244 51604 20254
rect 51660 20244 51716 20748
rect 51884 20690 51940 20702
rect 51884 20638 51886 20690
rect 51938 20638 51940 20690
rect 51548 20242 51716 20244
rect 51548 20190 51550 20242
rect 51602 20190 51716 20242
rect 51548 20188 51716 20190
rect 51772 20578 51828 20590
rect 51772 20526 51774 20578
rect 51826 20526 51828 20578
rect 51548 20178 51604 20188
rect 51772 20132 51828 20526
rect 51884 20244 51940 20638
rect 51884 20178 51940 20188
rect 51772 20066 51828 20076
rect 51884 20020 51940 20030
rect 51884 19926 51940 19964
rect 51324 19852 51716 19908
rect 51548 19684 51604 19694
rect 51436 19236 51492 19246
rect 51436 19142 51492 19180
rect 51548 19124 51604 19628
rect 51660 19348 51716 19852
rect 51660 19346 51828 19348
rect 51660 19294 51662 19346
rect 51714 19294 51828 19346
rect 51660 19292 51828 19294
rect 51660 19282 51716 19292
rect 51212 18956 51492 19012
rect 51324 18788 51380 18798
rect 51324 18564 51380 18732
rect 51324 18498 51380 18508
rect 51436 18452 51492 18956
rect 51548 18674 51604 19068
rect 51548 18622 51550 18674
rect 51602 18622 51604 18674
rect 51548 18610 51604 18622
rect 51436 18396 51716 18452
rect 50988 17836 51156 17892
rect 50876 17778 51044 17780
rect 50876 17726 50878 17778
rect 50930 17726 51044 17778
rect 50876 17724 51044 17726
rect 50876 17714 50932 17724
rect 50204 17266 50260 17276
rect 50316 17668 50372 17678
rect 50316 16770 50372 17612
rect 50428 17444 50484 17454
rect 50428 17350 50484 17388
rect 50876 17444 50932 17454
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50540 16884 50596 16894
rect 50540 16790 50596 16828
rect 50316 16718 50318 16770
rect 50370 16718 50372 16770
rect 50316 16660 50372 16718
rect 50316 16604 50484 16660
rect 50204 16212 50260 16222
rect 49980 16210 50260 16212
rect 49980 16158 50206 16210
rect 50258 16158 50260 16210
rect 49980 16156 50260 16158
rect 49980 13748 50036 16156
rect 50204 16146 50260 16156
rect 50092 15874 50148 15886
rect 50092 15822 50094 15874
rect 50146 15822 50148 15874
rect 50092 15540 50148 15822
rect 50316 15874 50372 15886
rect 50316 15822 50318 15874
rect 50370 15822 50372 15874
rect 50316 15764 50372 15822
rect 50428 15876 50484 16604
rect 50764 16098 50820 16110
rect 50764 16046 50766 16098
rect 50818 16046 50820 16098
rect 50764 15988 50820 16046
rect 50764 15922 50820 15932
rect 50428 15810 50484 15820
rect 50316 15698 50372 15708
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 50092 15484 50372 15540
rect 50204 15202 50260 15214
rect 50204 15150 50206 15202
rect 50258 15150 50260 15202
rect 50204 13748 50260 15150
rect 50316 15092 50372 15484
rect 50428 15428 50484 15438
rect 50876 15428 50932 17388
rect 50428 15314 50484 15372
rect 50428 15262 50430 15314
rect 50482 15262 50484 15314
rect 50428 15250 50484 15262
rect 50764 15372 50932 15428
rect 50316 15026 50372 15036
rect 50316 14644 50372 14654
rect 50316 14550 50372 14588
rect 50652 14308 50708 14346
rect 50764 14308 50820 15372
rect 50876 15204 50932 15242
rect 50876 15138 50932 15148
rect 50988 14532 51044 17724
rect 50988 14466 51044 14476
rect 51100 14642 51156 17836
rect 51324 17890 51380 17902
rect 51324 17838 51326 17890
rect 51378 17838 51380 17890
rect 51324 17442 51380 17838
rect 51324 17390 51326 17442
rect 51378 17390 51380 17442
rect 51324 16772 51380 17390
rect 51548 16996 51604 17006
rect 51548 16902 51604 16940
rect 51324 16716 51604 16772
rect 51212 16100 51268 16138
rect 51212 16034 51268 16044
rect 51100 14590 51102 14642
rect 51154 14590 51156 14642
rect 50764 14252 51044 14308
rect 50652 14242 50708 14252
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50540 13748 50596 13758
rect 49980 13746 50148 13748
rect 49980 13694 49982 13746
rect 50034 13694 50148 13746
rect 49980 13692 50148 13694
rect 50204 13746 50596 13748
rect 50204 13694 50542 13746
rect 50594 13694 50596 13746
rect 50204 13692 50596 13694
rect 49980 13682 50036 13692
rect 49868 13570 49924 13580
rect 49756 13356 50036 13412
rect 49532 13074 49700 13076
rect 49532 13022 49534 13074
rect 49586 13022 49700 13074
rect 49532 13020 49700 13022
rect 49532 13010 49588 13020
rect 49196 12962 49252 12974
rect 49196 12910 49198 12962
rect 49250 12910 49252 12962
rect 49196 12852 49252 12910
rect 49196 12786 49252 12796
rect 49644 12852 49700 12862
rect 49644 12758 49700 12796
rect 49420 12738 49476 12750
rect 49420 12686 49422 12738
rect 49474 12686 49476 12738
rect 49420 11956 49476 12686
rect 49756 12628 49812 12638
rect 49644 12516 49700 12526
rect 49644 12178 49700 12460
rect 49644 12126 49646 12178
rect 49698 12126 49700 12178
rect 49644 12114 49700 12126
rect 49420 11890 49476 11900
rect 49420 11508 49476 11518
rect 49420 11414 49476 11452
rect 49084 11228 49476 11284
rect 48860 11190 48916 11228
rect 49420 10834 49476 11228
rect 49420 10782 49422 10834
rect 49474 10782 49476 10834
rect 49420 10770 49476 10782
rect 49756 10836 49812 12572
rect 49868 12292 49924 12302
rect 49868 12198 49924 12236
rect 49868 11620 49924 11630
rect 49868 11506 49924 11564
rect 49868 11454 49870 11506
rect 49922 11454 49924 11506
rect 49868 11442 49924 11454
rect 49868 10836 49924 10846
rect 49756 10834 49924 10836
rect 49756 10782 49870 10834
rect 49922 10782 49924 10834
rect 49756 10780 49924 10782
rect 48300 9940 48356 9950
rect 48300 9714 48356 9884
rect 48300 9662 48302 9714
rect 48354 9662 48356 9714
rect 48300 9650 48356 9662
rect 48300 9268 48356 9278
rect 48300 9174 48356 9212
rect 48636 9266 48692 10108
rect 49084 10052 49140 10062
rect 49084 9958 49140 9996
rect 49532 10052 49588 10062
rect 49420 9940 49476 9950
rect 49420 9846 49476 9884
rect 48636 9214 48638 9266
rect 48690 9214 48692 9266
rect 48636 9202 48692 9214
rect 49532 9266 49588 9996
rect 49532 9214 49534 9266
rect 49586 9214 49588 9266
rect 49532 9202 49588 9214
rect 49868 9268 49924 10780
rect 49980 10612 50036 13356
rect 50092 11732 50148 13692
rect 50540 13682 50596 13692
rect 50092 11666 50148 11676
rect 50204 13524 50260 13534
rect 50204 12068 50260 13468
rect 50428 13412 50484 13422
rect 50316 12738 50372 12750
rect 50316 12686 50318 12738
rect 50370 12686 50372 12738
rect 50316 12516 50372 12686
rect 50316 12450 50372 12460
rect 50428 12740 50484 13356
rect 50652 12740 50708 12750
rect 50428 12738 50708 12740
rect 50428 12686 50654 12738
rect 50706 12686 50708 12738
rect 50428 12684 50708 12686
rect 50316 12068 50372 12078
rect 50204 12066 50372 12068
rect 50204 12014 50318 12066
rect 50370 12014 50372 12066
rect 50204 12012 50372 12014
rect 50204 11396 50260 12012
rect 50316 12002 50372 12012
rect 50428 11956 50484 12684
rect 50652 12674 50708 12684
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 50876 12404 50932 12414
rect 50876 12310 50932 12348
rect 50540 11956 50596 11966
rect 50428 11900 50540 11956
rect 50540 11732 50596 11900
rect 50764 11844 50820 11854
rect 50764 11732 50932 11788
rect 50540 11666 50596 11676
rect 49980 10546 50036 10556
rect 50092 11340 50260 11396
rect 50652 11620 50708 11630
rect 49980 9268 50036 9278
rect 49868 9266 50036 9268
rect 49868 9214 49982 9266
rect 50034 9214 50036 9266
rect 49868 9212 50036 9214
rect 48188 8988 48580 9044
rect 48300 8034 48356 8046
rect 48300 7982 48302 8034
rect 48354 7982 48356 8034
rect 47852 7700 47908 7710
rect 47740 7698 47908 7700
rect 47740 7646 47854 7698
rect 47906 7646 47908 7698
rect 47740 7644 47908 7646
rect 47852 7634 47908 7644
rect 47628 6066 47684 6076
rect 48188 6916 48244 6926
rect 48188 6130 48244 6860
rect 48188 6078 48190 6130
rect 48242 6078 48244 6130
rect 47292 5794 47348 5806
rect 47292 5742 47294 5794
rect 47346 5742 47348 5794
rect 47292 5348 47348 5742
rect 48188 5796 48244 6078
rect 48188 5730 48244 5740
rect 48300 6578 48356 7982
rect 48300 6526 48302 6578
rect 48354 6526 48356 6578
rect 48300 5572 48356 6526
rect 48524 7698 48580 8988
rect 48524 7646 48526 7698
rect 48578 7646 48580 7698
rect 48524 6580 48580 7646
rect 49084 8034 49140 8046
rect 49084 7982 49086 8034
rect 49138 7982 49140 8034
rect 49084 6692 49140 7982
rect 49420 8036 49476 8046
rect 49420 7252 49476 7980
rect 49532 7700 49588 7710
rect 49532 7606 49588 7644
rect 49868 7698 49924 9212
rect 49980 9202 50036 9212
rect 49980 8260 50036 8270
rect 49980 8166 50036 8204
rect 49868 7646 49870 7698
rect 49922 7646 49924 7698
rect 49868 7364 49924 7646
rect 50092 7588 50148 11340
rect 50316 11284 50372 11294
rect 50204 11172 50260 11182
rect 50204 11078 50260 11116
rect 50092 7522 50148 7532
rect 50204 10724 50260 10734
rect 49868 7298 49924 7308
rect 49420 7186 49476 7196
rect 50204 6692 50260 10668
rect 50316 10164 50372 11228
rect 50652 11172 50708 11564
rect 50652 11106 50708 11116
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50764 10836 50820 10846
rect 50876 10836 50932 11732
rect 50988 11508 51044 14252
rect 50988 11442 51044 11452
rect 51100 13524 51156 14590
rect 50764 10834 50932 10836
rect 50764 10782 50766 10834
rect 50818 10782 50932 10834
rect 50764 10780 50932 10782
rect 50988 10948 51044 10958
rect 50764 10770 50820 10780
rect 50428 10498 50484 10510
rect 50428 10446 50430 10498
rect 50482 10446 50484 10498
rect 50428 10386 50484 10446
rect 50428 10334 50430 10386
rect 50482 10334 50484 10386
rect 50428 10322 50484 10334
rect 50876 10164 50932 10174
rect 50316 10108 50484 10164
rect 50428 9156 50484 10108
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 50316 9100 50484 9156
rect 50316 8036 50372 9100
rect 50428 8932 50484 8942
rect 50428 8838 50484 8876
rect 50876 8708 50932 10108
rect 50428 8652 50932 8708
rect 50428 8370 50484 8652
rect 50428 8318 50430 8370
rect 50482 8318 50484 8370
rect 50428 8306 50484 8318
rect 50876 8484 50932 8494
rect 50876 8370 50932 8428
rect 50876 8318 50878 8370
rect 50930 8318 50932 8370
rect 50876 8306 50932 8318
rect 50316 7980 50484 8036
rect 50316 7700 50372 7710
rect 50316 7606 50372 7644
rect 50316 6692 50372 6702
rect 50204 6690 50372 6692
rect 50204 6638 50318 6690
rect 50370 6638 50372 6690
rect 50204 6636 50372 6638
rect 49084 6626 49140 6636
rect 48524 6514 48580 6524
rect 49420 6580 49476 6590
rect 49420 6486 49476 6524
rect 49868 6580 49924 6590
rect 49084 6466 49140 6478
rect 49084 6414 49086 6466
rect 49138 6414 49140 6466
rect 48524 6132 48580 6142
rect 48524 6038 48580 6076
rect 48972 6132 49028 6142
rect 47292 5282 47348 5292
rect 48076 5516 48356 5572
rect 47740 4900 47796 4910
rect 47068 3614 47070 3666
rect 47122 3614 47124 3666
rect 47068 3602 47124 3614
rect 47516 4788 47572 4798
rect 47516 3666 47572 4732
rect 47740 4564 47796 4844
rect 48076 4564 48132 5516
rect 48972 5348 49028 6076
rect 49084 5684 49140 6414
rect 49868 6132 49924 6524
rect 49868 6066 49924 6076
rect 49980 6020 50036 6030
rect 49420 5908 49476 5918
rect 49084 5618 49140 5628
rect 49308 5906 49476 5908
rect 49308 5854 49422 5906
rect 49474 5854 49476 5906
rect 49308 5852 49476 5854
rect 49084 5348 49140 5358
rect 48972 5346 49140 5348
rect 48972 5294 49086 5346
rect 49138 5294 49140 5346
rect 48972 5292 49140 5294
rect 49084 5282 49140 5292
rect 47740 4562 48020 4564
rect 47740 4510 47742 4562
rect 47794 4510 48020 4562
rect 47740 4508 48020 4510
rect 47740 4498 47796 4508
rect 47516 3614 47518 3666
rect 47570 3614 47572 3666
rect 47516 3602 47572 3614
rect 47964 3668 48020 4508
rect 48076 4432 48132 4508
rect 48524 4900 48580 4910
rect 48524 3892 48580 4844
rect 48524 3826 48580 3836
rect 48748 4226 48804 4238
rect 48748 4174 48750 4226
rect 48802 4174 48804 4226
rect 48748 3780 48804 4174
rect 48748 3714 48804 3724
rect 48076 3668 48132 3678
rect 47964 3666 48132 3668
rect 47964 3614 48078 3666
rect 48130 3614 48132 3666
rect 47964 3612 48132 3614
rect 48076 3556 48132 3612
rect 48860 3668 48916 3678
rect 48860 3574 48916 3612
rect 49308 3668 49364 5852
rect 49420 5842 49476 5852
rect 49980 5906 50036 5964
rect 49980 5854 49982 5906
rect 50034 5854 50036 5906
rect 49868 5460 49924 5470
rect 49868 5234 49924 5404
rect 49868 5182 49870 5234
rect 49922 5182 49924 5234
rect 49868 5170 49924 5182
rect 49980 5236 50036 5854
rect 49980 5170 50036 5180
rect 50316 5234 50372 6636
rect 50316 5182 50318 5234
rect 50370 5182 50372 5234
rect 50316 5170 50372 5182
rect 49644 4676 49700 4686
rect 49420 4114 49476 4126
rect 49420 4062 49422 4114
rect 49474 4062 49476 4114
rect 49420 3780 49476 4062
rect 49420 3714 49476 3724
rect 49644 3780 49700 4620
rect 49980 4564 50036 4574
rect 49980 4470 50036 4508
rect 49644 3714 49700 3724
rect 49756 4004 49812 4014
rect 49308 3574 49364 3612
rect 48076 3490 48132 3500
rect 49756 3556 49812 3948
rect 50428 3892 50484 7980
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 50876 7476 50932 7486
rect 50764 7364 50820 7374
rect 50764 6690 50820 7308
rect 50876 7362 50932 7420
rect 50876 7310 50878 7362
rect 50930 7310 50932 7362
rect 50876 6804 50932 7310
rect 50876 6738 50932 6748
rect 50764 6638 50766 6690
rect 50818 6638 50820 6690
rect 50764 6626 50820 6638
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 50764 5346 50820 5358
rect 50764 5294 50766 5346
rect 50818 5294 50820 5346
rect 50764 5234 50820 5294
rect 50764 5182 50766 5234
rect 50818 5182 50820 5234
rect 50764 5170 50820 5182
rect 50988 5236 51044 10892
rect 51100 9940 51156 13468
rect 51212 15876 51268 15886
rect 51212 12292 51268 15820
rect 51324 15764 51380 15774
rect 51324 15538 51380 15708
rect 51324 15486 51326 15538
rect 51378 15486 51380 15538
rect 51324 15474 51380 15486
rect 51324 14418 51380 14430
rect 51324 14366 51326 14418
rect 51378 14366 51380 14418
rect 51324 13970 51380 14366
rect 51324 13918 51326 13970
rect 51378 13918 51380 13970
rect 51324 13906 51380 13918
rect 51436 12852 51492 12862
rect 51436 12758 51492 12796
rect 51548 12404 51604 16716
rect 51660 14418 51716 18396
rect 51772 18340 51828 19292
rect 51996 19012 52052 21756
rect 52220 21586 52276 21598
rect 52220 21534 52222 21586
rect 52274 21534 52276 21586
rect 52220 20580 52276 21534
rect 52220 20514 52276 20524
rect 52332 20578 52388 20590
rect 52332 20526 52334 20578
rect 52386 20526 52388 20578
rect 52332 20356 52388 20526
rect 52332 20290 52388 20300
rect 51996 18946 52052 18956
rect 52108 19908 52164 19918
rect 52108 19122 52164 19852
rect 52108 19070 52110 19122
rect 52162 19070 52164 19122
rect 51884 18564 51940 18574
rect 51884 18470 51940 18508
rect 51772 18274 51828 18284
rect 51884 18004 51940 18014
rect 51772 17442 51828 17454
rect 51772 17390 51774 17442
rect 51826 17390 51828 17442
rect 51772 17108 51828 17390
rect 51772 17042 51828 17052
rect 51884 17108 51940 17948
rect 51996 17108 52052 17118
rect 51884 17106 52052 17108
rect 51884 17054 51998 17106
rect 52050 17054 52052 17106
rect 51884 17052 52052 17054
rect 51884 15764 51940 17052
rect 51996 17042 52052 17052
rect 52108 16098 52164 19070
rect 52220 19234 52276 19246
rect 52220 19182 52222 19234
rect 52274 19182 52276 19234
rect 52220 19124 52276 19182
rect 52220 19058 52276 19068
rect 52444 18900 52500 22204
rect 52108 16046 52110 16098
rect 52162 16046 52164 16098
rect 52108 16034 52164 16046
rect 52220 18844 52500 18900
rect 52220 16212 52276 18844
rect 52444 18564 52500 18574
rect 52444 18470 52500 18508
rect 52332 17780 52388 17790
rect 52332 17686 52388 17724
rect 51884 15698 51940 15708
rect 52220 15764 52276 16156
rect 52556 15988 52612 23436
rect 52668 23380 52724 29260
rect 52780 28308 52836 30604
rect 53228 29876 53284 37324
rect 53452 36370 53508 38612
rect 53564 37380 53620 37390
rect 53564 37286 53620 37324
rect 53452 36318 53454 36370
rect 53506 36318 53508 36370
rect 53452 35476 53508 36318
rect 53452 35410 53508 35420
rect 53676 36372 53732 38612
rect 53788 37826 53844 37838
rect 53788 37774 53790 37826
rect 53842 37774 53844 37826
rect 53788 37716 53844 37774
rect 53788 37650 53844 37660
rect 53900 37380 53956 39900
rect 54012 38276 54068 41804
rect 54124 41858 54180 41870
rect 54124 41806 54126 41858
rect 54178 41806 54180 41858
rect 54124 41746 54180 41806
rect 54124 41694 54126 41746
rect 54178 41694 54180 41746
rect 54124 41682 54180 41694
rect 54124 41412 54180 41422
rect 54124 41186 54180 41356
rect 54124 41134 54126 41186
rect 54178 41134 54180 41186
rect 54124 40402 54180 41134
rect 54124 40350 54126 40402
rect 54178 40350 54180 40402
rect 54124 40338 54180 40350
rect 54236 40292 54292 42588
rect 54348 41188 54404 42700
rect 54572 42690 54628 42700
rect 54572 41858 54628 41870
rect 54572 41806 54574 41858
rect 54626 41806 54628 41858
rect 54572 41636 54628 41806
rect 54348 41132 54516 41188
rect 54348 40964 54404 40974
rect 54348 40626 54404 40908
rect 54348 40574 54350 40626
rect 54402 40574 54404 40626
rect 54348 40562 54404 40574
rect 54236 40236 54404 40292
rect 54236 39732 54292 39742
rect 54124 39060 54180 39070
rect 54124 38834 54180 39004
rect 54124 38782 54126 38834
rect 54178 38782 54180 38834
rect 54124 38770 54180 38782
rect 54236 38668 54292 39676
rect 54348 38946 54404 40236
rect 54460 39508 54516 41132
rect 54460 39060 54516 39452
rect 54460 38994 54516 39004
rect 54572 39058 54628 41580
rect 54908 40180 54964 44380
rect 55020 44994 55076 45006
rect 55020 44942 55022 44994
rect 55074 44942 55076 44994
rect 55020 43540 55076 44942
rect 55020 43474 55076 43484
rect 55132 44210 55188 44222
rect 55132 44158 55134 44210
rect 55186 44158 55188 44210
rect 55020 42756 55076 42766
rect 55132 42756 55188 44158
rect 55356 43652 55412 45612
rect 55356 43586 55412 43596
rect 55468 44434 55524 46732
rect 55580 48130 55636 48142
rect 55580 48078 55582 48130
rect 55634 48078 55636 48130
rect 55580 45892 55636 48078
rect 56028 48132 56084 48142
rect 56028 48038 56084 48076
rect 56476 48130 56532 48142
rect 56476 48078 56478 48130
rect 56530 48078 56532 48130
rect 56476 47684 56532 48078
rect 56476 47618 56532 47628
rect 55692 47236 55748 47246
rect 55692 47142 55748 47180
rect 56140 47236 56196 47246
rect 56140 47234 56308 47236
rect 56140 47182 56142 47234
rect 56194 47182 56308 47234
rect 56140 47180 56308 47182
rect 56140 47170 56196 47180
rect 56028 47124 56084 47134
rect 55692 46900 55748 46910
rect 56028 46900 56084 47068
rect 56252 47012 56308 47180
rect 56252 46946 56308 46956
rect 56588 47234 56644 47246
rect 56588 47182 56590 47234
rect 56642 47182 56644 47234
rect 56140 46900 56196 46910
rect 56028 46898 56196 46900
rect 56028 46846 56142 46898
rect 56194 46846 56196 46898
rect 56028 46844 56196 46846
rect 55692 46806 55748 46844
rect 56140 46834 56196 46844
rect 56588 46788 56644 47182
rect 56588 46722 56644 46732
rect 56812 47124 56868 47134
rect 56588 46564 56644 46574
rect 56588 46470 56644 46508
rect 55580 45826 55636 45836
rect 55804 45668 55860 45678
rect 56252 45668 56308 45678
rect 56588 45668 56644 45678
rect 55804 45574 55860 45612
rect 56028 45666 56308 45668
rect 56028 45614 56254 45666
rect 56306 45614 56308 45666
rect 56028 45612 56308 45614
rect 55580 44994 55636 45006
rect 55580 44942 55582 44994
rect 55634 44942 55636 44994
rect 55580 44884 55636 44942
rect 55580 44818 55636 44828
rect 55916 44994 55972 45006
rect 55916 44942 55918 44994
rect 55970 44942 55972 44994
rect 55468 44382 55470 44434
rect 55522 44382 55524 44434
rect 55356 43426 55412 43438
rect 55356 43374 55358 43426
rect 55410 43374 55412 43426
rect 55356 43092 55412 43374
rect 55468 43316 55524 44382
rect 55916 44436 55972 44942
rect 55916 44370 55972 44380
rect 55580 44324 55636 44334
rect 55580 44230 55636 44268
rect 55468 43250 55524 43260
rect 55356 43026 55412 43036
rect 55020 42754 55132 42756
rect 55020 42702 55022 42754
rect 55074 42702 55132 42754
rect 55020 42700 55132 42702
rect 55020 42690 55076 42700
rect 55132 42690 55188 42700
rect 55356 42812 55972 42868
rect 55132 42530 55188 42542
rect 55132 42478 55134 42530
rect 55186 42478 55188 42530
rect 55020 41746 55076 41758
rect 55020 41694 55022 41746
rect 55074 41694 55076 41746
rect 55020 40740 55076 41694
rect 55132 41188 55188 42478
rect 55244 42532 55300 42542
rect 55356 42532 55412 42812
rect 55916 42754 55972 42812
rect 55916 42702 55918 42754
rect 55970 42702 55972 42754
rect 55916 42690 55972 42702
rect 55244 42530 55412 42532
rect 55244 42478 55246 42530
rect 55298 42478 55412 42530
rect 55244 42476 55412 42478
rect 55244 42466 55300 42476
rect 55356 42084 55412 42476
rect 55804 42642 55860 42654
rect 55804 42590 55806 42642
rect 55858 42590 55860 42642
rect 55468 42084 55524 42094
rect 55356 42082 55524 42084
rect 55356 42030 55470 42082
rect 55522 42030 55524 42082
rect 55356 42028 55524 42030
rect 55132 41122 55188 41132
rect 55244 41972 55300 41982
rect 55244 41186 55300 41916
rect 55244 41134 55246 41186
rect 55298 41134 55300 41186
rect 55244 41076 55300 41134
rect 55244 41010 55300 41020
rect 55356 40962 55412 40974
rect 55356 40910 55358 40962
rect 55410 40910 55412 40962
rect 55020 40684 55300 40740
rect 55132 40516 55188 40526
rect 55132 40422 55188 40460
rect 55020 40404 55076 40414
rect 55020 40310 55076 40348
rect 55244 40180 55300 40684
rect 55356 40404 55412 40910
rect 55468 40964 55524 42028
rect 55580 42084 55636 42094
rect 55580 41858 55636 42028
rect 55580 41806 55582 41858
rect 55634 41806 55636 41858
rect 55580 41794 55636 41806
rect 55468 40898 55524 40908
rect 55580 41636 55636 41646
rect 55356 40338 55412 40348
rect 55468 40740 55524 40750
rect 54908 40124 55188 40180
rect 55244 40124 55412 40180
rect 54908 39508 54964 39518
rect 54908 39414 54964 39452
rect 54572 39006 54574 39058
rect 54626 39006 54628 39058
rect 54572 38994 54628 39006
rect 55020 39394 55076 39406
rect 55020 39342 55022 39394
rect 55074 39342 55076 39394
rect 55020 39060 55076 39342
rect 55020 38994 55076 39004
rect 54348 38894 54350 38946
rect 54402 38894 54404 38946
rect 54348 38882 54404 38894
rect 54012 38210 54068 38220
rect 54124 38612 54292 38668
rect 54908 38724 54964 38762
rect 54908 38658 54964 38668
rect 55132 38668 55188 40124
rect 55244 39620 55300 39630
rect 55244 39526 55300 39564
rect 55244 38948 55300 38958
rect 55244 38854 55300 38892
rect 53676 35140 53732 36316
rect 53788 37324 53956 37380
rect 53788 36258 53844 37324
rect 54124 36820 54180 38612
rect 55020 38610 55076 38622
rect 55132 38612 55300 38668
rect 55020 38558 55022 38610
rect 55074 38558 55076 38610
rect 55020 38500 55076 38558
rect 55020 38444 55188 38500
rect 53900 36484 53956 36494
rect 53900 36390 53956 36428
rect 53788 36206 53790 36258
rect 53842 36206 53844 36258
rect 53788 36194 53844 36206
rect 54012 35924 54068 35934
rect 54012 35810 54068 35868
rect 54012 35758 54014 35810
rect 54066 35758 54068 35810
rect 54012 35746 54068 35758
rect 53340 35084 53732 35140
rect 53340 33348 53396 35084
rect 53788 34916 53844 34926
rect 53788 34822 53844 34860
rect 53452 34802 53508 34814
rect 53452 34750 53454 34802
rect 53506 34750 53508 34802
rect 53452 34244 53508 34750
rect 53564 34804 53620 34814
rect 53564 34710 53620 34748
rect 54124 34692 54180 36764
rect 54684 38276 54740 38286
rect 54348 36708 54404 36718
rect 54236 36706 54404 36708
rect 54236 36654 54350 36706
rect 54402 36654 54404 36706
rect 54236 36652 54404 36654
rect 54236 36482 54292 36652
rect 54348 36642 54404 36652
rect 54236 36430 54238 36482
rect 54290 36430 54292 36482
rect 54236 36418 54292 36430
rect 54460 34916 54516 34926
rect 54684 34916 54740 38220
rect 54908 38052 54964 38062
rect 54908 37958 54964 37996
rect 55020 37940 55076 37950
rect 55020 37846 55076 37884
rect 54796 37828 54852 37838
rect 54796 37734 54852 37772
rect 55132 36484 55188 38444
rect 55244 36706 55300 38612
rect 55244 36654 55246 36706
rect 55298 36654 55300 36706
rect 55244 36642 55300 36654
rect 55020 36428 55188 36484
rect 54796 36258 54852 36270
rect 54796 36206 54798 36258
rect 54850 36206 54852 36258
rect 54796 35364 54852 36206
rect 54796 35298 54852 35308
rect 54684 34860 54852 34916
rect 54460 34822 54516 34860
rect 53788 34636 54180 34692
rect 54684 34692 54740 34702
rect 53676 34244 53732 34254
rect 53452 34242 53732 34244
rect 53452 34190 53678 34242
rect 53730 34190 53732 34242
rect 53452 34188 53732 34190
rect 53564 33572 53620 34188
rect 53676 34178 53732 34188
rect 53788 34130 53844 34636
rect 53788 34078 53790 34130
rect 53842 34078 53844 34130
rect 53676 33906 53732 33918
rect 53676 33854 53678 33906
rect 53730 33854 53732 33906
rect 53676 33796 53732 33854
rect 53676 33730 53732 33740
rect 53564 33506 53620 33516
rect 53340 33292 53620 33348
rect 53340 33124 53396 33134
rect 53340 33030 53396 33068
rect 53452 32788 53508 32798
rect 53452 32674 53508 32732
rect 53452 32622 53454 32674
rect 53506 32622 53508 32674
rect 53452 32610 53508 32622
rect 53340 32004 53396 32014
rect 53340 30212 53396 31948
rect 53452 31666 53508 31678
rect 53452 31614 53454 31666
rect 53506 31614 53508 31666
rect 53452 31556 53508 31614
rect 53452 31490 53508 31500
rect 53564 30772 53620 33292
rect 53788 33124 53844 34078
rect 53900 34468 53956 34478
rect 53900 33346 53956 34412
rect 54684 34356 54740 34636
rect 54460 34300 54740 34356
rect 54348 33906 54404 33918
rect 54348 33854 54350 33906
rect 54402 33854 54404 33906
rect 54348 33460 54404 33854
rect 54348 33366 54404 33404
rect 53900 33294 53902 33346
rect 53954 33294 53956 33346
rect 53900 33282 53956 33294
rect 54012 33348 54068 33358
rect 53788 33068 53956 33124
rect 53676 32562 53732 32574
rect 53676 32510 53678 32562
rect 53730 32510 53732 32562
rect 53676 32452 53732 32510
rect 53676 32386 53732 32396
rect 53788 32450 53844 32462
rect 53788 32398 53790 32450
rect 53842 32398 53844 32450
rect 53676 32004 53732 32014
rect 53676 31890 53732 31948
rect 53676 31838 53678 31890
rect 53730 31838 53732 31890
rect 53676 31826 53732 31838
rect 53676 31668 53732 31678
rect 53676 31574 53732 31612
rect 53676 30996 53732 31006
rect 53788 30996 53844 32398
rect 53900 31780 53956 33068
rect 54012 32562 54068 33292
rect 54012 32510 54014 32562
rect 54066 32510 54068 32562
rect 54012 32116 54068 32510
rect 54012 32050 54068 32060
rect 54236 33346 54292 33358
rect 54236 33294 54238 33346
rect 54290 33294 54292 33346
rect 54236 32338 54292 33294
rect 54236 32286 54238 32338
rect 54290 32286 54292 32338
rect 53900 31714 53956 31724
rect 54236 31778 54292 32286
rect 54236 31726 54238 31778
rect 54290 31726 54292 31778
rect 54236 31714 54292 31726
rect 53676 30994 53844 30996
rect 53676 30942 53678 30994
rect 53730 30942 53844 30994
rect 53676 30940 53844 30942
rect 53676 30930 53732 30940
rect 54124 30884 54180 30894
rect 53564 30716 53732 30772
rect 53340 30156 53620 30212
rect 52780 28242 52836 28252
rect 53004 29820 53284 29876
rect 53340 29988 53396 29998
rect 53004 28082 53060 29820
rect 53228 29426 53284 29438
rect 53228 29374 53230 29426
rect 53282 29374 53284 29426
rect 53228 28868 53284 29374
rect 53228 28802 53284 28812
rect 53004 28030 53006 28082
rect 53058 28030 53060 28082
rect 53004 28018 53060 28030
rect 53116 28308 53172 28318
rect 53116 27970 53172 28252
rect 53116 27918 53118 27970
rect 53170 27918 53172 27970
rect 53004 27858 53060 27870
rect 53004 27806 53006 27858
rect 53058 27806 53060 27858
rect 53004 27300 53060 27806
rect 53116 27860 53172 27918
rect 53116 27794 53172 27804
rect 53004 27234 53060 27244
rect 53340 26908 53396 29932
rect 53564 29538 53620 30156
rect 53564 29486 53566 29538
rect 53618 29486 53620 29538
rect 53564 29316 53620 29486
rect 53564 29250 53620 29260
rect 53676 28754 53732 30716
rect 53788 30324 53844 30334
rect 53788 30210 53844 30268
rect 53788 30158 53790 30210
rect 53842 30158 53844 30210
rect 53788 30146 53844 30158
rect 54124 29652 54180 30828
rect 54236 30548 54292 30558
rect 54236 30212 54292 30492
rect 54236 30210 54404 30212
rect 54236 30158 54238 30210
rect 54290 30158 54404 30210
rect 54236 30156 54404 30158
rect 54236 30146 54292 30156
rect 54236 29652 54292 29662
rect 54124 29650 54292 29652
rect 54124 29598 54238 29650
rect 54290 29598 54292 29650
rect 54124 29596 54292 29598
rect 54236 29586 54292 29596
rect 53676 28702 53678 28754
rect 53730 28702 53732 28754
rect 53676 28690 53732 28702
rect 54012 28644 54068 28654
rect 54012 28642 54180 28644
rect 54012 28590 54014 28642
rect 54066 28590 54180 28642
rect 54012 28588 54180 28590
rect 54012 28578 54068 28588
rect 53564 28420 53620 28430
rect 53564 28326 53620 28364
rect 53788 28418 53844 28430
rect 53788 28366 53790 28418
rect 53842 28366 53844 28418
rect 53564 27300 53620 27310
rect 53564 27206 53620 27244
rect 53676 27074 53732 27086
rect 53676 27022 53678 27074
rect 53730 27022 53732 27074
rect 53340 26852 53620 26908
rect 52780 26516 52836 26526
rect 52780 26514 53172 26516
rect 52780 26462 52782 26514
rect 52834 26462 53172 26514
rect 52780 26460 53172 26462
rect 52780 26450 52836 26460
rect 52892 26290 52948 26302
rect 52892 26238 52894 26290
rect 52946 26238 52948 26290
rect 52780 26068 52836 26078
rect 52780 25974 52836 26012
rect 52892 25956 52948 26238
rect 52892 25890 52948 25900
rect 53004 25732 53060 25742
rect 52780 24722 52836 24734
rect 52780 24670 52782 24722
rect 52834 24670 52836 24722
rect 52780 23940 52836 24670
rect 52780 23874 52836 23884
rect 53004 24722 53060 25676
rect 53004 24670 53006 24722
rect 53058 24670 53060 24722
rect 52668 23324 52948 23380
rect 52780 23154 52836 23166
rect 52780 23102 52782 23154
rect 52834 23102 52836 23154
rect 52780 22260 52836 23102
rect 52780 22194 52836 22204
rect 52668 21476 52724 21486
rect 52668 20916 52724 21420
rect 52892 21364 52948 23324
rect 52892 21298 52948 21308
rect 52668 20850 52724 20860
rect 53004 20580 53060 24670
rect 53004 20130 53060 20524
rect 53116 20188 53172 26460
rect 53228 26404 53284 26414
rect 53228 25396 53284 26348
rect 53340 26180 53396 26190
rect 53452 26180 53508 26190
rect 53396 26178 53508 26180
rect 53396 26126 53454 26178
rect 53506 26126 53508 26178
rect 53396 26124 53508 26126
rect 53340 25620 53396 26124
rect 53452 26114 53508 26124
rect 53340 25554 53396 25564
rect 53452 25508 53508 25518
rect 53228 25340 53396 25396
rect 53228 23044 53284 23054
rect 53228 22950 53284 22988
rect 53340 22820 53396 25340
rect 53452 24946 53508 25452
rect 53564 25060 53620 26852
rect 53676 26852 53732 27022
rect 53676 26786 53732 26796
rect 53788 26628 53844 28366
rect 53676 26572 53844 26628
rect 53900 27860 53956 27870
rect 53676 25732 53732 26572
rect 53900 26516 53956 27804
rect 54124 27076 54180 28588
rect 54236 28642 54292 28654
rect 54236 28590 54238 28642
rect 54290 28590 54292 28642
rect 54236 27972 54292 28590
rect 54236 27906 54292 27916
rect 54348 27636 54404 30156
rect 54460 28308 54516 34300
rect 54684 34132 54740 34142
rect 54684 34038 54740 34076
rect 54572 33346 54628 33358
rect 54572 33294 54574 33346
rect 54626 33294 54628 33346
rect 54572 33236 54628 33294
rect 54572 32116 54628 33180
rect 54796 32340 54852 34860
rect 54908 34018 54964 34030
rect 54908 33966 54910 34018
rect 54962 33966 54964 34018
rect 54908 33908 54964 33966
rect 54908 33842 54964 33852
rect 55020 32562 55076 36428
rect 55132 36260 55188 36270
rect 55132 36166 55188 36204
rect 55356 35140 55412 40124
rect 55468 36484 55524 40684
rect 55580 38668 55636 41580
rect 55804 40628 55860 42590
rect 56028 40740 56084 45612
rect 56252 45602 56308 45612
rect 56476 45666 56644 45668
rect 56476 45614 56590 45666
rect 56642 45614 56644 45666
rect 56476 45612 56644 45614
rect 56364 44996 56420 45006
rect 56364 44902 56420 44940
rect 56140 44100 56196 44110
rect 56140 43538 56196 44044
rect 56140 43486 56142 43538
rect 56194 43486 56196 43538
rect 56140 43474 56196 43486
rect 56364 43316 56420 43326
rect 56252 42756 56308 42766
rect 56252 42662 56308 42700
rect 56364 42194 56420 43260
rect 56364 42142 56366 42194
rect 56418 42142 56420 42194
rect 56364 42130 56420 42142
rect 56140 42084 56196 42094
rect 56140 41990 56196 42028
rect 56252 41860 56308 41870
rect 56252 41858 56420 41860
rect 56252 41806 56254 41858
rect 56306 41806 56420 41858
rect 56252 41804 56420 41806
rect 56252 41794 56308 41804
rect 56028 40674 56084 40684
rect 56140 41188 56196 41198
rect 56364 41188 56420 41804
rect 56476 41636 56532 45612
rect 56588 45602 56644 45612
rect 56588 44098 56644 44110
rect 56588 44046 56590 44098
rect 56642 44046 56644 44098
rect 56588 43764 56644 44046
rect 56588 43698 56644 43708
rect 56588 43428 56644 43438
rect 56588 43334 56644 43372
rect 56700 41972 56756 41982
rect 56476 41570 56532 41580
rect 56588 41970 56756 41972
rect 56588 41918 56702 41970
rect 56754 41918 56756 41970
rect 56588 41916 56756 41918
rect 56364 41132 56532 41188
rect 55804 40572 55972 40628
rect 55692 40516 55748 40526
rect 55692 39618 55748 40460
rect 55804 40404 55860 40414
rect 55804 40310 55860 40348
rect 55916 39956 55972 40572
rect 56140 40402 56196 41132
rect 56252 41076 56308 41086
rect 56252 40982 56308 41020
rect 56364 40964 56420 40974
rect 56364 40870 56420 40908
rect 56140 40350 56142 40402
rect 56194 40350 56196 40402
rect 55916 39900 56084 39956
rect 55692 39566 55694 39618
rect 55746 39566 55748 39618
rect 55692 38948 55748 39566
rect 55916 39732 55972 39742
rect 55916 39618 55972 39676
rect 55916 39566 55918 39618
rect 55970 39566 55972 39618
rect 55916 39554 55972 39566
rect 55804 39508 55860 39518
rect 55804 39414 55860 39452
rect 55692 38882 55748 38892
rect 56028 38834 56084 39900
rect 56140 39732 56196 40350
rect 56476 40180 56532 41132
rect 56588 41186 56644 41916
rect 56700 41906 56756 41916
rect 56812 41412 56868 47068
rect 56924 43428 56980 55244
rect 57148 53844 57204 53854
rect 57036 49700 57092 49710
rect 57036 47570 57092 49644
rect 57036 47518 57038 47570
rect 57090 47518 57092 47570
rect 57036 47506 57092 47518
rect 57148 44660 57204 53788
rect 57932 50820 57988 50830
rect 57484 48132 57540 48142
rect 57484 48130 57652 48132
rect 57484 48078 57486 48130
rect 57538 48078 57652 48130
rect 57484 48076 57652 48078
rect 57484 48066 57540 48076
rect 57484 47796 57540 47806
rect 57484 47570 57540 47740
rect 57484 47518 57486 47570
rect 57538 47518 57540 47570
rect 57484 47506 57540 47518
rect 57372 46564 57428 46574
rect 57372 46470 57428 46508
rect 57260 46114 57316 46126
rect 57260 46062 57262 46114
rect 57314 46062 57316 46114
rect 57260 46002 57316 46062
rect 57260 45950 57262 46002
rect 57314 45950 57316 46002
rect 57260 45938 57316 45950
rect 57596 46004 57652 48076
rect 57932 47572 57988 50764
rect 57596 45938 57652 45948
rect 57708 47570 57988 47572
rect 57708 47518 57934 47570
rect 57986 47518 57988 47570
rect 57708 47516 57988 47518
rect 57596 45666 57652 45678
rect 57596 45614 57598 45666
rect 57650 45614 57652 45666
rect 57484 45220 57540 45230
rect 57484 45126 57540 45164
rect 57148 44594 57204 44604
rect 57596 44548 57652 45614
rect 57596 44482 57652 44492
rect 57484 44324 57540 44334
rect 57708 44324 57764 47516
rect 57932 47506 57988 47516
rect 57820 46788 57876 46798
rect 57820 46694 57876 46732
rect 58044 46114 58100 46126
rect 58044 46062 58046 46114
rect 58098 46062 58100 46114
rect 57820 46004 57876 46014
rect 57820 45218 57876 45948
rect 58044 45666 58100 46062
rect 58044 45614 58046 45666
rect 58098 45614 58100 45666
rect 58044 45556 58100 45614
rect 58828 45668 58884 45678
rect 57820 45166 57822 45218
rect 57874 45166 57876 45218
rect 57820 45154 57876 45166
rect 57932 45500 58660 45556
rect 57932 44324 57988 45500
rect 57484 44322 57764 44324
rect 57484 44270 57486 44322
rect 57538 44270 57764 44322
rect 57484 44268 57764 44270
rect 57820 44268 57988 44324
rect 58044 45220 58100 45230
rect 57484 44258 57540 44268
rect 57820 44212 57876 44268
rect 57708 44156 57876 44212
rect 57148 44100 57204 44110
rect 57148 44006 57204 44044
rect 57372 43540 57428 43550
rect 57708 43540 57764 44156
rect 57932 44100 57988 44110
rect 57372 43538 57764 43540
rect 57372 43486 57374 43538
rect 57426 43486 57764 43538
rect 57372 43484 57764 43486
rect 57820 44098 57988 44100
rect 57820 44046 57934 44098
rect 57986 44046 57988 44098
rect 57820 44044 57988 44046
rect 57372 43474 57428 43484
rect 56924 43362 56980 43372
rect 57820 43428 57876 44044
rect 57932 44034 57988 44044
rect 57820 43362 57876 43372
rect 57932 43426 57988 43438
rect 57932 43374 57934 43426
rect 57986 43374 57988 43426
rect 56812 41346 56868 41356
rect 57148 42978 57204 42990
rect 57148 42926 57150 42978
rect 57202 42926 57204 42978
rect 56588 41134 56590 41186
rect 56642 41134 56644 41186
rect 56588 41122 56644 41134
rect 57036 40962 57092 40974
rect 57036 40910 57038 40962
rect 57090 40910 57092 40962
rect 56700 40292 56756 40302
rect 56700 40290 56980 40292
rect 56700 40238 56702 40290
rect 56754 40238 56980 40290
rect 56700 40236 56980 40238
rect 56700 40226 56756 40236
rect 56476 40114 56532 40124
rect 56812 40068 56868 40078
rect 56140 39172 56196 39676
rect 56700 39844 56756 39854
rect 56364 39620 56420 39630
rect 56364 39618 56644 39620
rect 56364 39566 56366 39618
rect 56418 39566 56644 39618
rect 56364 39564 56644 39566
rect 56364 39554 56420 39564
rect 56140 39106 56196 39116
rect 56364 39396 56420 39406
rect 56028 38782 56030 38834
rect 56082 38782 56084 38834
rect 55580 38612 55748 38668
rect 55692 37492 55748 38612
rect 55804 38612 55860 38622
rect 55804 38162 55860 38556
rect 55804 38110 55806 38162
rect 55858 38110 55860 38162
rect 55804 38098 55860 38110
rect 56028 38050 56084 38782
rect 56252 38612 56308 38622
rect 56252 38518 56308 38556
rect 56028 37998 56030 38050
rect 56082 37998 56084 38050
rect 56028 37986 56084 37998
rect 56140 38274 56196 38286
rect 56140 38222 56142 38274
rect 56194 38222 56196 38274
rect 56140 37828 56196 38222
rect 55692 37436 55972 37492
rect 55804 37268 55860 37278
rect 55692 37154 55748 37166
rect 55692 37102 55694 37154
rect 55746 37102 55748 37154
rect 55692 37044 55748 37102
rect 55692 36978 55748 36988
rect 55468 36428 55748 36484
rect 55580 36258 55636 36270
rect 55580 36206 55582 36258
rect 55634 36206 55636 36258
rect 55580 35588 55636 36206
rect 55580 35522 55636 35532
rect 55244 35084 55412 35140
rect 55468 35476 55524 35486
rect 55020 32510 55022 32562
rect 55074 32510 55076 32562
rect 55020 32498 55076 32510
rect 55132 35028 55188 35038
rect 55132 34356 55188 34972
rect 54796 32284 55076 32340
rect 54572 32050 54628 32060
rect 54908 31778 54964 31790
rect 54908 31726 54910 31778
rect 54962 31726 54964 31778
rect 54908 31444 54964 31726
rect 54796 31106 54852 31118
rect 54796 31054 54798 31106
rect 54850 31054 54852 31106
rect 54796 30436 54852 31054
rect 54796 30370 54852 30380
rect 54684 30212 54740 30222
rect 54684 30118 54740 30156
rect 54684 29988 54740 29998
rect 54684 29092 54740 29932
rect 54908 29652 54964 31388
rect 54684 29026 54740 29036
rect 54796 29596 54964 29652
rect 55020 29650 55076 32284
rect 55132 30212 55188 34300
rect 55244 34132 55300 35084
rect 55356 34916 55412 34926
rect 55468 34916 55524 35420
rect 55692 35028 55748 36428
rect 55692 34962 55748 34972
rect 55412 34860 55524 34916
rect 55804 34916 55860 37212
rect 55356 34784 55412 34860
rect 55804 34850 55860 34860
rect 55580 34804 55636 34814
rect 55468 34748 55580 34804
rect 55468 34242 55524 34748
rect 55580 34738 55636 34748
rect 55692 34692 55748 34702
rect 55468 34190 55470 34242
rect 55522 34190 55524 34242
rect 55244 34076 55412 34132
rect 55244 33908 55300 33918
rect 55244 31892 55300 33852
rect 55244 31778 55300 31836
rect 55244 31726 55246 31778
rect 55298 31726 55300 31778
rect 55244 31714 55300 31726
rect 55356 31890 55412 34076
rect 55468 33796 55524 34190
rect 55580 34356 55636 34366
rect 55692 34356 55748 34636
rect 55580 34354 55748 34356
rect 55580 34302 55582 34354
rect 55634 34302 55748 34354
rect 55580 34300 55748 34302
rect 55580 34244 55636 34300
rect 55580 34178 55636 34188
rect 55468 33730 55524 33740
rect 55356 31838 55358 31890
rect 55410 31838 55412 31890
rect 55356 31220 55412 31838
rect 55356 31154 55412 31164
rect 55356 30994 55412 31006
rect 55356 30942 55358 30994
rect 55410 30942 55412 30994
rect 55356 30212 55412 30942
rect 55132 30156 55412 30212
rect 55132 29988 55188 29998
rect 55132 29894 55188 29932
rect 55020 29598 55022 29650
rect 55074 29598 55076 29650
rect 54460 28242 54516 28252
rect 54348 27570 54404 27580
rect 54460 28084 54516 28094
rect 54124 27010 54180 27020
rect 54348 27188 54404 27198
rect 54348 27074 54404 27132
rect 54348 27022 54350 27074
rect 54402 27022 54404 27074
rect 54348 27010 54404 27022
rect 54236 26964 54292 26974
rect 53676 25666 53732 25676
rect 53788 26460 53956 26516
rect 54124 26852 54292 26908
rect 54460 26964 54516 28028
rect 54684 27972 54740 27982
rect 54460 26898 54516 26908
rect 54572 27858 54628 27870
rect 54572 27806 54574 27858
rect 54626 27806 54628 27858
rect 54348 26852 54404 26862
rect 53676 25506 53732 25518
rect 53676 25454 53678 25506
rect 53730 25454 53732 25506
rect 53676 25284 53732 25454
rect 53676 25218 53732 25228
rect 53788 25394 53844 26460
rect 53788 25342 53790 25394
rect 53842 25342 53844 25394
rect 53564 25004 53732 25060
rect 53452 24894 53454 24946
rect 53506 24894 53508 24946
rect 53452 24882 53508 24894
rect 53564 24724 53620 24734
rect 53564 24630 53620 24668
rect 53452 23940 53508 23950
rect 53452 23380 53508 23884
rect 53676 23492 53732 25004
rect 53676 23426 53732 23436
rect 53788 24722 53844 25342
rect 54012 26290 54068 26302
rect 54012 26238 54014 26290
rect 54066 26238 54068 26290
rect 54012 25172 54068 26238
rect 53788 24670 53790 24722
rect 53842 24670 53844 24722
rect 53452 23314 53508 23324
rect 53228 22764 53396 22820
rect 53452 23156 53508 23166
rect 53228 21140 53284 22764
rect 53452 22258 53508 23100
rect 53788 22932 53844 24670
rect 53900 25116 54012 25172
rect 53900 23940 53956 25116
rect 54012 25106 54068 25116
rect 54124 25060 54180 26852
rect 54124 24994 54180 25004
rect 54012 24948 54068 24958
rect 54012 24854 54068 24892
rect 53900 23154 53956 23884
rect 54124 24722 54180 24734
rect 54124 24670 54126 24722
rect 54178 24670 54180 24722
rect 53900 23102 53902 23154
rect 53954 23102 53956 23154
rect 53900 23090 53956 23102
rect 54012 23826 54068 23838
rect 54012 23774 54014 23826
rect 54066 23774 54068 23826
rect 54012 22932 54068 23774
rect 53788 22876 54068 22932
rect 53452 22206 53454 22258
rect 53506 22206 53508 22258
rect 53452 21588 53508 22206
rect 53788 22148 53844 22158
rect 53788 21812 53844 22092
rect 53452 21522 53508 21532
rect 53676 21756 53844 21812
rect 53340 21476 53396 21486
rect 53340 21382 53396 21420
rect 53676 21364 53732 21756
rect 53788 21588 53844 21598
rect 53788 21494 53844 21532
rect 53676 21308 53844 21364
rect 53340 21140 53396 21150
rect 53228 21084 53340 21140
rect 53340 20914 53396 21084
rect 53340 20862 53342 20914
rect 53394 20862 53396 20914
rect 53340 20850 53396 20862
rect 53564 20244 53620 20254
rect 53116 20132 53396 20188
rect 53564 20150 53620 20188
rect 53004 20078 53006 20130
rect 53058 20078 53060 20130
rect 52780 20018 52836 20030
rect 52780 19966 52782 20018
rect 52834 19966 52836 20018
rect 52780 18788 52836 19966
rect 52780 18674 52836 18732
rect 52780 18622 52782 18674
rect 52834 18622 52836 18674
rect 52780 18610 52836 18622
rect 53004 18340 53060 20078
rect 53228 20018 53284 20030
rect 53228 19966 53230 20018
rect 53282 19966 53284 20018
rect 52892 18284 53060 18340
rect 53116 19908 53172 19918
rect 52668 18004 52724 18014
rect 52668 17778 52724 17948
rect 52668 17726 52670 17778
rect 52722 17726 52724 17778
rect 52668 17714 52724 17726
rect 52892 16212 52948 18284
rect 52892 16146 52948 16156
rect 53004 17780 53060 17790
rect 53004 16996 53060 17724
rect 53004 16882 53060 16940
rect 53004 16830 53006 16882
rect 53058 16830 53060 16882
rect 52556 15986 52948 15988
rect 52556 15934 52558 15986
rect 52610 15934 52948 15986
rect 52556 15932 52948 15934
rect 52556 15922 52612 15932
rect 52220 15698 52276 15708
rect 52780 15764 52836 15774
rect 51884 15540 51940 15550
rect 51884 15446 51940 15484
rect 52220 15428 52276 15438
rect 52276 15372 52612 15428
rect 52220 15314 52276 15372
rect 52220 15262 52222 15314
rect 52274 15262 52276 15314
rect 52220 14642 52276 15262
rect 52444 15204 52500 15242
rect 52556 15204 52612 15372
rect 52556 15148 52724 15204
rect 52220 14590 52222 14642
rect 52274 14590 52276 14642
rect 52220 14578 52276 14590
rect 52332 15092 52388 15102
rect 52332 14530 52388 15036
rect 52332 14478 52334 14530
rect 52386 14478 52388 14530
rect 51660 14366 51662 14418
rect 51714 14366 51716 14418
rect 51660 14354 51716 14366
rect 51772 14418 51828 14430
rect 51772 14366 51774 14418
rect 51826 14366 51828 14418
rect 51772 13972 51828 14366
rect 51772 13906 51828 13916
rect 52108 14196 52164 14206
rect 52108 13748 52164 14140
rect 52108 13682 52164 13692
rect 52332 13748 52388 14478
rect 51660 13636 51716 13646
rect 51996 13636 52052 13646
rect 51716 13580 51940 13636
rect 51660 13542 51716 13580
rect 51772 12964 51828 12974
rect 51772 12870 51828 12908
rect 51660 12404 51716 12414
rect 51548 12402 51716 12404
rect 51548 12350 51662 12402
rect 51714 12350 51716 12402
rect 51548 12348 51716 12350
rect 51660 12338 51716 12348
rect 51212 12236 51604 12292
rect 51212 12068 51268 12078
rect 51212 11172 51268 12012
rect 51324 11396 51380 11406
rect 51324 11302 51380 11340
rect 51212 11116 51380 11172
rect 51212 10612 51268 10622
rect 51212 10518 51268 10556
rect 51324 10052 51380 11116
rect 51324 9986 51380 9996
rect 51436 10164 51492 10174
rect 51100 9884 51268 9940
rect 51100 9268 51156 9278
rect 51100 9174 51156 9212
rect 51100 9044 51156 9054
rect 51100 6468 51156 8988
rect 51212 8484 51268 9884
rect 51436 9268 51492 10108
rect 51548 9492 51604 12236
rect 51660 11732 51716 11742
rect 51660 11282 51716 11676
rect 51660 11230 51662 11282
rect 51714 11230 51716 11282
rect 51660 11218 51716 11230
rect 51660 11060 51716 11070
rect 51660 10386 51716 11004
rect 51772 10836 51828 10846
rect 51772 10742 51828 10780
rect 51660 10334 51662 10386
rect 51714 10334 51716 10386
rect 51660 10322 51716 10334
rect 51884 9940 51940 13580
rect 52332 13616 52388 13692
rect 51996 10836 52052 13580
rect 52332 12852 52388 12862
rect 52332 12758 52388 12796
rect 52108 12740 52164 12750
rect 52108 12180 52164 12684
rect 52332 12628 52388 12638
rect 52220 12180 52276 12190
rect 52108 12178 52276 12180
rect 52108 12126 52222 12178
rect 52274 12126 52276 12178
rect 52108 12124 52276 12126
rect 51996 10770 52052 10780
rect 52108 11620 52164 11630
rect 52108 11506 52164 11564
rect 52108 11454 52110 11506
rect 52162 11454 52164 11506
rect 52108 10724 52164 11454
rect 52108 10658 52164 10668
rect 51884 9874 51940 9884
rect 52108 10498 52164 10510
rect 52108 10446 52110 10498
rect 52162 10446 52164 10498
rect 51884 9716 51940 9726
rect 51884 9714 52052 9716
rect 51884 9662 51886 9714
rect 51938 9662 52052 9714
rect 51884 9660 52052 9662
rect 51884 9650 51940 9660
rect 51884 9492 51940 9502
rect 51548 9436 51716 9492
rect 51548 9268 51604 9278
rect 51436 9266 51604 9268
rect 51436 9214 51550 9266
rect 51602 9214 51604 9266
rect 51436 9212 51604 9214
rect 51548 9202 51604 9212
rect 51212 8418 51268 8428
rect 51548 8932 51604 8942
rect 51212 8260 51268 8270
rect 51212 8166 51268 8204
rect 51548 7700 51604 8876
rect 51660 8370 51716 9436
rect 51660 8318 51662 8370
rect 51714 8318 51716 8370
rect 51660 8148 51716 8318
rect 51660 8082 51716 8092
rect 51884 8930 51940 9436
rect 51884 8878 51886 8930
rect 51938 8878 51940 8930
rect 51660 7700 51716 7710
rect 51548 7698 51716 7700
rect 51548 7646 51662 7698
rect 51714 7646 51716 7698
rect 51548 7644 51716 7646
rect 51212 6692 51268 6702
rect 51212 6598 51268 6636
rect 51100 6412 51268 6468
rect 51212 5346 51268 6412
rect 51212 5294 51214 5346
rect 51266 5294 51268 5346
rect 51212 5282 51268 5294
rect 51100 5236 51156 5246
rect 50988 5234 51156 5236
rect 50988 5182 51102 5234
rect 51154 5182 51156 5234
rect 50988 5180 51156 5182
rect 51100 5170 51156 5180
rect 51660 5234 51716 7644
rect 51772 7700 51828 7710
rect 51772 6802 51828 7644
rect 51772 6750 51774 6802
rect 51826 6750 51828 6802
rect 51772 6738 51828 6750
rect 51884 6692 51940 8878
rect 51884 6626 51940 6636
rect 51660 5182 51662 5234
rect 51714 5182 51716 5234
rect 51660 5170 51716 5182
rect 51436 4900 51492 4910
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50428 3826 50484 3836
rect 49756 3462 49812 3500
rect 50204 3780 50260 3790
rect 50204 3554 50260 3724
rect 51100 3668 51156 3678
rect 51100 3574 51156 3612
rect 51436 3666 51492 4844
rect 51996 4116 52052 9660
rect 52108 9604 52164 10446
rect 52108 9538 52164 9548
rect 52220 9156 52276 12124
rect 52332 9716 52388 12572
rect 52444 12404 52500 15148
rect 52668 12964 52724 15148
rect 52668 12850 52724 12908
rect 52668 12798 52670 12850
rect 52722 12798 52724 12850
rect 52668 12786 52724 12798
rect 52780 13746 52836 15708
rect 52780 13694 52782 13746
rect 52834 13694 52836 13746
rect 52556 12404 52612 12414
rect 52444 12402 52612 12404
rect 52444 12350 52558 12402
rect 52610 12350 52612 12402
rect 52444 12348 52612 12350
rect 52556 12338 52612 12348
rect 52780 11788 52836 13694
rect 52444 11732 52836 11788
rect 52444 10276 52500 11732
rect 52892 11508 52948 15932
rect 53004 15876 53060 16830
rect 53116 16884 53172 19852
rect 53228 19236 53284 19966
rect 53228 19170 53284 19180
rect 53340 18564 53396 20132
rect 53676 20132 53732 20142
rect 53452 20020 53508 20030
rect 53452 20018 53620 20020
rect 53452 19966 53454 20018
rect 53506 19966 53620 20018
rect 53452 19964 53620 19966
rect 53452 19954 53508 19964
rect 53452 19460 53508 19470
rect 53452 19366 53508 19404
rect 53228 18508 53396 18564
rect 53452 19236 53508 19246
rect 53228 18452 53284 18508
rect 53228 17780 53284 18396
rect 53340 18340 53396 18350
rect 53340 18246 53396 18284
rect 53452 18116 53508 19180
rect 53228 17714 53284 17724
rect 53340 18060 53508 18116
rect 53564 19234 53620 19964
rect 53564 19182 53566 19234
rect 53618 19182 53620 19234
rect 53340 17444 53396 18060
rect 53564 17892 53620 19182
rect 53676 18564 53732 20076
rect 53788 19684 53844 21308
rect 54012 21140 54068 22876
rect 54012 21074 54068 21084
rect 54012 20804 54068 20814
rect 54012 20710 54068 20748
rect 54124 20244 54180 24670
rect 54236 23380 54292 23390
rect 54236 23286 54292 23324
rect 54236 22146 54292 22158
rect 54236 22094 54238 22146
rect 54290 22094 54292 22146
rect 54236 21924 54292 22094
rect 54236 21858 54292 21868
rect 54348 21810 54404 26796
rect 54460 26740 54516 26750
rect 54460 26180 54516 26684
rect 54460 24050 54516 26124
rect 54572 25618 54628 27806
rect 54572 25566 54574 25618
rect 54626 25566 54628 25618
rect 54572 25554 54628 25566
rect 54460 23998 54462 24050
rect 54514 23998 54516 24050
rect 54460 23986 54516 23998
rect 54348 21758 54350 21810
rect 54402 21758 54404 21810
rect 54348 21746 54404 21758
rect 54460 23266 54516 23278
rect 54460 23214 54462 23266
rect 54514 23214 54516 23266
rect 54348 20690 54404 20702
rect 54348 20638 54350 20690
rect 54402 20638 54404 20690
rect 54124 20178 54180 20188
rect 54236 20578 54292 20590
rect 54236 20526 54238 20578
rect 54290 20526 54292 20578
rect 54236 20020 54292 20526
rect 54348 20244 54404 20638
rect 54348 20178 54404 20188
rect 54348 20020 54404 20030
rect 54236 19964 54348 20020
rect 54348 19926 54404 19964
rect 54460 19908 54516 23214
rect 54572 23156 54628 23166
rect 54572 23062 54628 23100
rect 54684 22372 54740 27916
rect 54796 27076 54852 29596
rect 55020 29586 55076 29598
rect 54908 29428 54964 29438
rect 54908 29334 54964 29372
rect 55132 29428 55188 29466
rect 55132 29362 55188 29372
rect 55132 28418 55188 28430
rect 55132 28366 55134 28418
rect 55186 28366 55188 28418
rect 55132 28084 55188 28366
rect 55132 28018 55188 28028
rect 55244 27188 55300 30156
rect 55580 30100 55636 30110
rect 55580 30006 55636 30044
rect 55468 29428 55524 29438
rect 55356 29314 55412 29326
rect 55356 29262 55358 29314
rect 55410 29262 55412 29314
rect 55356 28644 55412 29262
rect 55356 28578 55412 28588
rect 55244 27122 55300 27132
rect 55468 28418 55524 29372
rect 55580 29204 55636 29214
rect 55580 29110 55636 29148
rect 55692 29092 55748 34300
rect 55804 34356 55860 34366
rect 55916 34356 55972 37436
rect 56140 36594 56196 37772
rect 56364 37266 56420 39340
rect 56364 37214 56366 37266
rect 56418 37214 56420 37266
rect 56364 37202 56420 37214
rect 56588 39058 56644 39564
rect 56588 39006 56590 39058
rect 56642 39006 56644 39058
rect 56588 37156 56644 39006
rect 56588 37090 56644 37100
rect 56140 36542 56142 36594
rect 56194 36542 56196 36594
rect 56140 36530 56196 36542
rect 56252 36258 56308 36270
rect 56252 36206 56254 36258
rect 56306 36206 56308 36258
rect 56252 35700 56308 36206
rect 56588 35812 56644 35822
rect 56588 35718 56644 35756
rect 56252 35634 56308 35644
rect 55804 34354 55972 34356
rect 55804 34302 55806 34354
rect 55858 34302 55972 34354
rect 55804 34300 55972 34302
rect 56028 35588 56084 35598
rect 55804 33684 55860 34300
rect 55804 29316 55860 33628
rect 55916 33236 55972 33246
rect 55916 33142 55972 33180
rect 56028 32900 56084 35532
rect 56252 35476 56308 35486
rect 56252 35382 56308 35420
rect 56588 34804 56644 34814
rect 56588 34710 56644 34748
rect 56252 34580 56308 34590
rect 56252 33458 56308 34524
rect 56700 34356 56756 39788
rect 56812 39842 56868 40012
rect 56812 39790 56814 39842
rect 56866 39790 56868 39842
rect 56812 39778 56868 39790
rect 56924 37940 56980 40236
rect 57036 39844 57092 40910
rect 57036 39778 57092 39788
rect 57036 39618 57092 39630
rect 57036 39566 57038 39618
rect 57090 39566 57092 39618
rect 57036 39508 57092 39566
rect 57036 39442 57092 39452
rect 56924 37716 56980 37884
rect 57148 37828 57204 42926
rect 57708 42980 57764 42990
rect 57932 42980 57988 43374
rect 57708 42978 57988 42980
rect 57708 42926 57710 42978
rect 57762 42926 57988 42978
rect 57708 42924 57988 42926
rect 57708 42866 57764 42924
rect 57708 42814 57710 42866
rect 57762 42814 57764 42866
rect 57708 42802 57764 42814
rect 57372 42532 57428 42542
rect 57372 42438 57428 42476
rect 57372 41860 57428 41870
rect 57372 41766 57428 41804
rect 57820 41860 57876 41870
rect 57820 41766 57876 41804
rect 58044 41636 58100 45164
rect 58156 43764 58212 43774
rect 58156 41748 58212 43708
rect 58156 41692 58548 41748
rect 58044 41580 58436 41636
rect 57372 40964 57428 40974
rect 57820 40964 57876 40974
rect 57372 40962 57764 40964
rect 57372 40910 57374 40962
rect 57426 40910 57764 40962
rect 57372 40908 57764 40910
rect 57372 40898 57428 40908
rect 57708 40516 57764 40908
rect 57820 40962 58324 40964
rect 57820 40910 57822 40962
rect 57874 40910 58324 40962
rect 57820 40908 58324 40910
rect 57820 40898 57876 40908
rect 57708 40460 58212 40516
rect 57372 40292 57428 40302
rect 57372 40290 57876 40292
rect 57372 40238 57374 40290
rect 57426 40238 57876 40290
rect 57372 40236 57876 40238
rect 57372 40226 57428 40236
rect 57260 39618 57316 39630
rect 57260 39566 57262 39618
rect 57314 39566 57316 39618
rect 57260 38274 57316 39566
rect 57708 39620 57764 39630
rect 57708 39526 57764 39564
rect 57484 39394 57540 39406
rect 57484 39342 57486 39394
rect 57538 39342 57540 39394
rect 57372 39060 57428 39070
rect 57372 38966 57428 39004
rect 57484 38836 57540 39342
rect 57596 39396 57652 39406
rect 57596 39302 57652 39340
rect 57596 39172 57652 39182
rect 57596 39058 57652 39116
rect 57596 39006 57598 39058
rect 57650 39006 57652 39058
rect 57596 38994 57652 39006
rect 57708 38948 57764 38958
rect 57708 38854 57764 38892
rect 57484 38770 57540 38780
rect 57820 38668 57876 40236
rect 57260 38222 57262 38274
rect 57314 38222 57316 38274
rect 57260 38210 57316 38222
rect 57708 38612 57876 38668
rect 57932 40290 57988 40302
rect 57932 40238 57934 40290
rect 57986 40238 57988 40290
rect 57596 38052 57652 38062
rect 57596 37958 57652 37996
rect 57148 37772 57316 37828
rect 56924 37660 57204 37716
rect 57148 36484 57204 37660
rect 57260 36932 57316 37772
rect 57372 37380 57428 37390
rect 57372 37378 57652 37380
rect 57372 37326 57374 37378
rect 57426 37326 57652 37378
rect 57372 37324 57652 37326
rect 57372 37314 57428 37324
rect 57484 37156 57540 37166
rect 57260 36876 57428 36932
rect 57260 36484 57316 36494
rect 57148 36482 57316 36484
rect 57148 36430 57262 36482
rect 57314 36430 57316 36482
rect 57148 36428 57316 36430
rect 57260 36418 57316 36428
rect 56812 36372 56868 36382
rect 56812 36278 56868 36316
rect 57260 36148 57316 36158
rect 57036 35700 57092 35710
rect 56924 35028 56980 35038
rect 56924 34934 56980 34972
rect 57036 34914 57092 35644
rect 57036 34862 57038 34914
rect 57090 34862 57092 34914
rect 57036 34850 57092 34862
rect 56700 34300 56868 34356
rect 56364 34244 56420 34254
rect 56364 34242 56532 34244
rect 56364 34190 56366 34242
rect 56418 34190 56532 34242
rect 56364 34188 56532 34190
rect 56364 34178 56420 34188
rect 56252 33406 56254 33458
rect 56306 33406 56308 33458
rect 56252 33394 56308 33406
rect 56476 33572 56532 34188
rect 56588 34132 56644 34142
rect 56588 34038 56644 34076
rect 55916 32844 56084 32900
rect 56140 33122 56196 33134
rect 56364 33124 56420 33134
rect 56140 33070 56142 33122
rect 56194 33070 56196 33122
rect 55916 30996 55972 32844
rect 56028 32450 56084 32462
rect 56028 32398 56030 32450
rect 56082 32398 56084 32450
rect 56028 31668 56084 32398
rect 56140 32004 56196 33070
rect 56140 31938 56196 31948
rect 56252 33122 56420 33124
rect 56252 33070 56366 33122
rect 56418 33070 56420 33122
rect 56252 33068 56420 33070
rect 56028 31602 56084 31612
rect 55916 30930 55972 30940
rect 56252 30324 56308 33068
rect 56364 33058 56420 33068
rect 56476 31778 56532 33516
rect 56588 32564 56644 32574
rect 56588 32470 56644 32508
rect 56812 32452 56868 34300
rect 57260 33460 57316 36092
rect 57260 33394 57316 33404
rect 56812 32004 56868 32396
rect 56476 31726 56478 31778
rect 56530 31726 56532 31778
rect 56476 31714 56532 31726
rect 56700 31948 56868 32004
rect 56924 33236 56980 33246
rect 56700 31890 56756 31948
rect 56700 31838 56702 31890
rect 56754 31838 56756 31890
rect 56700 31220 56756 31838
rect 56812 31780 56868 31790
rect 56812 31666 56868 31724
rect 56812 31614 56814 31666
rect 56866 31614 56868 31666
rect 56812 31602 56868 31614
rect 56700 31164 56868 31220
rect 56364 31108 56420 31118
rect 56364 31106 56644 31108
rect 56364 31054 56366 31106
rect 56418 31054 56644 31106
rect 56364 31052 56644 31054
rect 56364 31042 56420 31052
rect 56252 30268 56532 30324
rect 56252 30098 56308 30110
rect 56252 30046 56254 30098
rect 56306 30046 56308 30098
rect 56028 29428 56084 29438
rect 56028 29334 56084 29372
rect 55804 29250 55860 29260
rect 56140 29204 56196 29214
rect 55692 29036 55860 29092
rect 55468 28366 55470 28418
rect 55522 28366 55524 28418
rect 54908 27076 54964 27086
rect 54796 27074 54964 27076
rect 54796 27022 54910 27074
rect 54962 27022 54964 27074
rect 54796 27020 54964 27022
rect 54908 26964 54964 27020
rect 54908 26898 54964 26908
rect 55132 26964 55188 26974
rect 55468 26908 55524 28366
rect 55804 28196 55860 29036
rect 56028 28980 56084 28990
rect 55804 27300 55860 28140
rect 55916 28756 55972 28766
rect 55916 27412 55972 28700
rect 56028 28642 56084 28924
rect 56140 28754 56196 29148
rect 56140 28702 56142 28754
rect 56194 28702 56196 28754
rect 56140 28690 56196 28702
rect 56252 28756 56308 30046
rect 56364 29652 56420 29662
rect 56476 29652 56532 30268
rect 56364 29650 56532 29652
rect 56364 29598 56366 29650
rect 56418 29598 56532 29650
rect 56364 29596 56532 29598
rect 56364 29586 56420 29596
rect 56476 29428 56532 29438
rect 56476 29334 56532 29372
rect 56252 28700 56420 28756
rect 56028 28590 56030 28642
rect 56082 28590 56084 28642
rect 56028 28578 56084 28590
rect 56252 28530 56308 28542
rect 56252 28478 56254 28530
rect 56306 28478 56308 28530
rect 56252 28308 56308 28478
rect 56252 28242 56308 28252
rect 56028 28084 56084 28094
rect 56028 27858 56084 28028
rect 56028 27806 56030 27858
rect 56082 27806 56084 27858
rect 56028 27794 56084 27806
rect 55916 27300 55972 27356
rect 56140 27300 56196 27310
rect 55916 27298 56196 27300
rect 55916 27246 56142 27298
rect 56194 27246 56196 27298
rect 55916 27244 56196 27246
rect 55804 27168 55860 27244
rect 56140 27234 56196 27244
rect 55132 26870 55188 26908
rect 55356 26852 55524 26908
rect 55580 27076 55636 27086
rect 54908 26292 54964 26302
rect 54908 26198 54964 26236
rect 55244 25508 55300 25518
rect 55244 25414 55300 25452
rect 54796 25172 54852 25182
rect 54796 24946 54852 25116
rect 54796 24894 54798 24946
rect 54850 24894 54852 24946
rect 54796 24882 54852 24894
rect 55132 24834 55188 24846
rect 55132 24782 55134 24834
rect 55186 24782 55188 24834
rect 55132 24500 55188 24782
rect 55132 24434 55188 24444
rect 55356 24164 55412 26852
rect 55580 24164 55636 27020
rect 56028 27076 56084 27086
rect 56364 27076 56420 28700
rect 56588 27972 56644 31052
rect 56700 30994 56756 31006
rect 56700 30942 56702 30994
rect 56754 30942 56756 30994
rect 56700 30660 56756 30942
rect 56700 30594 56756 30604
rect 56700 30210 56756 30222
rect 56700 30158 56702 30210
rect 56754 30158 56756 30210
rect 56700 30100 56756 30158
rect 56700 30034 56756 30044
rect 56700 29428 56756 29438
rect 56700 29334 56756 29372
rect 56700 28756 56756 28766
rect 56700 28642 56756 28700
rect 56700 28590 56702 28642
rect 56754 28590 56756 28642
rect 56700 28578 56756 28590
rect 56812 28084 56868 31164
rect 56924 30322 56980 33180
rect 57148 33236 57204 33246
rect 57372 33236 57428 36876
rect 57484 35810 57540 37100
rect 57484 35758 57486 35810
rect 57538 35758 57540 35810
rect 57484 35746 57540 35758
rect 57484 35476 57540 35486
rect 57484 34242 57540 35420
rect 57484 34190 57486 34242
rect 57538 34190 57540 34242
rect 57484 34178 57540 34190
rect 57596 34132 57652 37324
rect 57708 36708 57764 38612
rect 57820 38500 57876 38510
rect 57820 38164 57876 38444
rect 57932 38388 57988 40238
rect 57932 38322 57988 38332
rect 58156 38164 58212 40460
rect 57820 38162 58100 38164
rect 57820 38110 57822 38162
rect 57874 38110 58100 38162
rect 57820 38108 58100 38110
rect 57820 38098 57876 38108
rect 57820 37156 57876 37166
rect 57820 37154 57988 37156
rect 57820 37102 57822 37154
rect 57874 37102 57988 37154
rect 57820 37100 57988 37102
rect 57820 37090 57876 37100
rect 57708 36652 57876 36708
rect 57708 36482 57764 36494
rect 57708 36430 57710 36482
rect 57762 36430 57764 36482
rect 57708 35924 57764 36430
rect 57820 36148 57876 36652
rect 57820 36082 57876 36092
rect 57820 35924 57876 35934
rect 57708 35922 57876 35924
rect 57708 35870 57822 35922
rect 57874 35870 57876 35922
rect 57708 35868 57876 35870
rect 57820 35858 57876 35868
rect 57708 35700 57764 35710
rect 57708 35606 57764 35644
rect 57596 34076 57764 34132
rect 57148 33234 57428 33236
rect 57148 33182 57150 33234
rect 57202 33182 57428 33234
rect 57148 33180 57428 33182
rect 57596 33906 57652 33918
rect 57596 33854 57598 33906
rect 57650 33854 57652 33906
rect 57148 32564 57204 33180
rect 57484 33124 57540 33134
rect 57148 32498 57204 32508
rect 57260 33122 57540 33124
rect 57260 33070 57486 33122
rect 57538 33070 57540 33122
rect 57260 33068 57540 33070
rect 56924 30270 56926 30322
rect 56978 30270 56980 30322
rect 56924 30258 56980 30270
rect 57148 32116 57204 32126
rect 56812 28018 56868 28028
rect 57148 28530 57204 32060
rect 57260 29428 57316 33068
rect 57484 33058 57540 33068
rect 57484 32676 57540 32686
rect 57372 32674 57540 32676
rect 57372 32622 57486 32674
rect 57538 32622 57540 32674
rect 57372 32620 57540 32622
rect 57372 31892 57428 32620
rect 57484 32610 57540 32620
rect 57372 31826 57428 31836
rect 57484 31780 57540 31790
rect 57596 31780 57652 33854
rect 57708 31892 57764 34076
rect 57932 33348 57988 37100
rect 58044 35810 58100 38108
rect 58156 38098 58212 38108
rect 58268 37268 58324 40908
rect 58268 37202 58324 37212
rect 58044 35758 58046 35810
rect 58098 35758 58100 35810
rect 58044 35028 58100 35758
rect 58044 34962 58100 34972
rect 58156 36372 58212 36382
rect 58044 34692 58100 34702
rect 58044 34598 58100 34636
rect 58044 34020 58100 34030
rect 58044 33926 58100 33964
rect 57932 33282 57988 33292
rect 57932 33122 57988 33134
rect 57932 33070 57934 33122
rect 57986 33070 57988 33122
rect 57932 32676 57988 33070
rect 57932 32610 57988 32620
rect 57820 32564 57876 32574
rect 57820 32470 57876 32508
rect 57708 31836 57876 31892
rect 57540 31724 57764 31780
rect 57484 31556 57540 31724
rect 57372 31500 57540 31556
rect 57372 30210 57428 31500
rect 57484 31106 57540 31118
rect 57484 31054 57486 31106
rect 57538 31054 57540 31106
rect 57484 30324 57540 31054
rect 57484 30258 57540 30268
rect 57596 30996 57652 31006
rect 57372 30158 57374 30210
rect 57426 30158 57428 30210
rect 57372 30146 57428 30158
rect 57596 30100 57652 30940
rect 57708 30994 57764 31724
rect 57820 31556 57876 31836
rect 57932 31780 57988 31790
rect 57932 31778 58100 31780
rect 57932 31726 57934 31778
rect 57986 31726 58100 31778
rect 57932 31724 58100 31726
rect 57932 31714 57988 31724
rect 57820 31490 57876 31500
rect 57708 30942 57710 30994
rect 57762 30942 57764 30994
rect 57708 30930 57764 30942
rect 57484 30044 57652 30100
rect 57484 29650 57540 30044
rect 57820 29988 57876 29998
rect 57820 29986 57988 29988
rect 57820 29934 57822 29986
rect 57874 29934 57988 29986
rect 57820 29932 57988 29934
rect 57820 29922 57876 29932
rect 57484 29598 57486 29650
rect 57538 29598 57540 29650
rect 57484 29586 57540 29598
rect 57260 29362 57316 29372
rect 57708 29426 57764 29438
rect 57708 29374 57710 29426
rect 57762 29374 57764 29426
rect 57708 28644 57764 29374
rect 57484 28642 57764 28644
rect 57484 28590 57710 28642
rect 57762 28590 57764 28642
rect 57484 28588 57764 28590
rect 57372 28532 57428 28542
rect 57148 28478 57150 28530
rect 57202 28478 57204 28530
rect 57148 28420 57204 28478
rect 57148 28084 57204 28364
rect 57148 28018 57204 28028
rect 57260 28530 57428 28532
rect 57260 28478 57374 28530
rect 57426 28478 57428 28530
rect 57260 28476 57428 28478
rect 56588 27906 56644 27916
rect 57260 27748 57316 28476
rect 57372 28466 57428 28476
rect 57484 28196 57540 28588
rect 57708 28578 57764 28588
rect 57596 28420 57652 28430
rect 57596 28326 57652 28364
rect 57932 28196 57988 29932
rect 58044 28756 58100 31724
rect 58044 28690 58100 28700
rect 57484 28140 57652 28196
rect 57036 27692 57316 27748
rect 57484 27972 57540 27982
rect 56028 27074 56420 27076
rect 56028 27022 56030 27074
rect 56082 27022 56420 27074
rect 56028 27020 56420 27022
rect 56476 27412 56532 27422
rect 55692 26962 55748 26974
rect 55692 26910 55694 26962
rect 55746 26910 55748 26962
rect 55692 24948 55748 26910
rect 56028 26964 56084 27020
rect 56028 26852 56196 26908
rect 56028 26178 56084 26190
rect 56028 26126 56030 26178
rect 56082 26126 56084 26178
rect 56028 25620 56084 26126
rect 56028 25554 56084 25564
rect 55692 24882 55748 24892
rect 56140 24946 56196 26852
rect 56140 24894 56142 24946
rect 56194 24894 56196 24946
rect 56140 24882 56196 24894
rect 55804 24836 55860 24846
rect 56476 24836 56532 27356
rect 56812 27300 56868 27310
rect 56588 26180 56644 26190
rect 56588 26086 56644 26124
rect 56588 25508 56644 25518
rect 56588 25414 56644 25452
rect 56588 25284 56644 25294
rect 56588 24946 56644 25228
rect 56588 24894 56590 24946
rect 56642 24894 56644 24946
rect 56588 24882 56644 24894
rect 55804 24742 55860 24780
rect 56364 24780 56532 24836
rect 55132 24108 55412 24164
rect 55468 24108 55636 24164
rect 55916 24164 55972 24174
rect 54684 22306 54740 22316
rect 54908 24052 54964 24062
rect 54684 21476 54740 21486
rect 54684 21382 54740 21420
rect 54572 20580 54628 20590
rect 54572 20242 54628 20524
rect 54572 20190 54574 20242
rect 54626 20190 54628 20242
rect 54572 20178 54628 20190
rect 54460 19842 54516 19852
rect 53788 19628 54180 19684
rect 54124 19458 54180 19628
rect 54124 19406 54126 19458
rect 54178 19406 54180 19458
rect 54124 19394 54180 19406
rect 54012 19348 54068 19358
rect 53900 19292 54012 19348
rect 53788 19236 53844 19246
rect 53788 19142 53844 19180
rect 53676 18498 53732 18508
rect 53788 18340 53844 18350
rect 53788 18246 53844 18284
rect 53564 17826 53620 17836
rect 53452 17780 53508 17790
rect 53452 17666 53508 17724
rect 53452 17614 53454 17666
rect 53506 17614 53508 17666
rect 53452 17602 53508 17614
rect 53788 17556 53844 17566
rect 53900 17556 53956 19292
rect 54012 19254 54068 19292
rect 54684 19012 54740 19022
rect 54684 18918 54740 18956
rect 54908 18788 54964 23996
rect 55132 23716 55188 24108
rect 55244 23938 55300 23950
rect 55244 23886 55246 23938
rect 55298 23886 55300 23938
rect 55244 23828 55300 23886
rect 55468 23828 55524 24108
rect 55916 24050 55972 24108
rect 55916 23998 55918 24050
rect 55970 23998 55972 24050
rect 55244 23772 55524 23828
rect 55132 23660 55412 23716
rect 55244 23380 55300 23390
rect 55244 23286 55300 23324
rect 55132 23154 55188 23166
rect 55132 23102 55134 23154
rect 55186 23102 55188 23154
rect 55132 23044 55188 23102
rect 55132 22596 55188 22988
rect 55244 22932 55300 22942
rect 55356 22932 55412 23660
rect 55244 22930 55412 22932
rect 55244 22878 55246 22930
rect 55298 22878 55412 22930
rect 55244 22876 55412 22878
rect 55244 22866 55300 22876
rect 55468 22596 55524 23772
rect 55580 23938 55636 23950
rect 55580 23886 55582 23938
rect 55634 23886 55636 23938
rect 55580 23156 55636 23886
rect 55580 23090 55636 23100
rect 55916 23154 55972 23998
rect 55916 23102 55918 23154
rect 55970 23102 55972 23154
rect 55916 23044 55972 23102
rect 55916 22978 55972 22988
rect 55132 22540 55412 22596
rect 55020 22372 55076 22382
rect 55244 22372 55300 22382
rect 55020 22278 55076 22316
rect 55132 22370 55300 22372
rect 55132 22318 55246 22370
rect 55298 22318 55300 22370
rect 55132 22316 55300 22318
rect 55020 20804 55076 20814
rect 55020 20710 55076 20748
rect 54908 18722 54964 18732
rect 54796 18676 54852 18686
rect 54796 18582 54852 18620
rect 53788 17554 53956 17556
rect 53788 17502 53790 17554
rect 53842 17502 53956 17554
rect 53788 17500 53956 17502
rect 54012 18564 54068 18574
rect 53788 17490 53844 17500
rect 53340 17388 53508 17444
rect 53228 16884 53284 16894
rect 53116 16882 53284 16884
rect 53116 16830 53230 16882
rect 53282 16830 53284 16882
rect 53116 16828 53284 16830
rect 53228 16324 53284 16828
rect 53228 16258 53284 16268
rect 53340 16772 53396 16782
rect 53004 15820 53172 15876
rect 53004 15428 53060 15466
rect 53004 15362 53060 15372
rect 53116 15148 53172 15820
rect 53340 15538 53396 16716
rect 53340 15486 53342 15538
rect 53394 15486 53396 15538
rect 53340 15474 53396 15486
rect 52668 11452 52948 11508
rect 53004 15092 53172 15148
rect 53452 15148 53508 17388
rect 53900 17332 53956 17342
rect 53564 17108 53620 17146
rect 53564 17042 53620 17052
rect 53564 16884 53620 16894
rect 53564 16770 53620 16828
rect 53564 16718 53566 16770
rect 53618 16718 53620 16770
rect 53564 16706 53620 16718
rect 53676 16772 53732 16782
rect 53564 16212 53620 16222
rect 53564 15764 53620 16156
rect 53676 16098 53732 16716
rect 53676 16046 53678 16098
rect 53730 16046 53732 16098
rect 53676 16034 53732 16046
rect 53788 16436 53844 16446
rect 53676 15764 53732 15774
rect 53564 15708 53676 15764
rect 53452 15092 53620 15148
rect 52668 10836 52724 11452
rect 52780 11284 52836 11294
rect 53004 11284 53060 15092
rect 53340 14308 53396 14318
rect 53228 13860 53284 13870
rect 53228 13766 53284 13804
rect 53116 13748 53172 13758
rect 53116 12402 53172 13692
rect 53340 13074 53396 14252
rect 53564 14306 53620 15092
rect 53564 14254 53566 14306
rect 53618 14254 53620 14306
rect 53564 14196 53620 14254
rect 53340 13022 53342 13074
rect 53394 13022 53396 13074
rect 53340 13010 53396 13022
rect 53452 14140 53564 14196
rect 53116 12350 53118 12402
rect 53170 12350 53172 12402
rect 53116 12338 53172 12350
rect 53340 12178 53396 12190
rect 53340 12126 53342 12178
rect 53394 12126 53396 12178
rect 53340 12068 53396 12126
rect 53340 11732 53396 12012
rect 53340 11666 53396 11676
rect 52780 11282 53060 11284
rect 52780 11230 52782 11282
rect 52834 11230 53060 11282
rect 52780 11228 53060 11230
rect 53340 11284 53396 11294
rect 52780 11218 52836 11228
rect 52668 10704 52724 10780
rect 52444 10220 52612 10276
rect 52444 9940 52500 9950
rect 52444 9846 52500 9884
rect 52332 9650 52388 9660
rect 52556 9492 52612 10220
rect 52892 9940 52948 11228
rect 53340 11190 53396 11228
rect 53004 10498 53060 10510
rect 53004 10446 53006 10498
rect 53058 10446 53060 10498
rect 53004 10276 53060 10446
rect 53004 10210 53060 10220
rect 53452 10164 53508 14140
rect 53564 14130 53620 14140
rect 53564 10836 53620 10846
rect 53564 10742 53620 10780
rect 53116 10108 53508 10164
rect 52892 9884 53060 9940
rect 52556 9426 52612 9436
rect 52892 9716 52948 9726
rect 52556 9268 52612 9278
rect 52220 9100 52500 9156
rect 52332 8932 52388 8942
rect 52220 8930 52388 8932
rect 52220 8878 52334 8930
rect 52386 8878 52388 8930
rect 52220 8876 52388 8878
rect 52220 8484 52276 8876
rect 52332 8866 52388 8876
rect 52220 8418 52276 8428
rect 52332 8708 52388 8718
rect 52108 8148 52164 8158
rect 52108 7700 52164 8092
rect 52108 7634 52164 7644
rect 52332 7698 52388 8652
rect 52332 7646 52334 7698
rect 52386 7646 52388 7698
rect 52332 7634 52388 7646
rect 52108 6468 52164 6478
rect 52108 5234 52164 6412
rect 52108 5182 52110 5234
rect 52162 5182 52164 5234
rect 52108 5170 52164 5182
rect 52220 6466 52276 6478
rect 52220 6414 52222 6466
rect 52274 6414 52276 6466
rect 51996 4050 52052 4060
rect 51436 3614 51438 3666
rect 51490 3614 51492 3666
rect 51436 3602 51492 3614
rect 51996 3892 52052 3902
rect 51996 3666 52052 3836
rect 51996 3614 51998 3666
rect 52050 3614 52052 3666
rect 51996 3602 52052 3614
rect 50204 3502 50206 3554
rect 50258 3502 50260 3554
rect 50204 3490 50260 3502
rect 50540 3556 50596 3566
rect 50540 3330 50596 3500
rect 50540 3278 50542 3330
rect 50594 3278 50596 3330
rect 50540 3266 50596 3278
rect 51772 3444 51828 3454
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51772 800 51828 3388
rect 52220 2772 52276 6414
rect 52332 6018 52388 6030
rect 52332 5966 52334 6018
rect 52386 5966 52388 6018
rect 52332 4564 52388 5966
rect 52444 5348 52500 9100
rect 52556 8370 52612 9212
rect 52892 9266 52948 9660
rect 52892 9214 52894 9266
rect 52946 9214 52948 9266
rect 52892 9202 52948 9214
rect 52556 8318 52558 8370
rect 52610 8318 52612 8370
rect 52556 8306 52612 8318
rect 52780 8036 52836 8046
rect 52780 7698 52836 7980
rect 52780 7646 52782 7698
rect 52834 7646 52836 7698
rect 52780 7634 52836 7646
rect 52556 6804 52612 6814
rect 52556 6710 52612 6748
rect 53004 6580 53060 9884
rect 53116 8036 53172 10108
rect 53340 9940 53396 9950
rect 53676 9940 53732 15708
rect 53788 15538 53844 16380
rect 53788 15486 53790 15538
rect 53842 15486 53844 15538
rect 53788 15474 53844 15486
rect 53788 14532 53844 14542
rect 53788 10836 53844 14476
rect 53900 14420 53956 17276
rect 54012 16884 54068 18508
rect 54908 18564 54964 18574
rect 54908 18470 54964 18508
rect 54236 18452 54292 18462
rect 54236 18358 54292 18396
rect 54684 18452 54740 18462
rect 54684 18228 54740 18396
rect 54460 18172 54740 18228
rect 54460 17444 54516 18172
rect 54796 17892 54852 17902
rect 54684 17556 54740 17566
rect 54572 17444 54628 17482
rect 54460 17388 54572 17444
rect 54572 17378 54628 17388
rect 54572 17220 54628 17230
rect 54460 17108 54516 17118
rect 54460 16994 54516 17052
rect 54460 16942 54462 16994
rect 54514 16942 54516 16994
rect 54460 16930 54516 16942
rect 54012 16818 54068 16828
rect 54124 16548 54180 16558
rect 54124 16324 54180 16492
rect 54012 16322 54180 16324
rect 54012 16270 54126 16322
rect 54178 16270 54180 16322
rect 54012 16268 54180 16270
rect 54012 15540 54068 16268
rect 54124 16258 54180 16268
rect 54012 15474 54068 15484
rect 54124 16100 54180 16110
rect 54124 14868 54180 16044
rect 54572 15538 54628 17164
rect 54684 16994 54740 17500
rect 54684 16942 54686 16994
rect 54738 16942 54740 16994
rect 54684 16930 54740 16942
rect 54684 16212 54740 16222
rect 54684 16118 54740 16156
rect 54572 15486 54574 15538
rect 54626 15486 54628 15538
rect 54572 15474 54628 15486
rect 54684 15428 54740 15438
rect 54684 15334 54740 15372
rect 54236 15314 54292 15326
rect 54236 15262 54238 15314
rect 54290 15262 54292 15314
rect 54236 15092 54292 15262
rect 54236 15026 54292 15036
rect 54684 14980 54740 14990
rect 54124 14812 54628 14868
rect 53900 14418 54068 14420
rect 53900 14366 53902 14418
rect 53954 14366 54068 14418
rect 53900 14364 54068 14366
rect 53900 14354 53956 14364
rect 53900 13524 53956 13534
rect 53900 13430 53956 13468
rect 54012 11788 54068 14364
rect 54348 14306 54404 14318
rect 54348 14254 54350 14306
rect 54402 14254 54404 14306
rect 54236 13636 54292 13646
rect 54236 13542 54292 13580
rect 54124 12850 54180 12862
rect 54124 12798 54126 12850
rect 54178 12798 54180 12850
rect 54124 12740 54180 12798
rect 54124 12180 54180 12684
rect 54348 12628 54404 14254
rect 54460 13748 54516 13758
rect 54460 12850 54516 13692
rect 54460 12798 54462 12850
rect 54514 12798 54516 12850
rect 54460 12786 54516 12798
rect 54348 12562 54404 12572
rect 54236 12180 54292 12190
rect 54124 12178 54292 12180
rect 54124 12126 54238 12178
rect 54290 12126 54292 12178
rect 54124 12124 54292 12126
rect 54236 12114 54292 12124
rect 54348 12068 54404 12078
rect 53900 11732 54068 11788
rect 54236 11956 54292 11966
rect 53900 11396 53956 11732
rect 53900 11340 54180 11396
rect 54124 11282 54180 11340
rect 54124 11230 54126 11282
rect 54178 11230 54180 11282
rect 53900 10836 53956 10846
rect 53788 10834 53956 10836
rect 53788 10782 53902 10834
rect 53954 10782 53956 10834
rect 53788 10780 53956 10782
rect 53900 10386 53956 10780
rect 53900 10334 53902 10386
rect 53954 10334 53956 10386
rect 53900 10322 53956 10334
rect 53340 9938 53732 9940
rect 53340 9886 53342 9938
rect 53394 9886 53732 9938
rect 53340 9884 53732 9886
rect 53340 9874 53396 9884
rect 53676 9268 53732 9884
rect 53676 9136 53732 9212
rect 53788 10052 53844 10062
rect 53788 9938 53844 9996
rect 53788 9886 53790 9938
rect 53842 9886 53844 9938
rect 53788 9044 53844 9886
rect 54012 9268 54068 9278
rect 53788 8988 53956 9044
rect 53228 8932 53284 8942
rect 53228 8930 53396 8932
rect 53228 8878 53230 8930
rect 53282 8878 53396 8930
rect 53228 8876 53396 8878
rect 53228 8866 53284 8876
rect 53340 8820 53396 8876
rect 53788 8820 53844 8830
rect 53340 8764 53620 8820
rect 53116 7970 53172 7980
rect 53228 8708 53284 8718
rect 53004 6514 53060 6524
rect 53116 7812 53172 7822
rect 53116 6130 53172 7756
rect 53228 7698 53284 8652
rect 53340 8372 53396 8382
rect 53340 8278 53396 8316
rect 53228 7646 53230 7698
rect 53282 7646 53284 7698
rect 53228 7634 53284 7646
rect 53452 8260 53508 8270
rect 53452 6690 53508 8204
rect 53564 7700 53620 8764
rect 53788 8370 53844 8764
rect 53788 8318 53790 8370
rect 53842 8318 53844 8370
rect 53788 8306 53844 8318
rect 53564 7634 53620 7644
rect 53452 6638 53454 6690
rect 53506 6638 53508 6690
rect 53452 6626 53508 6638
rect 53564 6692 53620 6702
rect 53116 6078 53118 6130
rect 53170 6078 53172 6130
rect 53116 6066 53172 6078
rect 53564 6130 53620 6636
rect 53564 6078 53566 6130
rect 53618 6078 53620 6130
rect 53564 6066 53620 6078
rect 52444 5282 52500 5292
rect 53340 5348 53396 5358
rect 53340 5234 53396 5292
rect 53340 5182 53342 5234
rect 53394 5182 53396 5234
rect 53340 5170 53396 5182
rect 53788 5348 53844 5358
rect 52444 5124 52500 5134
rect 52444 5030 52500 5068
rect 52332 4498 52388 4508
rect 53788 4562 53844 5292
rect 53788 4510 53790 4562
rect 53842 4510 53844 4562
rect 53788 4498 53844 4510
rect 52556 4340 52612 4350
rect 52556 4004 52612 4284
rect 52556 3938 52612 3948
rect 52892 4338 52948 4350
rect 52892 4286 52894 4338
rect 52946 4286 52948 4338
rect 52892 4228 52948 4286
rect 52892 3668 52948 4172
rect 52892 3602 52948 3612
rect 53452 3666 53508 3678
rect 53452 3614 53454 3666
rect 53506 3614 53508 3666
rect 52780 3556 52836 3566
rect 52780 3462 52836 3500
rect 53452 3444 53508 3614
rect 53452 3378 53508 3388
rect 52220 2706 52276 2716
rect 53900 1540 53956 8988
rect 54012 7698 54068 9212
rect 54012 7646 54014 7698
rect 54066 7646 54068 7698
rect 54012 7634 54068 7646
rect 54012 6692 54068 6702
rect 54124 6692 54180 11230
rect 54236 10836 54292 11900
rect 54348 11394 54404 12012
rect 54348 11342 54350 11394
rect 54402 11342 54404 11394
rect 54348 11330 54404 11342
rect 54348 10836 54404 10846
rect 54236 10834 54404 10836
rect 54236 10782 54350 10834
rect 54402 10782 54404 10834
rect 54236 10780 54404 10782
rect 54348 10770 54404 10780
rect 54460 10386 54516 10398
rect 54460 10334 54462 10386
rect 54514 10334 54516 10386
rect 54236 9602 54292 9614
rect 54236 9550 54238 9602
rect 54290 9550 54292 9602
rect 54236 8260 54292 9550
rect 54348 9268 54404 9278
rect 54348 9174 54404 9212
rect 54236 8194 54292 8204
rect 54236 8036 54292 8046
rect 54236 7942 54292 7980
rect 54348 7700 54404 7710
rect 54460 7700 54516 10334
rect 54572 9268 54628 14812
rect 54684 12852 54740 14924
rect 54684 9828 54740 12796
rect 54796 11396 54852 17836
rect 55132 17556 55188 22316
rect 55244 22306 55300 22316
rect 55244 21586 55300 21598
rect 55244 21534 55246 21586
rect 55298 21534 55300 21586
rect 55244 19908 55300 21534
rect 55244 19842 55300 19852
rect 55356 19684 55412 22540
rect 55468 22530 55524 22540
rect 55692 22596 55748 22606
rect 55468 22370 55524 22382
rect 55468 22318 55470 22370
rect 55522 22318 55524 22370
rect 55468 20244 55524 22318
rect 55692 22370 55748 22540
rect 55804 22484 55860 22494
rect 55804 22390 55860 22428
rect 55692 22318 55694 22370
rect 55746 22318 55748 22370
rect 55692 22306 55748 22318
rect 55692 22148 55748 22158
rect 55580 21698 55636 21710
rect 55580 21646 55582 21698
rect 55634 21646 55636 21698
rect 55580 20692 55636 21646
rect 55580 20626 55636 20636
rect 55692 21588 55748 22092
rect 55916 22146 55972 22158
rect 55916 22094 55918 22146
rect 55970 22094 55972 22146
rect 55916 22036 55972 22094
rect 55916 21970 55972 21980
rect 56364 21868 56420 24780
rect 56588 23940 56644 23950
rect 56588 23846 56644 23884
rect 56476 23268 56532 23278
rect 56476 23154 56532 23212
rect 56476 23102 56478 23154
rect 56530 23102 56532 23154
rect 56476 23044 56532 23102
rect 56476 22978 56532 22988
rect 56588 22596 56644 22606
rect 56588 22502 56644 22540
rect 56700 22148 56756 22158
rect 56700 22054 56756 22092
rect 56364 21812 56532 21868
rect 56364 21700 56420 21710
rect 56364 21606 56420 21644
rect 55580 20244 55636 20254
rect 55468 20242 55636 20244
rect 55468 20190 55582 20242
rect 55634 20190 55636 20242
rect 55468 20188 55636 20190
rect 55580 20178 55636 20188
rect 55020 17500 55188 17556
rect 55244 19628 55412 19684
rect 55468 20018 55524 20030
rect 55468 19966 55470 20018
rect 55522 19966 55524 20018
rect 55468 19908 55524 19966
rect 54908 17444 54964 17454
rect 54908 17350 54964 17388
rect 54908 17108 54964 17118
rect 55020 17108 55076 17500
rect 54908 17106 55076 17108
rect 54908 17054 54910 17106
rect 54962 17054 55076 17106
rect 54908 17052 55076 17054
rect 54908 17042 54964 17052
rect 55020 16882 55076 16894
rect 55020 16830 55022 16882
rect 55074 16830 55076 16882
rect 55020 16660 55076 16830
rect 54908 15876 54964 15886
rect 54908 15426 54964 15820
rect 54908 15374 54910 15426
rect 54962 15374 54964 15426
rect 54908 15362 54964 15374
rect 55020 15148 55076 16604
rect 55020 15092 55188 15148
rect 54908 14532 54964 14542
rect 54908 13746 54964 14476
rect 54908 13694 54910 13746
rect 54962 13694 54964 13746
rect 54908 13636 54964 13694
rect 54908 12628 54964 13580
rect 55020 13748 55076 13758
rect 55020 12852 55076 13692
rect 55132 13186 55188 15092
rect 55132 13134 55134 13186
rect 55186 13134 55188 13186
rect 55132 13122 55188 13134
rect 55244 13076 55300 19628
rect 55468 19236 55524 19852
rect 55356 19180 55524 19236
rect 55692 19794 55748 21532
rect 56028 20690 56084 20702
rect 56028 20638 56030 20690
rect 56082 20638 56084 20690
rect 56028 20244 56084 20638
rect 56028 20178 56084 20188
rect 56364 20580 56420 20590
rect 55692 19742 55694 19794
rect 55746 19742 55748 19794
rect 55356 17220 55412 19180
rect 55468 19012 55524 19050
rect 55468 18946 55524 18956
rect 55692 18340 55748 19742
rect 55804 20020 55860 20030
rect 55804 19796 55860 19964
rect 55916 19796 55972 19806
rect 55804 19794 55972 19796
rect 55804 19742 55918 19794
rect 55970 19742 55972 19794
rect 55804 19740 55972 19742
rect 55804 19124 55860 19740
rect 55916 19730 55972 19740
rect 55804 19030 55860 19068
rect 56252 19012 56308 19022
rect 55356 17154 55412 17164
rect 55468 18284 55748 18340
rect 55804 18564 55860 18574
rect 55804 18450 55860 18508
rect 55804 18398 55806 18450
rect 55858 18398 55860 18450
rect 55468 16996 55524 18284
rect 55580 18116 55636 18126
rect 55580 17890 55636 18060
rect 55580 17838 55582 17890
rect 55634 17838 55636 17890
rect 55580 17826 55636 17838
rect 55692 17556 55748 17566
rect 55804 17556 55860 18398
rect 55916 18562 55972 18574
rect 55916 18510 55918 18562
rect 55970 18510 55972 18562
rect 55916 18452 55972 18510
rect 55916 18386 55972 18396
rect 56252 18004 56308 18956
rect 56252 17938 56308 17948
rect 56364 18450 56420 20524
rect 56476 20132 56532 21812
rect 56700 21588 56756 21598
rect 56700 21494 56756 21532
rect 56588 21364 56644 21374
rect 56588 20914 56644 21308
rect 56588 20862 56590 20914
rect 56642 20862 56644 20914
rect 56588 20850 56644 20862
rect 56476 18676 56532 20076
rect 56700 20132 56756 20142
rect 56700 20038 56756 20076
rect 56588 19906 56644 19918
rect 56588 19854 56590 19906
rect 56642 19854 56644 19906
rect 56588 19236 56644 19854
rect 56812 19348 56868 27244
rect 57036 24052 57092 27692
rect 57148 26852 57204 26862
rect 57148 26758 57204 26796
rect 57484 26852 57540 27916
rect 57484 26758 57540 26796
rect 57484 26066 57540 26078
rect 57484 26014 57486 26066
rect 57538 26014 57540 26066
rect 57484 25060 57540 26014
rect 57484 24994 57540 25004
rect 57484 24834 57540 24846
rect 57484 24782 57486 24834
rect 57538 24782 57540 24834
rect 57260 24724 57316 24734
rect 57148 24052 57204 24062
rect 57036 24050 57204 24052
rect 57036 23998 57150 24050
rect 57202 23998 57204 24050
rect 57036 23996 57204 23998
rect 57148 23986 57204 23996
rect 57036 23882 57092 23894
rect 57036 23830 57038 23882
rect 57090 23830 57092 23882
rect 56924 22260 56980 22270
rect 56924 22166 56980 22204
rect 56812 19282 56868 19292
rect 56588 19170 56644 19180
rect 56924 19124 56980 19134
rect 56924 19030 56980 19068
rect 57036 18676 57092 23830
rect 57148 23716 57204 23726
rect 57148 23622 57204 23660
rect 57260 23548 57316 24668
rect 57484 24164 57540 24782
rect 57596 24834 57652 28140
rect 57708 28140 57988 28196
rect 57708 26628 57764 28140
rect 57820 27972 57876 27982
rect 57820 27878 57876 27916
rect 57932 27188 57988 27198
rect 57932 27094 57988 27132
rect 57708 25508 57764 26572
rect 57820 26852 57876 26862
rect 57820 26066 57876 26796
rect 58044 26178 58100 26190
rect 58044 26126 58046 26178
rect 58098 26126 58100 26178
rect 57820 26014 57822 26066
rect 57874 26014 57876 26066
rect 57820 25956 57876 26014
rect 57820 25890 57876 25900
rect 57932 26068 57988 26078
rect 57708 25452 57876 25508
rect 57708 25284 57764 25294
rect 57708 25190 57764 25228
rect 57596 24782 57598 24834
rect 57650 24782 57652 24834
rect 57596 24770 57652 24782
rect 57484 24098 57540 24108
rect 57708 24722 57764 24734
rect 57708 24670 57710 24722
rect 57762 24670 57764 24722
rect 57484 23940 57540 23950
rect 56476 18544 56532 18620
rect 56812 18620 57036 18676
rect 56700 18564 56756 18574
rect 56364 18398 56366 18450
rect 56418 18398 56420 18450
rect 55748 17500 55860 17556
rect 56252 17554 56308 17566
rect 56252 17502 56254 17554
rect 56306 17502 56308 17554
rect 55692 17462 55748 17500
rect 55356 16940 55524 16996
rect 55580 17444 55636 17454
rect 55356 16100 55412 16940
rect 55356 15874 55412 16044
rect 55356 15822 55358 15874
rect 55410 15822 55412 15874
rect 55356 15810 55412 15822
rect 55468 16098 55524 16110
rect 55468 16046 55470 16098
rect 55522 16046 55524 16098
rect 55468 15428 55524 16046
rect 55580 16100 55636 17388
rect 56252 17444 56308 17502
rect 56252 17378 56308 17388
rect 55916 16994 55972 17006
rect 55916 16942 55918 16994
rect 55970 16942 55972 16994
rect 55916 16884 55972 16942
rect 55916 16818 55972 16828
rect 56252 16882 56308 16894
rect 56252 16830 56254 16882
rect 56306 16830 56308 16882
rect 55804 16100 55860 16110
rect 55580 16098 55860 16100
rect 55580 16046 55806 16098
rect 55858 16046 55860 16098
rect 55580 16044 55860 16046
rect 55468 15296 55524 15372
rect 55580 15540 55636 15550
rect 55580 15148 55636 15484
rect 55468 15092 55636 15148
rect 55692 15092 55748 15102
rect 55356 14642 55412 14654
rect 55356 14590 55358 14642
rect 55410 14590 55412 14642
rect 55356 14196 55412 14590
rect 55356 14130 55412 14140
rect 55468 13076 55524 15092
rect 55692 14998 55748 15036
rect 55692 14420 55748 14430
rect 55692 13748 55748 14364
rect 55804 13748 55860 16044
rect 56252 15876 56308 16830
rect 56252 15810 56308 15820
rect 55916 15316 55972 15326
rect 55916 15222 55972 15260
rect 56364 15316 56420 18398
rect 56476 17668 56532 17678
rect 56476 17666 56644 17668
rect 56476 17614 56478 17666
rect 56530 17614 56644 17666
rect 56476 17612 56644 17614
rect 56476 17556 56532 17612
rect 56476 17490 56532 17500
rect 56588 15986 56644 17612
rect 56588 15934 56590 15986
rect 56642 15934 56644 15986
rect 56588 15922 56644 15934
rect 56700 17106 56756 18508
rect 56812 17890 56868 18620
rect 57036 18610 57092 18620
rect 57148 23492 57316 23548
rect 57372 23714 57428 23726
rect 57372 23662 57374 23714
rect 57426 23662 57428 23714
rect 57148 18564 57204 23492
rect 57372 23380 57428 23662
rect 57372 22820 57428 23324
rect 57484 23378 57540 23884
rect 57484 23326 57486 23378
rect 57538 23326 57540 23378
rect 57484 23314 57540 23326
rect 57708 23380 57764 24670
rect 57820 24050 57876 25452
rect 57932 25506 57988 26012
rect 57932 25454 57934 25506
rect 57986 25454 57988 25506
rect 57932 25442 57988 25454
rect 58044 24948 58100 26126
rect 57820 23998 57822 24050
rect 57874 23998 57876 24050
rect 57820 23986 57876 23998
rect 57932 24892 58100 24948
rect 57372 22754 57428 22764
rect 57484 23156 57540 23166
rect 57484 21810 57540 23100
rect 57484 21758 57486 21810
rect 57538 21758 57540 21810
rect 57484 21746 57540 21758
rect 57596 22370 57652 22382
rect 57596 22318 57598 22370
rect 57650 22318 57652 22370
rect 57260 21588 57316 21598
rect 57260 21026 57316 21532
rect 57596 21588 57652 22318
rect 57708 22260 57764 23324
rect 57820 23268 57876 23278
rect 57932 23268 57988 24892
rect 57820 23266 57988 23268
rect 57820 23214 57822 23266
rect 57874 23214 57988 23266
rect 57820 23212 57988 23214
rect 57820 23202 57876 23212
rect 57820 22260 57876 22270
rect 57708 22258 57876 22260
rect 57708 22206 57822 22258
rect 57874 22206 57876 22258
rect 57708 22204 57876 22206
rect 57820 22194 57876 22204
rect 57708 21588 57764 21598
rect 57652 21586 57764 21588
rect 57652 21534 57710 21586
rect 57762 21534 57764 21586
rect 57652 21532 57764 21534
rect 57596 21456 57652 21532
rect 57708 21522 57764 21532
rect 57260 20974 57262 21026
rect 57314 20974 57316 21026
rect 57260 20962 57316 20974
rect 57708 21028 57764 21038
rect 57372 20804 57428 20814
rect 57372 20710 57428 20748
rect 57484 20132 57540 20142
rect 57484 20038 57540 20076
rect 57708 19346 57764 20972
rect 57820 20916 57876 20926
rect 57820 20822 57876 20860
rect 57932 20580 57988 23212
rect 57932 20514 57988 20524
rect 58044 24722 58100 24734
rect 58044 24670 58046 24722
rect 58098 24670 58100 24722
rect 58044 24052 58100 24670
rect 58044 20356 58100 23996
rect 57820 20300 58100 20356
rect 57820 20242 57876 20300
rect 57820 20190 57822 20242
rect 57874 20190 57876 20242
rect 57820 20178 57876 20190
rect 57708 19294 57710 19346
rect 57762 19294 57764 19346
rect 57260 19124 57316 19134
rect 57260 19030 57316 19068
rect 57484 18564 57540 18574
rect 57148 18562 57540 18564
rect 57148 18510 57486 18562
rect 57538 18510 57540 18562
rect 57148 18508 57540 18510
rect 57484 18228 57540 18508
rect 57708 18564 57764 19294
rect 58044 20132 58100 20142
rect 57820 18676 57876 18686
rect 57820 18582 57876 18620
rect 57708 18498 57764 18508
rect 57484 18162 57540 18172
rect 56812 17838 56814 17890
rect 56866 17838 56868 17890
rect 56812 17826 56868 17838
rect 57372 17668 57428 17678
rect 57372 17554 57428 17612
rect 57372 17502 57374 17554
rect 57426 17502 57428 17554
rect 57372 17490 57428 17502
rect 56700 17054 56702 17106
rect 56754 17054 56756 17106
rect 56588 15540 56644 15550
rect 56588 15446 56644 15484
rect 56364 15250 56420 15260
rect 56140 15202 56196 15214
rect 56140 15150 56142 15202
rect 56194 15150 56196 15202
rect 56028 14530 56084 14542
rect 56028 14478 56030 14530
rect 56082 14478 56084 14530
rect 56028 14308 56084 14478
rect 56140 14532 56196 15150
rect 56700 15148 56756 17054
rect 57708 17444 57764 17454
rect 57484 16996 57540 17006
rect 57484 16902 57540 16940
rect 57708 16884 57764 17388
rect 57596 16882 57764 16884
rect 57596 16830 57710 16882
rect 57762 16830 57764 16882
rect 57596 16828 57764 16830
rect 57372 16324 57428 16334
rect 57372 16210 57428 16268
rect 57372 16158 57374 16210
rect 57426 16158 57428 16210
rect 56924 15876 56980 15886
rect 56924 15782 56980 15820
rect 56140 14466 56196 14476
rect 56476 15092 56756 15148
rect 57260 15316 57316 15326
rect 56028 14242 56084 14252
rect 56364 13972 56420 13982
rect 56140 13860 56196 13870
rect 55804 13692 56084 13748
rect 55692 13616 55748 13692
rect 56028 13634 56084 13692
rect 56028 13582 56030 13634
rect 56082 13582 56084 13634
rect 55580 13524 55636 13534
rect 55580 13300 55636 13468
rect 55580 13234 55636 13244
rect 55916 13188 55972 13198
rect 55692 13076 55748 13086
rect 55244 13020 55412 13076
rect 55468 13074 55748 13076
rect 55468 13022 55694 13074
rect 55746 13022 55748 13074
rect 55468 13020 55748 13022
rect 55132 12852 55188 12862
rect 55020 12850 55188 12852
rect 55020 12798 55134 12850
rect 55186 12798 55188 12850
rect 55020 12796 55188 12798
rect 55132 12786 55188 12796
rect 55244 12850 55300 12862
rect 55244 12798 55246 12850
rect 55298 12798 55300 12850
rect 55244 12628 55300 12798
rect 54908 12572 55300 12628
rect 54796 10834 54852 11340
rect 55132 12292 55188 12302
rect 55356 12292 55412 13020
rect 55692 13010 55748 13020
rect 55804 13076 55860 13086
rect 55132 12290 55412 12292
rect 55132 12238 55134 12290
rect 55186 12238 55412 12290
rect 55132 12236 55412 12238
rect 54796 10782 54798 10834
rect 54850 10782 54852 10834
rect 54796 10770 54852 10782
rect 54908 11172 54964 11182
rect 54908 10500 54964 11116
rect 54908 10434 54964 10444
rect 55132 9940 55188 12236
rect 55692 12178 55748 12190
rect 55692 12126 55694 12178
rect 55746 12126 55748 12178
rect 55692 12068 55748 12126
rect 55692 12002 55748 12012
rect 55356 11620 55412 11630
rect 55356 11506 55412 11564
rect 55356 11454 55358 11506
rect 55410 11454 55412 11506
rect 55356 11442 55412 11454
rect 55692 11618 55748 11630
rect 55692 11566 55694 11618
rect 55746 11566 55748 11618
rect 55356 10836 55412 10846
rect 55356 10742 55412 10780
rect 55692 10834 55748 11566
rect 55804 11506 55860 13020
rect 55804 11454 55806 11506
rect 55858 11454 55860 11506
rect 55804 11442 55860 11454
rect 55692 10782 55694 10834
rect 55746 10782 55748 10834
rect 55692 10770 55748 10782
rect 55580 9940 55636 9950
rect 55132 9938 55580 9940
rect 55132 9886 55134 9938
rect 55186 9886 55580 9938
rect 55132 9884 55580 9886
rect 55636 9884 55748 9940
rect 55132 9874 55188 9884
rect 54684 9772 55076 9828
rect 55580 9808 55636 9884
rect 54684 9602 54740 9614
rect 54684 9550 54686 9602
rect 54738 9550 54740 9602
rect 54684 9492 54740 9550
rect 54684 9426 54740 9436
rect 54684 9268 54740 9278
rect 54572 9266 54740 9268
rect 54572 9214 54686 9266
rect 54738 9214 54740 9266
rect 54572 9212 54740 9214
rect 54684 8372 54740 9212
rect 54684 8306 54740 8316
rect 55020 9268 55076 9772
rect 55468 9380 55524 9390
rect 55132 9268 55188 9278
rect 55020 9266 55188 9268
rect 55020 9214 55134 9266
rect 55186 9214 55188 9266
rect 55020 9212 55188 9214
rect 54348 7698 54516 7700
rect 54348 7646 54350 7698
rect 54402 7646 54516 7698
rect 54348 7644 54516 7646
rect 54348 7634 54404 7644
rect 54460 6804 54516 7644
rect 54796 8036 54852 8046
rect 54796 7698 54852 7980
rect 54796 7646 54798 7698
rect 54850 7646 54852 7698
rect 54796 7634 54852 7646
rect 54460 6738 54516 6748
rect 54012 6690 54124 6692
rect 54012 6638 54014 6690
rect 54066 6638 54124 6690
rect 54012 6636 54124 6638
rect 54012 6626 54068 6636
rect 54124 5236 54180 6636
rect 54908 6692 54964 6702
rect 54908 6598 54964 6636
rect 54236 6580 54292 6590
rect 54236 6130 54292 6524
rect 54460 6580 54516 6590
rect 54460 6486 54516 6524
rect 55020 6468 55076 9212
rect 55132 9202 55188 9212
rect 55020 6402 55076 6412
rect 55132 8372 55188 8382
rect 54236 6078 54238 6130
rect 54290 6078 54292 6130
rect 54236 6066 54292 6078
rect 54684 6132 54740 6142
rect 54684 6038 54740 6076
rect 55132 6130 55188 8316
rect 55356 8370 55412 8382
rect 55356 8318 55358 8370
rect 55410 8318 55412 8370
rect 55356 8148 55412 8318
rect 55356 8082 55412 8092
rect 55244 7588 55300 7598
rect 55244 7494 55300 7532
rect 55356 6580 55412 6590
rect 55356 6486 55412 6524
rect 55132 6078 55134 6130
rect 55186 6078 55188 6130
rect 55132 6066 55188 6078
rect 54572 5348 54628 5358
rect 54236 5236 54292 5246
rect 54124 5234 54292 5236
rect 54124 5182 54238 5234
rect 54290 5182 54292 5234
rect 54124 5180 54292 5182
rect 54236 5170 54292 5180
rect 54572 5234 54628 5292
rect 54572 5182 54574 5234
rect 54626 5182 54628 5234
rect 54572 5170 54628 5182
rect 55020 4900 55076 4910
rect 54908 4898 55076 4900
rect 54908 4846 55022 4898
rect 55074 4846 55076 4898
rect 54908 4844 55076 4846
rect 54124 4228 54180 4238
rect 54124 4134 54180 4172
rect 54908 4228 54964 4844
rect 55020 4834 55076 4844
rect 54908 4162 54964 4172
rect 55356 4226 55412 4238
rect 55356 4174 55358 4226
rect 55410 4174 55412 4226
rect 55244 3668 55300 3678
rect 55244 3574 55300 3612
rect 55356 2772 55412 4174
rect 55356 2706 55412 2716
rect 55468 1652 55524 9324
rect 55692 9266 55748 9884
rect 55692 9214 55694 9266
rect 55746 9214 55748 9266
rect 55692 9202 55748 9214
rect 55916 9268 55972 13132
rect 56028 12402 56084 13582
rect 56140 13074 56196 13804
rect 56140 13022 56142 13074
rect 56194 13022 56196 13074
rect 56140 13010 56196 13022
rect 56028 12350 56030 12402
rect 56082 12350 56084 12402
rect 56028 12338 56084 12350
rect 56364 11618 56420 13916
rect 56364 11566 56366 11618
rect 56418 11566 56420 11618
rect 56364 11554 56420 11566
rect 56252 11508 56308 11518
rect 56252 11414 56308 11452
rect 56476 11060 56532 15092
rect 57036 14868 57092 14878
rect 56700 14420 56756 14430
rect 57036 14420 57092 14812
rect 56700 14326 56756 14364
rect 56924 14418 57092 14420
rect 56924 14366 57038 14418
rect 57090 14366 57092 14418
rect 56924 14364 57092 14366
rect 56588 12404 56644 12414
rect 56588 12310 56644 12348
rect 56924 11732 56980 14364
rect 57036 14354 57092 14364
rect 57148 14644 57204 14654
rect 57036 12852 57092 12862
rect 57036 12758 57092 12796
rect 57148 12068 57204 14588
rect 56924 11666 56980 11676
rect 57036 12012 57204 12068
rect 57260 12852 57316 15260
rect 57372 13076 57428 16158
rect 57484 15876 57540 15886
rect 57484 15538 57540 15820
rect 57484 15486 57486 15538
rect 57538 15486 57540 15538
rect 57484 15474 57540 15486
rect 57596 15316 57652 16828
rect 57708 16818 57764 16828
rect 57820 15874 57876 15886
rect 57820 15822 57822 15874
rect 57874 15822 57876 15874
rect 57820 15764 57876 15822
rect 57820 15698 57876 15708
rect 57932 15876 57988 15886
rect 57484 15260 57652 15316
rect 57708 15316 57764 15326
rect 57484 13970 57540 15260
rect 57708 14980 57764 15260
rect 57708 14914 57764 14924
rect 57596 14532 57652 14542
rect 57596 14418 57652 14476
rect 57932 14530 57988 15820
rect 57932 14478 57934 14530
rect 57986 14478 57988 14530
rect 57932 14466 57988 14478
rect 57596 14366 57598 14418
rect 57650 14366 57652 14418
rect 57596 14354 57652 14366
rect 57484 13918 57486 13970
rect 57538 13918 57540 13970
rect 57484 13906 57540 13918
rect 57820 13748 57876 13758
rect 57820 13746 57988 13748
rect 57820 13694 57822 13746
rect 57874 13694 57988 13746
rect 57820 13692 57988 13694
rect 57820 13682 57876 13692
rect 57820 13076 57876 13086
rect 57372 13020 57764 13076
rect 57372 12852 57428 12862
rect 57260 12850 57428 12852
rect 57260 12798 57374 12850
rect 57426 12798 57428 12850
rect 57260 12796 57428 12798
rect 56700 11396 56756 11406
rect 56700 11302 56756 11340
rect 56476 10994 56532 11004
rect 56588 10612 56644 10622
rect 56476 10500 56532 10510
rect 56476 10406 56532 10444
rect 56252 9940 56308 9950
rect 56252 9846 56308 9884
rect 55916 9202 55972 9212
rect 56140 9268 56196 9278
rect 56140 9174 56196 9212
rect 56588 8932 56644 10556
rect 57036 10052 57092 12012
rect 56700 9996 57092 10052
rect 57148 11844 57204 11854
rect 57148 11506 57204 11788
rect 57148 11454 57150 11506
rect 57202 11454 57204 11506
rect 56700 9938 56756 9996
rect 56700 9886 56702 9938
rect 56754 9886 56756 9938
rect 56700 9380 56756 9886
rect 56700 9314 56756 9324
rect 56700 8932 56756 8942
rect 56588 8930 56756 8932
rect 56588 8878 56702 8930
rect 56754 8878 56756 8930
rect 56588 8876 56756 8878
rect 56140 8708 56196 8718
rect 56140 8258 56196 8652
rect 56140 8206 56142 8258
rect 56194 8206 56196 8258
rect 56140 8194 56196 8206
rect 56252 8372 56308 8382
rect 55692 7362 55748 7374
rect 55692 7310 55694 7362
rect 55746 7310 55748 7362
rect 55692 7252 55748 7310
rect 55692 7186 55748 7196
rect 55580 6804 55636 6814
rect 55580 6130 55636 6748
rect 56252 6802 56308 8316
rect 56588 8372 56644 8382
rect 56588 8278 56644 8316
rect 56588 7700 56644 7710
rect 56588 7606 56644 7644
rect 56700 7364 56756 8876
rect 57148 8370 57204 11454
rect 57260 11618 57316 12796
rect 57372 12786 57428 12796
rect 57372 12404 57428 12414
rect 57372 12310 57428 12348
rect 57708 12404 57764 13020
rect 57820 12982 57876 13020
rect 57932 12852 57988 13692
rect 57932 12786 57988 12796
rect 57820 12404 57876 12414
rect 57708 12402 57876 12404
rect 57708 12350 57822 12402
rect 57874 12350 57876 12402
rect 57708 12348 57876 12350
rect 57260 11566 57262 11618
rect 57314 11566 57316 11618
rect 57260 10276 57316 11566
rect 57372 11508 57428 11518
rect 57372 11284 57428 11452
rect 57596 11508 57652 11518
rect 57596 11414 57652 11452
rect 57372 10834 57428 11228
rect 57372 10782 57374 10834
rect 57426 10782 57428 10834
rect 57372 10500 57428 10782
rect 57372 10434 57428 10444
rect 57484 11396 57540 11406
rect 57260 10220 57428 10276
rect 57260 10052 57316 10062
rect 57260 9938 57316 9996
rect 57260 9886 57262 9938
rect 57314 9886 57316 9938
rect 57260 9874 57316 9886
rect 57148 8318 57150 8370
rect 57202 8318 57204 8370
rect 57148 8306 57204 8318
rect 57260 8820 57316 8830
rect 56700 7298 56756 7308
rect 56252 6750 56254 6802
rect 56306 6750 56308 6802
rect 56252 6738 56308 6750
rect 55804 6692 55860 6702
rect 55804 6598 55860 6636
rect 56700 6692 56756 6702
rect 56700 6598 56756 6636
rect 57260 6690 57316 8764
rect 57260 6638 57262 6690
rect 57314 6638 57316 6690
rect 57260 6626 57316 6638
rect 57372 7698 57428 10220
rect 57484 9940 57540 11340
rect 57596 9940 57652 9950
rect 57484 9938 57652 9940
rect 57484 9886 57598 9938
rect 57650 9886 57652 9938
rect 57484 9884 57652 9886
rect 57596 9874 57652 9884
rect 57708 9268 57764 12348
rect 57820 12338 57876 12348
rect 58044 11844 58100 20076
rect 57820 11788 58100 11844
rect 57820 9828 57876 11788
rect 58044 11618 58100 11630
rect 58044 11566 58046 11618
rect 58098 11566 58100 11618
rect 57932 11506 57988 11518
rect 57932 11454 57934 11506
rect 57986 11454 57988 11506
rect 57932 10834 57988 11454
rect 58044 11506 58100 11566
rect 58044 11454 58046 11506
rect 58098 11454 58100 11506
rect 58044 11442 58100 11454
rect 57932 10782 57934 10834
rect 57986 10782 57988 10834
rect 57932 10770 57988 10782
rect 58044 9940 58100 9950
rect 57820 9772 57988 9828
rect 57596 9212 57764 9268
rect 57484 9154 57540 9166
rect 57484 9102 57486 9154
rect 57538 9102 57540 9154
rect 57484 8708 57540 9102
rect 57484 8642 57540 8652
rect 57596 8260 57652 9212
rect 57708 9042 57764 9054
rect 57708 8990 57710 9042
rect 57762 8990 57764 9042
rect 57708 8596 57764 8990
rect 57708 8530 57764 8540
rect 57372 7646 57374 7698
rect 57426 7646 57428 7698
rect 57372 6692 57428 7646
rect 57484 8204 57652 8260
rect 57820 8482 57876 8494
rect 57820 8430 57822 8482
rect 57874 8430 57876 8482
rect 57484 7700 57540 8204
rect 57596 8036 57652 8046
rect 57596 7942 57652 7980
rect 57484 7634 57540 7644
rect 57820 7588 57876 8430
rect 57708 7532 57876 7588
rect 57428 6636 57540 6692
rect 57372 6626 57428 6636
rect 55580 6078 55582 6130
rect 55634 6078 55636 6130
rect 55580 6066 55636 6078
rect 56476 6132 56532 6142
rect 56476 6038 56532 6076
rect 57484 6130 57540 6636
rect 57596 6468 57652 6478
rect 57596 6374 57652 6412
rect 57484 6078 57486 6130
rect 57538 6078 57540 6130
rect 57484 6066 57540 6078
rect 55916 5796 55972 5806
rect 55916 5702 55972 5740
rect 57148 5684 57204 5694
rect 56700 5236 56756 5246
rect 56700 5142 56756 5180
rect 57148 5236 57204 5628
rect 57708 5572 57764 7532
rect 57820 7364 57876 7374
rect 57820 7270 57876 7308
rect 57932 6692 57988 9772
rect 58044 8482 58100 9884
rect 58044 8430 58046 8482
rect 58098 8430 58100 8482
rect 58044 8418 58100 8430
rect 58044 8034 58100 8046
rect 58044 7982 58046 8034
rect 58098 7982 58100 8034
rect 58044 6916 58100 7982
rect 58044 6850 58100 6860
rect 58044 6692 58100 6702
rect 57932 6690 58100 6692
rect 57932 6638 58046 6690
rect 58098 6638 58100 6690
rect 57932 6636 58100 6638
rect 58044 6626 58100 6636
rect 57820 6468 57876 6478
rect 57820 6130 57876 6412
rect 57820 6078 57822 6130
rect 57874 6078 57876 6130
rect 57820 6066 57876 6078
rect 57708 5516 57876 5572
rect 57596 5236 57652 5246
rect 57148 5234 57652 5236
rect 57148 5182 57150 5234
rect 57202 5182 57598 5234
rect 57650 5182 57652 5234
rect 57148 5180 57652 5182
rect 57148 5170 57204 5180
rect 57596 5170 57652 5180
rect 56252 5012 56308 5022
rect 55916 4898 55972 4910
rect 55916 4846 55918 4898
rect 55970 4846 55972 4898
rect 55916 3554 55972 4846
rect 56140 4452 56196 4462
rect 56140 4338 56196 4396
rect 56140 4286 56142 4338
rect 56194 4286 56196 4338
rect 56140 4274 56196 4286
rect 55916 3502 55918 3554
rect 55970 3502 55972 3554
rect 55916 3490 55972 3502
rect 56252 2884 56308 4956
rect 57484 4452 57540 4462
rect 57484 4358 57540 4396
rect 57708 4338 57764 4350
rect 57708 4286 57710 4338
rect 57762 4286 57764 4338
rect 56588 4226 56644 4238
rect 56588 4174 56590 4226
rect 56642 4174 56644 4226
rect 56588 4116 56644 4174
rect 56588 4050 56644 4060
rect 56700 4228 56756 4238
rect 56700 3668 56756 4172
rect 57484 4004 57540 4014
rect 57036 3668 57092 3678
rect 56700 3666 57092 3668
rect 56700 3614 56702 3666
rect 56754 3614 57038 3666
rect 57090 3614 57092 3666
rect 56700 3612 57092 3614
rect 56700 3602 56756 3612
rect 57036 3602 57092 3612
rect 57148 3668 57204 3678
rect 56252 2818 56308 2828
rect 55468 1586 55524 1596
rect 53900 1474 53956 1484
rect 57148 800 57204 3612
rect 57484 3666 57540 3948
rect 57484 3614 57486 3666
rect 57538 3614 57540 3666
rect 57484 3602 57540 3614
rect 57708 3332 57764 4286
rect 57708 3266 57764 3276
rect 57820 2660 57876 5516
rect 58044 4900 58100 4910
rect 58044 4806 58100 4844
rect 57932 3780 57988 3790
rect 57932 3666 57988 3724
rect 57932 3614 57934 3666
rect 57986 3614 57988 3666
rect 57932 3602 57988 3614
rect 58156 3388 58212 36316
rect 58268 34804 58324 34814
rect 58268 21028 58324 34748
rect 58268 20962 58324 20972
rect 58268 16772 58324 16782
rect 58268 16212 58324 16716
rect 58268 11618 58324 16156
rect 58380 14308 58436 41580
rect 58492 31444 58548 41692
rect 58604 38500 58660 45500
rect 58604 38434 58660 38444
rect 58716 41860 58772 41870
rect 58716 37604 58772 41804
rect 58716 33236 58772 37548
rect 58716 33170 58772 33180
rect 58492 31378 58548 31388
rect 58716 32564 58772 32574
rect 58492 27972 58548 27982
rect 58492 16772 58548 27916
rect 58604 25284 58660 25294
rect 58604 25190 58660 25228
rect 58492 16706 58548 16716
rect 58604 21028 58660 21038
rect 58380 14242 58436 14252
rect 58492 16548 58548 16558
rect 58268 11566 58270 11618
rect 58322 11566 58324 11618
rect 58268 11554 58324 11566
rect 58380 12852 58436 12862
rect 58380 5684 58436 12796
rect 58492 12404 58548 16492
rect 58492 12338 58548 12348
rect 58380 5618 58436 5628
rect 58604 5012 58660 20972
rect 58716 20132 58772 32508
rect 58828 29540 58884 45612
rect 58940 42532 58996 42542
rect 58940 34692 58996 42476
rect 58940 34626 58996 34636
rect 58828 29474 58884 29484
rect 59500 29540 59556 29550
rect 59164 29428 59220 29438
rect 59052 28756 59108 28766
rect 58940 25956 58996 25966
rect 58716 20066 58772 20076
rect 58828 23044 58884 23054
rect 58828 18900 58884 22988
rect 58716 18228 58772 18238
rect 58716 10836 58772 18172
rect 58828 16548 58884 18844
rect 58828 16482 58884 16492
rect 58716 10770 58772 10780
rect 58828 14868 58884 14878
rect 58828 8036 58884 14812
rect 58940 11508 58996 25900
rect 59052 22036 59108 28700
rect 59052 21970 59108 21980
rect 59164 20804 59220 29372
rect 59052 20748 59220 20804
rect 59276 23716 59332 23726
rect 59052 20468 59108 20748
rect 59052 13076 59108 20412
rect 59052 13010 59108 13020
rect 59164 19012 59220 19022
rect 58940 11442 58996 11452
rect 59164 9940 59220 18956
rect 59276 14868 59332 23660
rect 59276 14802 59332 14812
rect 59500 13524 59556 29484
rect 59500 13458 59556 13468
rect 59612 25282 59668 25294
rect 59612 25230 59614 25282
rect 59666 25230 59668 25282
rect 59164 9874 59220 9884
rect 58828 7970 58884 7980
rect 59612 7924 59668 25230
rect 59612 7858 59668 7868
rect 58604 4946 58660 4956
rect 58156 3332 58324 3388
rect 58268 3266 58324 3276
rect 57820 2594 57876 2604
rect 34636 700 35140 756
rect 40320 200 40432 800
rect 45696 200 45808 800
rect 51744 200 51856 800
rect 57120 200 57232 800
<< via2 >>
rect 1932 57148 1988 57204
rect 4172 56252 4228 56308
rect 4732 56306 4788 56308
rect 4732 56254 4734 56306
rect 4734 56254 4786 56306
rect 4786 56254 4788 56306
rect 4732 56252 4788 56254
rect 4476 55690 4532 55692
rect 4476 55638 4478 55690
rect 4478 55638 4530 55690
rect 4530 55638 4532 55690
rect 4476 55636 4532 55638
rect 4580 55690 4636 55692
rect 4580 55638 4582 55690
rect 4582 55638 4634 55690
rect 4634 55638 4636 55690
rect 4580 55636 4636 55638
rect 4684 55690 4740 55692
rect 4684 55638 4686 55690
rect 4686 55638 4738 55690
rect 4738 55638 4740 55690
rect 4684 55636 4740 55638
rect 3052 55020 3108 55076
rect 3500 55074 3556 55076
rect 3500 55022 3502 55074
rect 3502 55022 3554 55074
rect 3554 55022 3556 55074
rect 3500 55020 3556 55022
rect 4060 55020 4116 55076
rect 2716 53618 2772 53620
rect 2716 53566 2718 53618
rect 2718 53566 2770 53618
rect 2770 53566 2772 53618
rect 2716 53564 2772 53566
rect 3164 53618 3220 53620
rect 3164 53566 3166 53618
rect 3166 53566 3218 53618
rect 3218 53566 3220 53618
rect 3164 53564 3220 53566
rect 1932 51772 1988 51828
rect 3276 49868 3332 49924
rect 1148 48076 1204 48132
rect 1036 41020 1092 41076
rect 1932 45778 1988 45780
rect 1932 45726 1934 45778
rect 1934 45726 1986 45778
rect 1986 45726 1988 45778
rect 1932 45724 1988 45726
rect 1260 27132 1316 27188
rect 1260 16156 1316 16212
rect 1260 15148 1316 15204
rect 1932 39676 1988 39732
rect 3388 46060 3444 46116
rect 3164 45612 3220 45668
rect 2716 45218 2772 45220
rect 2716 45166 2718 45218
rect 2718 45166 2770 45218
rect 2770 45166 2772 45218
rect 2716 45164 2772 45166
rect 2828 43538 2884 43540
rect 2828 43486 2830 43538
rect 2830 43486 2882 43538
rect 2882 43486 2884 43538
rect 2828 43484 2884 43486
rect 3500 45836 3556 45892
rect 3276 45164 3332 45220
rect 2940 41244 2996 41300
rect 2604 41186 2660 41188
rect 2604 41134 2606 41186
rect 2606 41134 2658 41186
rect 2658 41134 2660 41186
rect 2604 41132 2660 41134
rect 3164 42252 3220 42308
rect 3052 41074 3108 41076
rect 3052 41022 3054 41074
rect 3054 41022 3106 41074
rect 3106 41022 3108 41074
rect 3052 41020 3108 41022
rect 3276 41132 3332 41188
rect 3500 41020 3556 41076
rect 3164 40572 3220 40628
rect 2940 35756 2996 35812
rect 2268 34860 2324 34916
rect 2828 34914 2884 34916
rect 2828 34862 2830 34914
rect 2830 34862 2882 34914
rect 2882 34862 2884 34914
rect 2828 34860 2884 34862
rect 1932 34300 1988 34356
rect 1596 32508 1652 32564
rect 2492 32396 2548 32452
rect 2380 31554 2436 31556
rect 2380 31502 2382 31554
rect 2382 31502 2434 31554
rect 2434 31502 2436 31554
rect 2380 31500 2436 31502
rect 2268 31388 2324 31444
rect 2828 31554 2884 31556
rect 2828 31502 2830 31554
rect 2830 31502 2882 31554
rect 2882 31502 2884 31554
rect 2828 31500 2884 31502
rect 1932 28252 1988 28308
rect 1596 21644 1652 21700
rect 1708 27692 1764 27748
rect 1820 26236 1876 26292
rect 1820 25564 1876 25620
rect 1932 25506 1988 25508
rect 1932 25454 1934 25506
rect 1934 25454 1986 25506
rect 1986 25454 1988 25506
rect 1932 25452 1988 25454
rect 2156 29650 2212 29652
rect 2156 29598 2158 29650
rect 2158 29598 2210 29650
rect 2210 29598 2212 29650
rect 2156 29596 2212 29598
rect 2380 28028 2436 28084
rect 2268 26908 2324 26964
rect 2156 26850 2212 26852
rect 2156 26798 2158 26850
rect 2158 26798 2210 26850
rect 2210 26798 2212 26850
rect 2156 26796 2212 26798
rect 2156 26178 2212 26180
rect 2156 26126 2158 26178
rect 2158 26126 2210 26178
rect 2210 26126 2212 26178
rect 2156 26124 2212 26126
rect 2268 25618 2324 25620
rect 2268 25566 2270 25618
rect 2270 25566 2322 25618
rect 2322 25566 2324 25618
rect 2268 25564 2324 25566
rect 2716 28028 2772 28084
rect 2604 27074 2660 27076
rect 2604 27022 2606 27074
rect 2606 27022 2658 27074
rect 2658 27022 2660 27074
rect 2604 27020 2660 27022
rect 2716 26684 2772 26740
rect 3836 42700 3892 42756
rect 3724 42588 3780 42644
rect 3948 41692 4004 41748
rect 3724 41298 3780 41300
rect 3724 41246 3726 41298
rect 3726 41246 3778 41298
rect 3778 41246 3780 41298
rect 3724 41244 3780 41246
rect 3724 41074 3780 41076
rect 3724 41022 3726 41074
rect 3726 41022 3778 41074
rect 3778 41022 3780 41074
rect 3724 41020 3780 41022
rect 4476 54122 4532 54124
rect 4476 54070 4478 54122
rect 4478 54070 4530 54122
rect 4530 54070 4532 54122
rect 4476 54068 4532 54070
rect 4580 54122 4636 54124
rect 4580 54070 4582 54122
rect 4582 54070 4634 54122
rect 4634 54070 4636 54122
rect 4580 54068 4636 54070
rect 4684 54122 4740 54124
rect 4684 54070 4686 54122
rect 4686 54070 4738 54122
rect 4738 54070 4740 54122
rect 4684 54068 4740 54070
rect 4476 52554 4532 52556
rect 4476 52502 4478 52554
rect 4478 52502 4530 52554
rect 4530 52502 4532 52554
rect 4476 52500 4532 52502
rect 4580 52554 4636 52556
rect 4580 52502 4582 52554
rect 4582 52502 4634 52554
rect 4634 52502 4636 52554
rect 4580 52500 4636 52502
rect 4684 52554 4740 52556
rect 4684 52502 4686 52554
rect 4686 52502 4738 52554
rect 4738 52502 4740 52554
rect 4684 52500 4740 52502
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 19836 56474 19892 56476
rect 19836 56422 19838 56474
rect 19838 56422 19890 56474
rect 19890 56422 19892 56474
rect 19836 56420 19892 56422
rect 19940 56474 19996 56476
rect 19940 56422 19942 56474
rect 19942 56422 19994 56474
rect 19994 56422 19996 56474
rect 19940 56420 19996 56422
rect 20044 56474 20100 56476
rect 20044 56422 20046 56474
rect 20046 56422 20098 56474
rect 20098 56422 20100 56474
rect 20044 56420 20100 56422
rect 29932 56140 29988 56196
rect 14140 56028 14196 56084
rect 10108 55916 10164 55972
rect 9548 49532 9604 49588
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 8764 48188 8820 48244
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 7756 47628 7812 47684
rect 7196 47404 7252 47460
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 5852 46284 5908 46340
rect 6412 46284 6468 46340
rect 5628 45666 5684 45668
rect 5628 45614 5630 45666
rect 5630 45614 5682 45666
rect 5682 45614 5684 45666
rect 5628 45612 5684 45614
rect 5740 45276 5796 45332
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 5068 44098 5124 44100
rect 5068 44046 5070 44098
rect 5070 44046 5122 44098
rect 5122 44046 5124 44098
rect 5068 44044 5124 44046
rect 5404 43484 5460 43540
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4956 42978 5012 42980
rect 4956 42926 4958 42978
rect 4958 42926 5010 42978
rect 5010 42926 5012 42978
rect 4956 42924 5012 42926
rect 5964 44098 6020 44100
rect 5964 44046 5966 44098
rect 5966 44046 6018 44098
rect 6018 44046 6020 44098
rect 5964 44044 6020 44046
rect 6748 44098 6804 44100
rect 6748 44046 6750 44098
rect 6750 44046 6802 44098
rect 6802 44046 6804 44098
rect 6748 44044 6804 44046
rect 4844 42642 4900 42644
rect 4844 42590 4846 42642
rect 4846 42590 4898 42642
rect 4898 42590 4900 42642
rect 4844 42588 4900 42590
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 5964 41970 6020 41972
rect 5964 41918 5966 41970
rect 5966 41918 6018 41970
rect 6018 41918 6020 41970
rect 5964 41916 6020 41918
rect 5740 41804 5796 41860
rect 5516 41692 5572 41748
rect 4956 40796 5012 40852
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4060 39788 4116 39844
rect 5404 40290 5460 40292
rect 5404 40238 5406 40290
rect 5406 40238 5458 40290
rect 5458 40238 5460 40290
rect 5404 40236 5460 40238
rect 3724 39058 3780 39060
rect 3724 39006 3726 39058
rect 3726 39006 3778 39058
rect 3778 39006 3780 39058
rect 3724 39004 3780 39006
rect 3948 38780 4004 38836
rect 4284 38780 4340 38836
rect 4396 39618 4452 39620
rect 4396 39566 4398 39618
rect 4398 39566 4450 39618
rect 4450 39566 4452 39618
rect 4396 39564 4452 39566
rect 4732 39004 4788 39060
rect 4620 38834 4676 38836
rect 4620 38782 4622 38834
rect 4622 38782 4674 38834
rect 4674 38782 4676 38834
rect 4620 38780 4676 38782
rect 4396 38668 4452 38724
rect 3612 38050 3668 38052
rect 3612 37998 3614 38050
rect 3614 37998 3666 38050
rect 3666 37998 3668 38050
rect 3612 37996 3668 37998
rect 3500 34914 3556 34916
rect 3500 34862 3502 34914
rect 3502 34862 3554 34914
rect 3554 34862 3556 34914
rect 3500 34860 3556 34862
rect 3388 31724 3444 31780
rect 2492 26012 2548 26068
rect 2492 25228 2548 25284
rect 2604 25676 2660 25732
rect 2156 23996 2212 24052
rect 2492 24668 2548 24724
rect 2044 23660 2100 23716
rect 1820 23042 1876 23044
rect 1820 22990 1822 23042
rect 1822 22990 1874 23042
rect 1874 22990 1876 23042
rect 1820 22988 1876 22990
rect 1932 22876 1988 22932
rect 2268 23660 2324 23716
rect 2380 23772 2436 23828
rect 2156 23548 2212 23604
rect 2268 22876 2324 22932
rect 2268 21308 2324 21364
rect 2044 20748 2100 20804
rect 1708 20636 1764 20692
rect 1932 20076 1988 20132
rect 1932 18620 1988 18676
rect 1820 18172 1876 18228
rect 1596 17724 1652 17780
rect 1372 12908 1428 12964
rect 1484 13020 1540 13076
rect 1260 10780 1316 10836
rect 1148 6636 1204 6692
rect 1372 5292 1428 5348
rect 1036 4396 1092 4452
rect 2156 20188 2212 20244
rect 2380 19234 2436 19236
rect 2380 19182 2382 19234
rect 2382 19182 2434 19234
rect 2434 19182 2436 19234
rect 2380 19180 2436 19182
rect 1708 15148 1764 15204
rect 1708 14924 1764 14980
rect 2268 17836 2324 17892
rect 2940 25676 2996 25732
rect 2828 25394 2884 25396
rect 2828 25342 2830 25394
rect 2830 25342 2882 25394
rect 2882 25342 2884 25394
rect 2828 25340 2884 25342
rect 2716 25004 2772 25060
rect 2828 25116 2884 25172
rect 3948 38556 4004 38612
rect 3836 32562 3892 32564
rect 3836 32510 3838 32562
rect 3838 32510 3890 32562
rect 3890 32510 3892 32562
rect 3836 32508 3892 32510
rect 3500 31500 3556 31556
rect 4844 38556 4900 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4172 38220 4228 38276
rect 4732 38220 4788 38276
rect 4620 38050 4676 38052
rect 4620 37998 4622 38050
rect 4622 37998 4674 38050
rect 4674 37998 4676 38050
rect 4620 37996 4676 37998
rect 4284 37938 4340 37940
rect 4284 37886 4286 37938
rect 4286 37886 4338 37938
rect 4338 37886 4340 37938
rect 4284 37884 4340 37886
rect 4172 37660 4228 37716
rect 4060 34690 4116 34692
rect 4060 34638 4062 34690
rect 4062 34638 4114 34690
rect 4114 34638 4116 34690
rect 4060 34636 4116 34638
rect 4396 37772 4452 37828
rect 4508 37884 4564 37940
rect 5404 39004 5460 39060
rect 5740 41074 5796 41076
rect 5740 41022 5742 41074
rect 5742 41022 5794 41074
rect 5794 41022 5796 41074
rect 5740 41020 5796 41022
rect 5740 40684 5796 40740
rect 5852 40290 5908 40292
rect 5852 40238 5854 40290
rect 5854 40238 5906 40290
rect 5906 40238 5908 40290
rect 5852 40236 5908 40238
rect 6748 43372 6804 43428
rect 6972 43538 7028 43540
rect 6972 43486 6974 43538
rect 6974 43486 7026 43538
rect 7026 43486 7028 43538
rect 6972 43484 7028 43486
rect 6412 42978 6468 42980
rect 6412 42926 6414 42978
rect 6414 42926 6466 42978
rect 6466 42926 6468 42978
rect 6412 42924 6468 42926
rect 6300 42754 6356 42756
rect 6300 42702 6302 42754
rect 6302 42702 6354 42754
rect 6354 42702 6356 42754
rect 6300 42700 6356 42702
rect 7644 43426 7700 43428
rect 7644 43374 7646 43426
rect 7646 43374 7698 43426
rect 7698 43374 7700 43426
rect 7644 43372 7700 43374
rect 8988 47682 9044 47684
rect 8988 47630 8990 47682
rect 8990 47630 9042 47682
rect 9042 47630 9044 47682
rect 8988 47628 9044 47630
rect 8764 47404 8820 47460
rect 9324 47234 9380 47236
rect 9324 47182 9326 47234
rect 9326 47182 9378 47234
rect 9378 47182 9380 47234
rect 9324 47180 9380 47182
rect 9772 49196 9828 49252
rect 13916 55970 13972 55972
rect 13916 55918 13918 55970
rect 13918 55918 13970 55970
rect 13970 55918 13972 55970
rect 13916 55916 13972 55918
rect 14364 55916 14420 55972
rect 15148 56028 15204 56084
rect 13580 55020 13636 55076
rect 10108 49532 10164 49588
rect 9772 48242 9828 48244
rect 9772 48190 9774 48242
rect 9774 48190 9826 48242
rect 9826 48190 9828 48242
rect 9772 48188 9828 48190
rect 10332 48914 10388 48916
rect 10332 48862 10334 48914
rect 10334 48862 10386 48914
rect 10386 48862 10388 48914
rect 10332 48860 10388 48862
rect 13244 49532 13300 49588
rect 13468 49308 13524 49364
rect 10444 48354 10500 48356
rect 10444 48302 10446 48354
rect 10446 48302 10498 48354
rect 10498 48302 10500 48354
rect 10444 48300 10500 48302
rect 11452 48860 11508 48916
rect 9660 47180 9716 47236
rect 10220 47628 10276 47684
rect 12572 48972 12628 49028
rect 10332 47404 10388 47460
rect 9100 46284 9156 46340
rect 9100 45778 9156 45780
rect 9100 45726 9102 45778
rect 9102 45726 9154 45778
rect 9154 45726 9156 45778
rect 9100 45724 9156 45726
rect 7868 44322 7924 44324
rect 7868 44270 7870 44322
rect 7870 44270 7922 44322
rect 7922 44270 7924 44322
rect 7868 44268 7924 44270
rect 8428 45330 8484 45332
rect 8428 45278 8430 45330
rect 8430 45278 8482 45330
rect 8482 45278 8484 45330
rect 8428 45276 8484 45278
rect 9772 45276 9828 45332
rect 9660 45164 9716 45220
rect 8540 44322 8596 44324
rect 8540 44270 8542 44322
rect 8542 44270 8594 44322
rect 8594 44270 8596 44322
rect 8540 44268 8596 44270
rect 8764 44268 8820 44324
rect 8092 43596 8148 43652
rect 7084 42924 7140 42980
rect 7980 43372 8036 43428
rect 6860 42700 6916 42756
rect 6748 41804 6804 41860
rect 6300 41074 6356 41076
rect 6300 41022 6302 41074
rect 6302 41022 6354 41074
rect 6354 41022 6356 41074
rect 6300 41020 6356 41022
rect 6300 40684 6356 40740
rect 6972 41916 7028 41972
rect 6860 41020 6916 41076
rect 6748 40684 6804 40740
rect 6524 40460 6580 40516
rect 5964 39618 6020 39620
rect 5964 39566 5966 39618
rect 5966 39566 6018 39618
rect 6018 39566 6020 39618
rect 5964 39564 6020 39566
rect 7756 42530 7812 42532
rect 7756 42478 7758 42530
rect 7758 42478 7810 42530
rect 7810 42478 7812 42530
rect 7756 42476 7812 42478
rect 7084 41692 7140 41748
rect 7420 42364 7476 42420
rect 6972 40460 7028 40516
rect 7308 40348 7364 40404
rect 8092 43036 8148 43092
rect 8092 42476 8148 42532
rect 8988 44156 9044 44212
rect 9324 44210 9380 44212
rect 9324 44158 9326 44210
rect 9326 44158 9378 44210
rect 9378 44158 9380 44210
rect 9324 44156 9380 44158
rect 8428 43372 8484 43428
rect 8204 42364 8260 42420
rect 8316 43148 8372 43204
rect 7532 40684 7588 40740
rect 7644 40514 7700 40516
rect 7644 40462 7646 40514
rect 7646 40462 7698 40514
rect 7698 40462 7700 40514
rect 7644 40460 7700 40462
rect 5180 38610 5236 38612
rect 5180 38558 5182 38610
rect 5182 38558 5234 38610
rect 5234 38558 5236 38610
rect 5180 38556 5236 38558
rect 4956 38108 5012 38164
rect 5628 38162 5684 38164
rect 5628 38110 5630 38162
rect 5630 38110 5682 38162
rect 5682 38110 5684 38162
rect 5628 38108 5684 38110
rect 5852 38556 5908 38612
rect 4956 37772 5012 37828
rect 4620 37100 4676 37156
rect 5180 37100 5236 37156
rect 5628 37154 5684 37156
rect 5628 37102 5630 37154
rect 5630 37102 5682 37154
rect 5682 37102 5684 37154
rect 5628 37100 5684 37102
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4844 35138 4900 35140
rect 4844 35086 4846 35138
rect 4846 35086 4898 35138
rect 4898 35086 4900 35138
rect 4844 35084 4900 35086
rect 4956 34972 5012 35028
rect 4732 34690 4788 34692
rect 4732 34638 4734 34690
rect 4734 34638 4786 34690
rect 4786 34638 4788 34690
rect 4732 34636 4788 34638
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4508 33404 4564 33460
rect 5068 33404 5124 33460
rect 4284 32450 4340 32452
rect 4284 32398 4286 32450
rect 4286 32398 4338 32450
rect 4338 32398 4340 32450
rect 4284 32396 4340 32398
rect 5180 32396 5236 32452
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 5068 32060 5124 32116
rect 4844 31948 4900 32004
rect 4172 31666 4228 31668
rect 4172 31614 4174 31666
rect 4174 31614 4226 31666
rect 4226 31614 4228 31666
rect 4172 31612 4228 31614
rect 3948 31276 4004 31332
rect 3836 31164 3892 31220
rect 4620 31218 4676 31220
rect 4620 31166 4622 31218
rect 4622 31166 4674 31218
rect 4674 31166 4676 31218
rect 4620 31164 4676 31166
rect 5068 31388 5124 31444
rect 6412 38780 6468 38836
rect 6636 38668 6692 38724
rect 5964 37938 6020 37940
rect 5964 37886 5966 37938
rect 5966 37886 6018 37938
rect 6018 37886 6020 37938
rect 5964 37884 6020 37886
rect 6188 37826 6244 37828
rect 6188 37774 6190 37826
rect 6190 37774 6242 37826
rect 6242 37774 6244 37826
rect 6188 37772 6244 37774
rect 7532 40012 7588 40068
rect 6748 38556 6804 38612
rect 6300 37154 6356 37156
rect 6300 37102 6302 37154
rect 6302 37102 6354 37154
rect 6354 37102 6356 37154
rect 6300 37100 6356 37102
rect 6636 36876 6692 36932
rect 6300 36204 6356 36260
rect 6188 35026 6244 35028
rect 6188 34974 6190 35026
rect 6190 34974 6242 35026
rect 6242 34974 6244 35026
rect 6188 34972 6244 34974
rect 6972 36876 7028 36932
rect 6972 36258 7028 36260
rect 6972 36206 6974 36258
rect 6974 36206 7026 36258
rect 7026 36206 7028 36258
rect 6972 36204 7028 36206
rect 7196 37212 7252 37268
rect 7308 36876 7364 36932
rect 7196 35980 7252 36036
rect 6300 34914 6356 34916
rect 6300 34862 6302 34914
rect 6302 34862 6354 34914
rect 6354 34862 6356 34914
rect 6300 34860 6356 34862
rect 5852 33628 5908 33684
rect 6636 34300 6692 34356
rect 7308 35644 7364 35700
rect 6972 34354 7028 34356
rect 6972 34302 6974 34354
rect 6974 34302 7026 34354
rect 7026 34302 7028 34354
rect 6972 34300 7028 34302
rect 7196 35026 7252 35028
rect 7196 34974 7198 35026
rect 7198 34974 7250 35026
rect 7250 34974 7252 35026
rect 7196 34972 7252 34974
rect 6076 33964 6132 34020
rect 5740 32956 5796 33012
rect 5404 32396 5460 32452
rect 5628 32338 5684 32340
rect 5628 32286 5630 32338
rect 5630 32286 5682 32338
rect 5682 32286 5684 32338
rect 5628 32284 5684 32286
rect 7196 34188 7252 34244
rect 6300 33516 6356 33572
rect 5852 32396 5908 32452
rect 7308 33852 7364 33908
rect 7308 33404 7364 33460
rect 6524 32620 6580 32676
rect 6748 33346 6804 33348
rect 6748 33294 6750 33346
rect 6750 33294 6802 33346
rect 6802 33294 6804 33346
rect 6748 33292 6804 33294
rect 6300 32284 6356 32340
rect 5740 32060 5796 32116
rect 6188 32060 6244 32116
rect 5292 31948 5348 32004
rect 6076 31948 6132 32004
rect 5740 31554 5796 31556
rect 5740 31502 5742 31554
rect 5742 31502 5794 31554
rect 5794 31502 5796 31554
rect 5740 31500 5796 31502
rect 7196 33122 7252 33124
rect 7196 33070 7198 33122
rect 7198 33070 7250 33122
rect 7250 33070 7252 33122
rect 7196 33068 7252 33070
rect 6748 31948 6804 32004
rect 4172 30716 4228 30772
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 3724 30098 3780 30100
rect 3724 30046 3726 30098
rect 3726 30046 3778 30098
rect 3778 30046 3780 30098
rect 3724 30044 3780 30046
rect 3164 27970 3220 27972
rect 3164 27918 3166 27970
rect 3166 27918 3218 27970
rect 3218 27918 3220 27970
rect 3164 27916 3220 27918
rect 3836 29932 3892 29988
rect 3388 29596 3444 29652
rect 3164 27132 3220 27188
rect 3724 28812 3780 28868
rect 3724 28028 3780 28084
rect 3612 27580 3668 27636
rect 3500 27132 3556 27188
rect 3948 28252 4004 28308
rect 3948 27858 4004 27860
rect 3948 27806 3950 27858
rect 3950 27806 4002 27858
rect 4002 27806 4004 27858
rect 3948 27804 4004 27806
rect 3836 27132 3892 27188
rect 3612 26908 3668 26964
rect 3500 26572 3556 26628
rect 3836 26514 3892 26516
rect 3836 26462 3838 26514
rect 3838 26462 3890 26514
rect 3890 26462 3892 26514
rect 3836 26460 3892 26462
rect 3276 25282 3332 25284
rect 3276 25230 3278 25282
rect 3278 25230 3330 25282
rect 3330 25230 3332 25282
rect 3276 25228 3332 25230
rect 3052 24220 3108 24276
rect 3164 24162 3220 24164
rect 3164 24110 3166 24162
rect 3166 24110 3218 24162
rect 3218 24110 3220 24162
rect 3164 24108 3220 24110
rect 2940 23660 2996 23716
rect 2828 22370 2884 22372
rect 2828 22318 2830 22370
rect 2830 22318 2882 22370
rect 2882 22318 2884 22370
rect 2828 22316 2884 22318
rect 2828 21698 2884 21700
rect 2828 21646 2830 21698
rect 2830 21646 2882 21698
rect 2882 21646 2884 21698
rect 2828 21644 2884 21646
rect 2604 20076 2660 20132
rect 2716 21532 2772 21588
rect 2604 19740 2660 19796
rect 3052 22204 3108 22260
rect 3164 23884 3220 23940
rect 3052 20636 3108 20692
rect 3164 21644 3220 21700
rect 3052 20300 3108 20356
rect 2940 19292 2996 19348
rect 2828 18732 2884 18788
rect 2044 16828 2100 16884
rect 1932 15372 1988 15428
rect 1932 15036 1988 15092
rect 2492 16716 2548 16772
rect 2604 16268 2660 16324
rect 3052 18284 3108 18340
rect 3052 17778 3108 17780
rect 3052 17726 3054 17778
rect 3054 17726 3106 17778
rect 3106 17726 3108 17778
rect 3052 17724 3108 17726
rect 2044 14924 2100 14980
rect 2716 15708 2772 15764
rect 2604 15596 2660 15652
rect 2716 15260 2772 15316
rect 3052 17164 3108 17220
rect 3388 24498 3444 24500
rect 3388 24446 3390 24498
rect 3390 24446 3442 24498
rect 3442 24446 3444 24498
rect 3388 24444 3444 24446
rect 3276 21532 3332 21588
rect 3612 24892 3668 24948
rect 3612 24220 3668 24276
rect 3276 20578 3332 20580
rect 3276 20526 3278 20578
rect 3278 20526 3330 20578
rect 3330 20526 3332 20578
rect 3276 20524 3332 20526
rect 3500 23714 3556 23716
rect 3500 23662 3502 23714
rect 3502 23662 3554 23714
rect 3554 23662 3556 23714
rect 3500 23660 3556 23662
rect 3500 23100 3556 23156
rect 3724 24108 3780 24164
rect 3612 22540 3668 22596
rect 4172 29260 4228 29316
rect 4172 25282 4228 25284
rect 4172 25230 4174 25282
rect 4174 25230 4226 25282
rect 4226 25230 4228 25282
rect 4172 25228 4228 25230
rect 5068 29986 5124 29988
rect 5068 29934 5070 29986
rect 5070 29934 5122 29986
rect 5122 29934 5124 29986
rect 5068 29932 5124 29934
rect 4620 29596 4676 29652
rect 4844 29538 4900 29540
rect 4844 29486 4846 29538
rect 4846 29486 4898 29538
rect 4898 29486 4900 29538
rect 4844 29484 4900 29486
rect 4396 29314 4452 29316
rect 4396 29262 4398 29314
rect 4398 29262 4450 29314
rect 4450 29262 4452 29314
rect 4396 29260 4452 29262
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 5068 29036 5124 29092
rect 4844 28028 4900 28084
rect 4396 27746 4452 27748
rect 4396 27694 4398 27746
rect 4398 27694 4450 27746
rect 4450 27694 4452 27746
rect 4396 27692 4452 27694
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4396 26962 4452 26964
rect 4396 26910 4398 26962
rect 4398 26910 4450 26962
rect 4450 26910 4452 26962
rect 4396 26908 4452 26910
rect 5292 30380 5348 30436
rect 5740 30380 5796 30436
rect 8204 41074 8260 41076
rect 8204 41022 8206 41074
rect 8206 41022 8258 41074
rect 8258 41022 8260 41074
rect 8204 41020 8260 41022
rect 7980 40962 8036 40964
rect 7980 40910 7982 40962
rect 7982 40910 8034 40962
rect 8034 40910 8036 40962
rect 7980 40908 8036 40910
rect 8204 40684 8260 40740
rect 8092 40460 8148 40516
rect 7868 40290 7924 40292
rect 7868 40238 7870 40290
rect 7870 40238 7922 40290
rect 7922 40238 7924 40290
rect 7868 40236 7924 40238
rect 7980 40124 8036 40180
rect 7756 39730 7812 39732
rect 7756 39678 7758 39730
rect 7758 39678 7810 39730
rect 7810 39678 7812 39730
rect 7756 39676 7812 39678
rect 7868 38556 7924 38612
rect 7868 37436 7924 37492
rect 7756 35586 7812 35588
rect 7756 35534 7758 35586
rect 7758 35534 7810 35586
rect 7810 35534 7812 35586
rect 7756 35532 7812 35534
rect 8540 41186 8596 41188
rect 8540 41134 8542 41186
rect 8542 41134 8594 41186
rect 8594 41134 8596 41186
rect 8540 41132 8596 41134
rect 8764 40460 8820 40516
rect 8316 40012 8372 40068
rect 8428 40236 8484 40292
rect 8092 39452 8148 39508
rect 8428 39842 8484 39844
rect 8428 39790 8430 39842
rect 8430 39790 8482 39842
rect 8482 39790 8484 39842
rect 8428 39788 8484 39790
rect 8092 38668 8148 38724
rect 8652 39676 8708 39732
rect 8540 39340 8596 39396
rect 8428 36764 8484 36820
rect 7980 34242 8036 34244
rect 7980 34190 7982 34242
rect 7982 34190 8034 34242
rect 8034 34190 8036 34242
rect 7980 34188 8036 34190
rect 7756 33964 7812 34020
rect 7868 33516 7924 33572
rect 6860 31612 6916 31668
rect 6188 30434 6244 30436
rect 6188 30382 6190 30434
rect 6190 30382 6242 30434
rect 6242 30382 6244 30434
rect 6188 30380 6244 30382
rect 6636 30380 6692 30436
rect 6972 30828 7028 30884
rect 5964 30322 6020 30324
rect 5964 30270 5966 30322
rect 5966 30270 6018 30322
rect 6018 30270 6020 30322
rect 5964 30268 6020 30270
rect 6748 30268 6804 30324
rect 6636 30044 6692 30100
rect 5628 29932 5684 29988
rect 5516 29820 5572 29876
rect 5628 29484 5684 29540
rect 5964 29932 6020 29988
rect 5180 28028 5236 28084
rect 4956 27746 5012 27748
rect 4956 27694 4958 27746
rect 4958 27694 5010 27746
rect 5010 27694 5012 27746
rect 4956 27692 5012 27694
rect 5180 27468 5236 27524
rect 4956 27356 5012 27412
rect 4956 27186 5012 27188
rect 4956 27134 4958 27186
rect 4958 27134 5010 27186
rect 5010 27134 5012 27186
rect 4956 27132 5012 27134
rect 4844 26684 4900 26740
rect 4396 26572 4452 26628
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4284 24892 4340 24948
rect 4396 25564 4452 25620
rect 4172 24780 4228 24836
rect 3948 23324 4004 23380
rect 4060 23154 4116 23156
rect 4060 23102 4062 23154
rect 4062 23102 4114 23154
rect 4114 23102 4116 23154
rect 4060 23100 4116 23102
rect 3724 22482 3780 22484
rect 3724 22430 3726 22482
rect 3726 22430 3778 22482
rect 3778 22430 3780 22482
rect 3724 22428 3780 22430
rect 3948 22316 4004 22372
rect 3836 22258 3892 22260
rect 3836 22206 3838 22258
rect 3838 22206 3890 22258
rect 3890 22206 3892 22258
rect 3836 22204 3892 22206
rect 3500 21474 3556 21476
rect 3500 21422 3502 21474
rect 3502 21422 3554 21474
rect 3554 21422 3556 21474
rect 3500 21420 3556 21422
rect 3388 20412 3444 20468
rect 3388 20018 3444 20020
rect 3388 19966 3390 20018
rect 3390 19966 3442 20018
rect 3442 19966 3444 20018
rect 3388 19964 3444 19966
rect 3276 19122 3332 19124
rect 3276 19070 3278 19122
rect 3278 19070 3330 19122
rect 3330 19070 3332 19122
rect 3276 19068 3332 19070
rect 3724 19404 3780 19460
rect 3612 19234 3668 19236
rect 3612 19182 3614 19234
rect 3614 19182 3666 19234
rect 3666 19182 3668 19234
rect 3612 19180 3668 19182
rect 3612 18844 3668 18900
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 5404 26402 5460 26404
rect 5404 26350 5406 26402
rect 5406 26350 5458 26402
rect 5458 26350 5460 26402
rect 5404 26348 5460 26350
rect 5180 25788 5236 25844
rect 4732 25564 4788 25620
rect 4956 25618 5012 25620
rect 4956 25566 4958 25618
rect 4958 25566 5010 25618
rect 5010 25566 5012 25618
rect 4956 25564 5012 25566
rect 4844 24668 4900 24724
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23884 4340 23940
rect 4844 23938 4900 23940
rect 4844 23886 4846 23938
rect 4846 23886 4898 23938
rect 4898 23886 4900 23938
rect 4844 23884 4900 23886
rect 4508 23324 4564 23380
rect 4396 23212 4452 23268
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 21868 4228 21924
rect 3948 19180 4004 19236
rect 3500 18450 3556 18452
rect 3500 18398 3502 18450
rect 3502 18398 3554 18450
rect 3554 18398 3556 18450
rect 3500 18396 3556 18398
rect 4172 20300 4228 20356
rect 4060 19122 4116 19124
rect 4060 19070 4062 19122
rect 4062 19070 4114 19122
rect 4114 19070 4116 19122
rect 4060 19068 4116 19070
rect 5068 25228 5124 25284
rect 5068 24892 5124 24948
rect 5292 25228 5348 25284
rect 5068 23660 5124 23716
rect 5516 24668 5572 24724
rect 4956 22764 5012 22820
rect 4956 22370 5012 22372
rect 4956 22318 4958 22370
rect 4958 22318 5010 22370
rect 5010 22318 5012 22370
rect 4956 22316 5012 22318
rect 4508 21586 4564 21588
rect 4508 21534 4510 21586
rect 4510 21534 4562 21586
rect 4562 21534 4564 21586
rect 4508 21532 4564 21534
rect 4956 21420 5012 21476
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4396 20972 4452 21028
rect 4620 20690 4676 20692
rect 4620 20638 4622 20690
rect 4622 20638 4674 20690
rect 4674 20638 4676 20690
rect 4620 20636 4676 20638
rect 4956 20300 5012 20356
rect 4732 20076 4788 20132
rect 4172 17612 4228 17668
rect 4508 20018 4564 20020
rect 4508 19966 4510 20018
rect 4510 19966 4562 20018
rect 4562 19966 4564 20018
rect 4508 19964 4564 19966
rect 3500 17164 3556 17220
rect 3276 16940 3332 16996
rect 4956 20018 5012 20020
rect 4956 19966 4958 20018
rect 4958 19966 5010 20018
rect 5010 19966 5012 20018
rect 4956 19964 5012 19966
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4620 19010 4676 19012
rect 4620 18958 4622 19010
rect 4622 18958 4674 19010
rect 4674 18958 4676 19010
rect 4620 18956 4676 18958
rect 4956 19122 5012 19124
rect 4956 19070 4958 19122
rect 4958 19070 5010 19122
rect 5010 19070 5012 19122
rect 4956 19068 5012 19070
rect 4620 18450 4676 18452
rect 4620 18398 4622 18450
rect 4622 18398 4674 18450
rect 4674 18398 4676 18450
rect 4620 18396 4676 18398
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5068 17948 5124 18004
rect 4620 17442 4676 17444
rect 4620 17390 4622 17442
rect 4622 17390 4674 17442
rect 4674 17390 4676 17442
rect 4620 17388 4676 17390
rect 4284 17164 4340 17220
rect 2940 14588 2996 14644
rect 3052 15314 3108 15316
rect 3052 15262 3054 15314
rect 3054 15262 3106 15314
rect 3106 15262 3108 15314
rect 3052 15260 3108 15262
rect 2828 14476 2884 14532
rect 2492 14140 2548 14196
rect 2716 13970 2772 13972
rect 2716 13918 2718 13970
rect 2718 13918 2770 13970
rect 2770 13918 2772 13970
rect 2716 13916 2772 13918
rect 2380 13580 2436 13636
rect 2828 13468 2884 13524
rect 2940 14028 2996 14084
rect 1932 13132 1988 13188
rect 2380 12962 2436 12964
rect 2380 12910 2382 12962
rect 2382 12910 2434 12962
rect 2434 12910 2436 12962
rect 2380 12908 2436 12910
rect 1932 11452 1988 11508
rect 2268 11340 2324 11396
rect 1820 11282 1876 11284
rect 1820 11230 1822 11282
rect 1822 11230 1874 11282
rect 1874 11230 1876 11282
rect 1820 11228 1876 11230
rect 2156 10722 2212 10724
rect 2156 10670 2158 10722
rect 2158 10670 2210 10722
rect 2210 10670 2212 10722
rect 2156 10668 2212 10670
rect 1932 9154 1988 9156
rect 1932 9102 1934 9154
rect 1934 9102 1986 9154
rect 1986 9102 1988 9154
rect 1932 9100 1988 9102
rect 2044 7586 2100 7588
rect 2044 7534 2046 7586
rect 2046 7534 2098 7586
rect 2098 7534 2100 7586
rect 2044 7532 2100 7534
rect 1932 6860 1988 6916
rect 2380 9938 2436 9940
rect 2380 9886 2382 9938
rect 2382 9886 2434 9938
rect 2434 9886 2436 9938
rect 2380 9884 2436 9886
rect 2716 9436 2772 9492
rect 2828 9042 2884 9044
rect 2828 8990 2830 9042
rect 2830 8990 2882 9042
rect 2882 8990 2884 9042
rect 2828 8988 2884 8990
rect 2380 7868 2436 7924
rect 2492 7980 2548 8036
rect 2268 6860 2324 6916
rect 2604 6690 2660 6692
rect 2604 6638 2606 6690
rect 2606 6638 2658 6690
rect 2658 6638 2660 6690
rect 2604 6636 2660 6638
rect 2940 7698 2996 7700
rect 2940 7646 2942 7698
rect 2942 7646 2994 7698
rect 2994 7646 2996 7698
rect 2940 7644 2996 7646
rect 2716 6188 2772 6244
rect 1932 5404 1988 5460
rect 2156 5234 2212 5236
rect 2156 5182 2158 5234
rect 2158 5182 2210 5234
rect 2210 5182 2212 5234
rect 2156 5180 2212 5182
rect 2604 5122 2660 5124
rect 2604 5070 2606 5122
rect 2606 5070 2658 5122
rect 2658 5070 2660 5122
rect 2604 5068 2660 5070
rect 2716 4450 2772 4452
rect 2716 4398 2718 4450
rect 2718 4398 2770 4450
rect 2770 4398 2772 4450
rect 2716 4396 2772 4398
rect 1596 2716 1652 2772
rect 28 1820 84 1876
rect 2940 2940 2996 2996
rect 1932 1820 1988 1876
rect 4396 16828 4452 16884
rect 3612 16604 3668 16660
rect 3612 15820 3668 15876
rect 4060 16716 4116 16772
rect 3948 15538 4004 15540
rect 3948 15486 3950 15538
rect 3950 15486 4002 15538
rect 4002 15486 4004 15538
rect 3948 15484 4004 15486
rect 3836 15036 3892 15092
rect 4172 16098 4228 16100
rect 4172 16046 4174 16098
rect 4174 16046 4226 16098
rect 4226 16046 4228 16098
rect 4172 16044 4228 16046
rect 5852 29314 5908 29316
rect 5852 29262 5854 29314
rect 5854 29262 5906 29314
rect 5906 29262 5908 29314
rect 5852 29260 5908 29262
rect 6188 29372 6244 29428
rect 6076 29260 6132 29316
rect 6076 28418 6132 28420
rect 6076 28366 6078 28418
rect 6078 28366 6130 28418
rect 6130 28366 6132 28418
rect 6076 28364 6132 28366
rect 5852 27746 5908 27748
rect 5852 27694 5854 27746
rect 5854 27694 5906 27746
rect 5906 27694 5908 27746
rect 5852 27692 5908 27694
rect 6076 27132 6132 27188
rect 6524 29314 6580 29316
rect 6524 29262 6526 29314
rect 6526 29262 6578 29314
rect 6578 29262 6580 29314
rect 6524 29260 6580 29262
rect 6300 28252 6356 28308
rect 6524 28082 6580 28084
rect 6524 28030 6526 28082
rect 6526 28030 6578 28082
rect 6578 28030 6580 28082
rect 6524 28028 6580 28030
rect 7084 30044 7140 30100
rect 7084 29484 7140 29540
rect 6972 29426 7028 29428
rect 6972 29374 6974 29426
rect 6974 29374 7026 29426
rect 7026 29374 7028 29426
rect 6972 29372 7028 29374
rect 6300 27634 6356 27636
rect 6300 27582 6302 27634
rect 6302 27582 6354 27634
rect 6354 27582 6356 27634
rect 6300 27580 6356 27582
rect 6860 27804 6916 27860
rect 5740 26908 5796 26964
rect 6300 26460 6356 26516
rect 5740 26236 5796 26292
rect 5740 25282 5796 25284
rect 5740 25230 5742 25282
rect 5742 25230 5794 25282
rect 5794 25230 5796 25282
rect 5740 25228 5796 25230
rect 6076 25564 6132 25620
rect 6076 25004 6132 25060
rect 5964 24556 6020 24612
rect 6300 24556 6356 24612
rect 6412 25116 6468 25172
rect 5964 24332 6020 24388
rect 6188 24444 6244 24500
rect 6188 23772 6244 23828
rect 6300 24108 6356 24164
rect 6188 23548 6244 23604
rect 5852 22428 5908 22484
rect 6076 23324 6132 23380
rect 5852 22258 5908 22260
rect 5852 22206 5854 22258
rect 5854 22206 5906 22258
rect 5906 22206 5908 22258
rect 5852 22204 5908 22206
rect 5852 21868 5908 21924
rect 5404 20972 5460 21028
rect 4956 17164 5012 17220
rect 5404 20188 5460 20244
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4844 16492 4900 16548
rect 4620 16210 4676 16212
rect 4620 16158 4622 16210
rect 4622 16158 4674 16210
rect 4674 16158 4676 16210
rect 4620 16156 4676 16158
rect 4284 15932 4340 15988
rect 4172 15148 4228 15204
rect 4172 14924 4228 14980
rect 3612 14642 3668 14644
rect 3612 14590 3614 14642
rect 3614 14590 3666 14642
rect 3666 14590 3668 14642
rect 3612 14588 3668 14590
rect 3500 13916 3556 13972
rect 3836 14252 3892 14308
rect 3276 12908 3332 12964
rect 3612 12850 3668 12852
rect 3612 12798 3614 12850
rect 3614 12798 3666 12850
rect 3666 12798 3668 12850
rect 3612 12796 3668 12798
rect 3164 11452 3220 11508
rect 3388 11452 3444 11508
rect 3164 10722 3220 10724
rect 3164 10670 3166 10722
rect 3166 10670 3218 10722
rect 3218 10670 3220 10722
rect 3164 10668 3220 10670
rect 3164 10444 3220 10500
rect 3276 10332 3332 10388
rect 3164 9436 3220 9492
rect 3164 7532 3220 7588
rect 3164 6636 3220 6692
rect 3612 11004 3668 11060
rect 3388 7644 3444 7700
rect 3500 9884 3556 9940
rect 4172 13692 4228 13748
rect 3948 12460 4004 12516
rect 3724 9602 3780 9604
rect 3724 9550 3726 9602
rect 3726 9550 3778 9602
rect 3778 9550 3780 9602
rect 3724 9548 3780 9550
rect 3724 9324 3780 9380
rect 4060 11340 4116 11396
rect 4060 9938 4116 9940
rect 4060 9886 4062 9938
rect 4062 9886 4114 9938
rect 4114 9886 4116 9938
rect 4060 9884 4116 9886
rect 3948 9660 4004 9716
rect 3948 8988 4004 9044
rect 3612 7980 3668 8036
rect 3836 7362 3892 7364
rect 3836 7310 3838 7362
rect 3838 7310 3890 7362
rect 3890 7310 3892 7362
rect 3836 7308 3892 7310
rect 3836 6860 3892 6916
rect 3724 6300 3780 6356
rect 3500 5794 3556 5796
rect 3500 5742 3502 5794
rect 3502 5742 3554 5794
rect 3554 5742 3556 5794
rect 3500 5740 3556 5742
rect 4844 15484 4900 15540
rect 5180 16828 5236 16884
rect 4732 15372 4788 15428
rect 5068 16098 5124 16100
rect 5068 16046 5070 16098
rect 5070 16046 5122 16098
rect 5122 16046 5124 16098
rect 5068 16044 5124 16046
rect 5740 19906 5796 19908
rect 5740 19854 5742 19906
rect 5742 19854 5794 19906
rect 5794 19854 5796 19906
rect 5740 19852 5796 19854
rect 6860 26796 6916 26852
rect 6860 26460 6916 26516
rect 6748 26290 6804 26292
rect 6748 26238 6750 26290
rect 6750 26238 6802 26290
rect 6802 26238 6804 26290
rect 6748 26236 6804 26238
rect 6636 25564 6692 25620
rect 7532 31666 7588 31668
rect 7532 31614 7534 31666
rect 7534 31614 7586 31666
rect 7586 31614 7588 31666
rect 7532 31612 7588 31614
rect 7532 31052 7588 31108
rect 7532 30882 7588 30884
rect 7532 30830 7534 30882
rect 7534 30830 7586 30882
rect 7586 30830 7588 30882
rect 7532 30828 7588 30830
rect 7756 31388 7812 31444
rect 7420 30268 7476 30324
rect 7532 30604 7588 30660
rect 7644 29986 7700 29988
rect 7644 29934 7646 29986
rect 7646 29934 7698 29986
rect 7698 29934 7700 29986
rect 7644 29932 7700 29934
rect 7532 29538 7588 29540
rect 7532 29486 7534 29538
rect 7534 29486 7586 29538
rect 7586 29486 7588 29538
rect 7532 29484 7588 29486
rect 7196 29260 7252 29316
rect 7308 28700 7364 28756
rect 8652 38556 8708 38612
rect 8988 41916 9044 41972
rect 8988 41244 9044 41300
rect 8988 41020 9044 41076
rect 8988 38668 9044 38724
rect 8876 37996 8932 38052
rect 9100 37660 9156 37716
rect 8652 36876 8708 36932
rect 9772 42924 9828 42980
rect 9772 41970 9828 41972
rect 9772 41918 9774 41970
rect 9774 41918 9826 41970
rect 9826 41918 9828 41970
rect 9772 41916 9828 41918
rect 10332 47180 10388 47236
rect 10108 45106 10164 45108
rect 10108 45054 10110 45106
rect 10110 45054 10162 45106
rect 10162 45054 10164 45106
rect 10108 45052 10164 45054
rect 12460 48354 12516 48356
rect 12460 48302 12462 48354
rect 12462 48302 12514 48354
rect 12514 48302 12516 48354
rect 12460 48300 12516 48302
rect 12012 48242 12068 48244
rect 12012 48190 12014 48242
rect 12014 48190 12066 48242
rect 12066 48190 12068 48242
rect 12012 48188 12068 48190
rect 11788 47516 11844 47572
rect 12460 47516 12516 47572
rect 11676 47404 11732 47460
rect 12236 47458 12292 47460
rect 12236 47406 12238 47458
rect 12238 47406 12290 47458
rect 12290 47406 12292 47458
rect 12236 47404 12292 47406
rect 11788 47346 11844 47348
rect 11788 47294 11790 47346
rect 11790 47294 11842 47346
rect 11842 47294 11844 47346
rect 11788 47292 11844 47294
rect 10780 46172 10836 46228
rect 12796 49026 12852 49028
rect 12796 48974 12798 49026
rect 12798 48974 12850 49026
rect 12850 48974 12852 49026
rect 12796 48972 12852 48974
rect 12684 48914 12740 48916
rect 12684 48862 12686 48914
rect 12686 48862 12738 48914
rect 12738 48862 12740 48914
rect 12684 48860 12740 48862
rect 12908 48802 12964 48804
rect 12908 48750 12910 48802
rect 12910 48750 12962 48802
rect 12962 48750 12964 48802
rect 12908 48748 12964 48750
rect 13132 47964 13188 48020
rect 12684 47516 12740 47572
rect 13020 47292 13076 47348
rect 11116 45724 11172 45780
rect 10556 45052 10612 45108
rect 10668 44940 10724 44996
rect 10220 43538 10276 43540
rect 10220 43486 10222 43538
rect 10222 43486 10274 43538
rect 10274 43486 10276 43538
rect 10220 43484 10276 43486
rect 10556 43596 10612 43652
rect 10332 42700 10388 42756
rect 9996 41692 10052 41748
rect 9436 41186 9492 41188
rect 9436 41134 9438 41186
rect 9438 41134 9490 41186
rect 9490 41134 9492 41186
rect 9436 41132 9492 41134
rect 9884 41132 9940 41188
rect 9548 41074 9604 41076
rect 9548 41022 9550 41074
rect 9550 41022 9602 41074
rect 9602 41022 9604 41074
rect 9548 41020 9604 41022
rect 9660 40908 9716 40964
rect 11116 44210 11172 44212
rect 11116 44158 11118 44210
rect 11118 44158 11170 44210
rect 11170 44158 11172 44210
rect 11116 44156 11172 44158
rect 11116 43538 11172 43540
rect 11116 43486 11118 43538
rect 11118 43486 11170 43538
rect 11170 43486 11172 43538
rect 11116 43484 11172 43486
rect 11116 43036 11172 43092
rect 11004 42754 11060 42756
rect 11004 42702 11006 42754
rect 11006 42702 11058 42754
rect 11058 42702 11060 42754
rect 11004 42700 11060 42702
rect 10780 41858 10836 41860
rect 10780 41806 10782 41858
rect 10782 41806 10834 41858
rect 10834 41806 10836 41858
rect 10780 41804 10836 41806
rect 10220 41186 10276 41188
rect 10220 41134 10222 41186
rect 10222 41134 10274 41186
rect 10274 41134 10276 41186
rect 10220 41132 10276 41134
rect 9996 40796 10052 40852
rect 10220 40514 10276 40516
rect 10220 40462 10222 40514
rect 10222 40462 10274 40514
rect 10274 40462 10276 40514
rect 10220 40460 10276 40462
rect 9772 39788 9828 39844
rect 9548 36876 9604 36932
rect 9660 38050 9716 38052
rect 9660 37998 9662 38050
rect 9662 37998 9714 38050
rect 9714 37998 9716 38050
rect 9660 37996 9716 37998
rect 9324 36764 9380 36820
rect 9436 36204 9492 36260
rect 8652 35644 8708 35700
rect 8876 35084 8932 35140
rect 8428 34300 8484 34356
rect 8316 33458 8372 33460
rect 8316 33406 8318 33458
rect 8318 33406 8370 33458
rect 8370 33406 8372 33458
rect 8316 33404 8372 33406
rect 7980 33068 8036 33124
rect 8204 33122 8260 33124
rect 8204 33070 8206 33122
rect 8206 33070 8258 33122
rect 8258 33070 8260 33122
rect 8204 33068 8260 33070
rect 8540 33852 8596 33908
rect 8428 33068 8484 33124
rect 9324 35532 9380 35588
rect 9548 35980 9604 36036
rect 9100 35026 9156 35028
rect 9100 34974 9102 35026
rect 9102 34974 9154 35026
rect 9154 34974 9156 35026
rect 9100 34972 9156 34974
rect 8988 34300 9044 34356
rect 9100 34242 9156 34244
rect 9100 34190 9102 34242
rect 9102 34190 9154 34242
rect 9154 34190 9156 34242
rect 9100 34188 9156 34190
rect 8988 33740 9044 33796
rect 8764 32674 8820 32676
rect 8764 32622 8766 32674
rect 8766 32622 8818 32674
rect 8818 32622 8820 32674
rect 8764 32620 8820 32622
rect 8540 31836 8596 31892
rect 8428 31612 8484 31668
rect 9100 33516 9156 33572
rect 8316 31388 8372 31444
rect 8092 30994 8148 30996
rect 8092 30942 8094 30994
rect 8094 30942 8146 30994
rect 8146 30942 8148 30994
rect 8092 30940 8148 30942
rect 8092 30716 8148 30772
rect 7196 28530 7252 28532
rect 7196 28478 7198 28530
rect 7198 28478 7250 28530
rect 7250 28478 7252 28530
rect 7196 28476 7252 28478
rect 7196 27858 7252 27860
rect 7196 27806 7198 27858
rect 7198 27806 7250 27858
rect 7250 27806 7252 27858
rect 7196 27804 7252 27806
rect 7420 27858 7476 27860
rect 7420 27806 7422 27858
rect 7422 27806 7474 27858
rect 7474 27806 7476 27858
rect 7420 27804 7476 27806
rect 7420 27580 7476 27636
rect 7308 27074 7364 27076
rect 7308 27022 7310 27074
rect 7310 27022 7362 27074
rect 7362 27022 7364 27074
rect 7308 27020 7364 27022
rect 7196 26850 7252 26852
rect 7196 26798 7198 26850
rect 7198 26798 7250 26850
rect 7250 26798 7252 26850
rect 7196 26796 7252 26798
rect 7084 26684 7140 26740
rect 7196 26572 7252 26628
rect 7532 26460 7588 26516
rect 7308 25618 7364 25620
rect 7308 25566 7310 25618
rect 7310 25566 7362 25618
rect 7362 25566 7364 25618
rect 7308 25564 7364 25566
rect 7420 26124 7476 26180
rect 7420 25676 7476 25732
rect 7196 25340 7252 25396
rect 7532 25564 7588 25620
rect 7420 25340 7476 25396
rect 6748 25228 6804 25284
rect 7308 24780 7364 24836
rect 6972 24722 7028 24724
rect 6972 24670 6974 24722
rect 6974 24670 7026 24722
rect 7026 24670 7028 24722
rect 6972 24668 7028 24670
rect 7196 24668 7252 24724
rect 6300 22370 6356 22372
rect 6300 22318 6302 22370
rect 6302 22318 6354 22370
rect 6354 22318 6356 22370
rect 6300 22316 6356 22318
rect 6748 23938 6804 23940
rect 6748 23886 6750 23938
rect 6750 23886 6802 23938
rect 6802 23886 6804 23938
rect 6748 23884 6804 23886
rect 7868 27858 7924 27860
rect 7868 27806 7870 27858
rect 7870 27806 7922 27858
rect 7922 27806 7924 27858
rect 7868 27804 7924 27806
rect 8316 31106 8372 31108
rect 8316 31054 8318 31106
rect 8318 31054 8370 31106
rect 8370 31054 8372 31106
rect 8316 31052 8372 31054
rect 8428 30882 8484 30884
rect 8428 30830 8430 30882
rect 8430 30830 8482 30882
rect 8482 30830 8484 30882
rect 8428 30828 8484 30830
rect 8540 30604 8596 30660
rect 8652 30940 8708 30996
rect 9212 33346 9268 33348
rect 9212 33294 9214 33346
rect 9214 33294 9266 33346
rect 9266 33294 9268 33346
rect 9212 33292 9268 33294
rect 8876 30604 8932 30660
rect 8316 30322 8372 30324
rect 8316 30270 8318 30322
rect 8318 30270 8370 30322
rect 8370 30270 8372 30322
rect 8316 30268 8372 30270
rect 9100 30268 9156 30324
rect 7644 24780 7700 24836
rect 8428 29650 8484 29652
rect 8428 29598 8430 29650
rect 8430 29598 8482 29650
rect 8482 29598 8484 29650
rect 8428 29596 8484 29598
rect 7868 26572 7924 26628
rect 7980 26236 8036 26292
rect 8652 29708 8708 29764
rect 9100 28700 9156 28756
rect 8428 28588 8484 28644
rect 8652 28642 8708 28644
rect 8652 28590 8654 28642
rect 8654 28590 8706 28642
rect 8706 28590 8708 28642
rect 8652 28588 8708 28590
rect 9996 38722 10052 38724
rect 9996 38670 9998 38722
rect 9998 38670 10050 38722
rect 10050 38670 10052 38722
rect 9996 38668 10052 38670
rect 10668 41074 10724 41076
rect 10668 41022 10670 41074
rect 10670 41022 10722 41074
rect 10722 41022 10724 41074
rect 10668 41020 10724 41022
rect 10780 40908 10836 40964
rect 10668 39506 10724 39508
rect 10668 39454 10670 39506
rect 10670 39454 10722 39506
rect 10722 39454 10724 39506
rect 10668 39452 10724 39454
rect 10332 38668 10388 38724
rect 10220 38444 10276 38500
rect 10220 38220 10276 38276
rect 9884 37660 9940 37716
rect 10332 36764 10388 36820
rect 9772 36482 9828 36484
rect 9772 36430 9774 36482
rect 9774 36430 9826 36482
rect 9826 36430 9828 36482
rect 9772 36428 9828 36430
rect 10220 36258 10276 36260
rect 10220 36206 10222 36258
rect 10222 36206 10274 36258
rect 10274 36206 10276 36258
rect 10220 36204 10276 36206
rect 9996 35980 10052 36036
rect 9660 35756 9716 35812
rect 9884 35420 9940 35476
rect 9996 35084 10052 35140
rect 10556 38722 10612 38724
rect 10556 38670 10558 38722
rect 10558 38670 10610 38722
rect 10610 38670 10612 38722
rect 10556 38668 10612 38670
rect 10556 38108 10612 38164
rect 11116 40012 11172 40068
rect 11116 39394 11172 39396
rect 11116 39342 11118 39394
rect 11118 39342 11170 39394
rect 11170 39342 11172 39394
rect 11116 39340 11172 39342
rect 12012 45218 12068 45220
rect 12012 45166 12014 45218
rect 12014 45166 12066 45218
rect 12066 45166 12068 45218
rect 12012 45164 12068 45166
rect 11564 44994 11620 44996
rect 11564 44942 11566 44994
rect 11566 44942 11618 44994
rect 11618 44942 11620 44994
rect 11564 44940 11620 44942
rect 11452 44098 11508 44100
rect 11452 44046 11454 44098
rect 11454 44046 11506 44098
rect 11506 44046 11508 44098
rect 11452 44044 11508 44046
rect 11900 44044 11956 44100
rect 11788 43650 11844 43652
rect 11788 43598 11790 43650
rect 11790 43598 11842 43650
rect 11842 43598 11844 43650
rect 11788 43596 11844 43598
rect 12012 43484 12068 43540
rect 12124 43036 12180 43092
rect 11452 42700 11508 42756
rect 11340 40460 11396 40516
rect 12684 45276 12740 45332
rect 12572 45218 12628 45220
rect 12572 45166 12574 45218
rect 12574 45166 12626 45218
rect 12626 45166 12628 45218
rect 12572 45164 12628 45166
rect 19836 54906 19892 54908
rect 19836 54854 19838 54906
rect 19838 54854 19890 54906
rect 19890 54854 19892 54906
rect 19836 54852 19892 54854
rect 19940 54906 19996 54908
rect 19940 54854 19942 54906
rect 19942 54854 19994 54906
rect 19994 54854 19996 54906
rect 19940 54852 19996 54854
rect 20044 54906 20100 54908
rect 20044 54854 20046 54906
rect 20046 54854 20098 54906
rect 20098 54854 20100 54906
rect 20044 54852 20100 54854
rect 19836 53338 19892 53340
rect 19836 53286 19838 53338
rect 19838 53286 19890 53338
rect 19890 53286 19892 53338
rect 19836 53284 19892 53286
rect 19940 53338 19996 53340
rect 19940 53286 19942 53338
rect 19942 53286 19994 53338
rect 19994 53286 19996 53338
rect 19940 53284 19996 53286
rect 20044 53338 20100 53340
rect 20044 53286 20046 53338
rect 20046 53286 20098 53338
rect 20098 53286 20100 53338
rect 20044 53284 20100 53286
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 13692 49532 13748 49588
rect 13916 49308 13972 49364
rect 13692 49084 13748 49140
rect 17612 49644 17668 49700
rect 14476 49308 14532 49364
rect 13804 48802 13860 48804
rect 13804 48750 13806 48802
rect 13806 48750 13858 48802
rect 13858 48750 13860 48802
rect 13804 48748 13860 48750
rect 13804 48242 13860 48244
rect 13804 48190 13806 48242
rect 13806 48190 13858 48242
rect 13858 48190 13860 48242
rect 13804 48188 13860 48190
rect 14028 47964 14084 48020
rect 13804 47458 13860 47460
rect 13804 47406 13806 47458
rect 13806 47406 13858 47458
rect 13858 47406 13860 47458
rect 13804 47404 13860 47406
rect 14028 47458 14084 47460
rect 14028 47406 14030 47458
rect 14030 47406 14082 47458
rect 14082 47406 14084 47458
rect 14028 47404 14084 47406
rect 13916 47346 13972 47348
rect 13916 47294 13918 47346
rect 13918 47294 13970 47346
rect 13970 47294 13972 47346
rect 13916 47292 13972 47294
rect 14028 46674 14084 46676
rect 14028 46622 14030 46674
rect 14030 46622 14082 46674
rect 14082 46622 14084 46674
rect 14028 46620 14084 46622
rect 13132 45276 13188 45332
rect 13580 45330 13636 45332
rect 13580 45278 13582 45330
rect 13582 45278 13634 45330
rect 13634 45278 13636 45330
rect 13580 45276 13636 45278
rect 12796 44940 12852 44996
rect 13132 44156 13188 44212
rect 13580 43820 13636 43876
rect 12572 43538 12628 43540
rect 12572 43486 12574 43538
rect 12574 43486 12626 43538
rect 12626 43486 12628 43538
rect 12572 43484 12628 43486
rect 12684 42924 12740 42980
rect 12348 42700 12404 42756
rect 11564 40124 11620 40180
rect 12348 40178 12404 40180
rect 12348 40126 12350 40178
rect 12350 40126 12402 40178
rect 12402 40126 12404 40178
rect 12348 40124 12404 40126
rect 12124 40012 12180 40068
rect 12572 39900 12628 39956
rect 11340 38668 11396 38724
rect 10892 37996 10948 38052
rect 11116 37996 11172 38052
rect 11228 37938 11284 37940
rect 11228 37886 11230 37938
rect 11230 37886 11282 37938
rect 11282 37886 11284 37938
rect 11228 37884 11284 37886
rect 10892 37660 10948 37716
rect 11116 37548 11172 37604
rect 10220 35308 10276 35364
rect 9884 34412 9940 34468
rect 10668 36204 10724 36260
rect 11004 35308 11060 35364
rect 10668 34914 10724 34916
rect 10668 34862 10670 34914
rect 10670 34862 10722 34914
rect 10722 34862 10724 34914
rect 10668 34860 10724 34862
rect 11004 34354 11060 34356
rect 11004 34302 11006 34354
rect 11006 34302 11058 34354
rect 11058 34302 11060 34354
rect 11004 34300 11060 34302
rect 9660 34188 9716 34244
rect 9660 32956 9716 33012
rect 9772 32620 9828 32676
rect 9100 28364 9156 28420
rect 8764 27858 8820 27860
rect 8764 27806 8766 27858
rect 8766 27806 8818 27858
rect 8818 27806 8820 27858
rect 8764 27804 8820 27806
rect 9324 28252 9380 28308
rect 8428 27356 8484 27412
rect 8316 27298 8372 27300
rect 8316 27246 8318 27298
rect 8318 27246 8370 27298
rect 8370 27246 8372 27298
rect 8316 27244 8372 27246
rect 8316 27020 8372 27076
rect 12124 38892 12180 38948
rect 11676 38444 11732 38500
rect 11676 37436 11732 37492
rect 12460 38946 12516 38948
rect 12460 38894 12462 38946
rect 12462 38894 12514 38946
rect 12514 38894 12516 38946
rect 12460 38892 12516 38894
rect 14028 45276 14084 45332
rect 14028 44994 14084 44996
rect 14028 44942 14030 44994
rect 14030 44942 14082 44994
rect 14082 44942 14084 44994
rect 14028 44940 14084 44942
rect 15820 49196 15876 49252
rect 17052 49196 17108 49252
rect 16044 49026 16100 49028
rect 16044 48974 16046 49026
rect 16046 48974 16098 49026
rect 16098 48974 16100 49026
rect 16044 48972 16100 48974
rect 16940 49026 16996 49028
rect 16940 48974 16942 49026
rect 16942 48974 16994 49026
rect 16994 48974 16996 49026
rect 16940 48972 16996 48974
rect 16268 48412 16324 48468
rect 14364 46898 14420 46900
rect 14364 46846 14366 46898
rect 14366 46846 14418 46898
rect 14418 46846 14420 46898
rect 14364 46844 14420 46846
rect 15932 48130 15988 48132
rect 15932 48078 15934 48130
rect 15934 48078 15986 48130
rect 15986 48078 15988 48130
rect 15932 48076 15988 48078
rect 17276 48300 17332 48356
rect 16604 48242 16660 48244
rect 16604 48190 16606 48242
rect 16606 48190 16658 48242
rect 16658 48190 16660 48242
rect 16604 48188 16660 48190
rect 15148 47404 15204 47460
rect 14924 47068 14980 47124
rect 15148 47068 15204 47124
rect 16268 46844 16324 46900
rect 14476 46620 14532 46676
rect 17052 47180 17108 47236
rect 16828 46898 16884 46900
rect 16828 46846 16830 46898
rect 16830 46846 16882 46898
rect 16882 46846 16884 46898
rect 16828 46844 16884 46846
rect 14700 45276 14756 45332
rect 14252 44940 14308 44996
rect 14588 45052 14644 45108
rect 14252 44322 14308 44324
rect 14252 44270 14254 44322
rect 14254 44270 14306 44322
rect 14306 44270 14308 44322
rect 14252 44268 14308 44270
rect 14364 43708 14420 43764
rect 13692 42924 13748 42980
rect 12796 42140 12852 42196
rect 12908 42812 12964 42868
rect 13804 42866 13860 42868
rect 13804 42814 13806 42866
rect 13806 42814 13858 42866
rect 13858 42814 13860 42866
rect 13804 42812 13860 42814
rect 13132 42028 13188 42084
rect 13692 42588 13748 42644
rect 13356 42140 13412 42196
rect 13020 40236 13076 40292
rect 12796 40178 12852 40180
rect 12796 40126 12798 40178
rect 12798 40126 12850 40178
rect 12850 40126 12852 40178
rect 12796 40124 12852 40126
rect 13020 39228 13076 39284
rect 13020 38834 13076 38836
rect 13020 38782 13022 38834
rect 13022 38782 13074 38834
rect 13074 38782 13076 38834
rect 13020 38780 13076 38782
rect 12348 37826 12404 37828
rect 12348 37774 12350 37826
rect 12350 37774 12402 37826
rect 12402 37774 12404 37826
rect 12348 37772 12404 37774
rect 12236 37660 12292 37716
rect 12012 37436 12068 37492
rect 11452 37378 11508 37380
rect 11452 37326 11454 37378
rect 11454 37326 11506 37378
rect 11506 37326 11508 37378
rect 11452 37324 11508 37326
rect 11564 36316 11620 36372
rect 11228 35810 11284 35812
rect 11228 35758 11230 35810
rect 11230 35758 11282 35810
rect 11282 35758 11284 35810
rect 11228 35756 11284 35758
rect 11340 35308 11396 35364
rect 11340 34914 11396 34916
rect 11340 34862 11342 34914
rect 11342 34862 11394 34914
rect 11394 34862 11396 34914
rect 11340 34860 11396 34862
rect 11228 34242 11284 34244
rect 11228 34190 11230 34242
rect 11230 34190 11282 34242
rect 11282 34190 11284 34242
rect 11228 34188 11284 34190
rect 11228 33964 11284 34020
rect 10108 33404 10164 33460
rect 9660 30716 9716 30772
rect 10108 32508 10164 32564
rect 10892 32450 10948 32452
rect 10892 32398 10894 32450
rect 10894 32398 10946 32450
rect 10946 32398 10948 32450
rect 10892 32396 10948 32398
rect 10220 31948 10276 32004
rect 10332 31890 10388 31892
rect 10332 31838 10334 31890
rect 10334 31838 10386 31890
rect 10386 31838 10388 31890
rect 10332 31836 10388 31838
rect 10668 31836 10724 31892
rect 10332 31612 10388 31668
rect 10108 31388 10164 31444
rect 9884 30828 9940 30884
rect 10220 30716 10276 30772
rect 9548 29986 9604 29988
rect 9548 29934 9550 29986
rect 9550 29934 9602 29986
rect 9602 29934 9604 29986
rect 9548 29932 9604 29934
rect 9548 29596 9604 29652
rect 9884 29708 9940 29764
rect 9436 27580 9492 27636
rect 9548 29148 9604 29204
rect 8428 26684 8484 26740
rect 8316 26460 8372 26516
rect 8540 26460 8596 26516
rect 8428 26290 8484 26292
rect 8428 26238 8430 26290
rect 8430 26238 8482 26290
rect 8482 26238 8484 26290
rect 8428 26236 8484 26238
rect 7980 25506 8036 25508
rect 7980 25454 7982 25506
rect 7982 25454 8034 25506
rect 8034 25454 8036 25506
rect 7980 25452 8036 25454
rect 7756 24668 7812 24724
rect 7868 25116 7924 25172
rect 7980 24162 8036 24164
rect 7980 24110 7982 24162
rect 7982 24110 8034 24162
rect 8034 24110 8036 24162
rect 7980 24108 8036 24110
rect 8204 23884 8260 23940
rect 6636 23100 6692 23156
rect 6748 23548 6804 23604
rect 6748 22428 6804 22484
rect 6860 23436 6916 23492
rect 6636 22370 6692 22372
rect 6636 22318 6638 22370
rect 6638 22318 6690 22370
rect 6690 22318 6692 22370
rect 6636 22316 6692 22318
rect 6748 22092 6804 22148
rect 6412 21644 6468 21700
rect 6300 20802 6356 20804
rect 6300 20750 6302 20802
rect 6302 20750 6354 20802
rect 6354 20750 6356 20802
rect 6300 20748 6356 20750
rect 6300 20524 6356 20580
rect 6076 19628 6132 19684
rect 5516 18508 5572 18564
rect 5180 15372 5236 15428
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4508 14530 4564 14532
rect 4508 14478 4510 14530
rect 4510 14478 4562 14530
rect 4562 14478 4564 14530
rect 4508 14476 4564 14478
rect 4508 13970 4564 13972
rect 4508 13918 4510 13970
rect 4510 13918 4562 13970
rect 4562 13918 4564 13970
rect 4508 13916 4564 13918
rect 4956 14924 5012 14980
rect 4956 14306 5012 14308
rect 4956 14254 4958 14306
rect 4958 14254 5010 14306
rect 5010 14254 5012 14306
rect 4956 14252 5012 14254
rect 4844 13468 4900 13524
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4620 13132 4676 13188
rect 4620 12908 4676 12964
rect 4396 12460 4452 12516
rect 5068 13804 5124 13860
rect 5516 17948 5572 18004
rect 5628 17500 5684 17556
rect 5740 16994 5796 16996
rect 5740 16942 5742 16994
rect 5742 16942 5794 16994
rect 5794 16942 5796 16994
rect 5740 16940 5796 16942
rect 5964 19010 6020 19012
rect 5964 18958 5966 19010
rect 5966 18958 6018 19010
rect 6018 18958 6020 19010
rect 5964 18956 6020 18958
rect 6188 18562 6244 18564
rect 6188 18510 6190 18562
rect 6190 18510 6242 18562
rect 6242 18510 6244 18562
rect 6188 18508 6244 18510
rect 6636 20802 6692 20804
rect 6636 20750 6638 20802
rect 6638 20750 6690 20802
rect 6690 20750 6692 20802
rect 6636 20748 6692 20750
rect 6748 20524 6804 20580
rect 7196 23436 7252 23492
rect 7196 22988 7252 23044
rect 7084 22428 7140 22484
rect 6972 22370 7028 22372
rect 6972 22318 6974 22370
rect 6974 22318 7026 22370
rect 7026 22318 7028 22370
rect 6972 22316 7028 22318
rect 6412 20188 6468 20244
rect 6972 21420 7028 21476
rect 6636 19852 6692 19908
rect 6524 19180 6580 19236
rect 5964 17442 6020 17444
rect 5964 17390 5966 17442
rect 5966 17390 6018 17442
rect 6018 17390 6020 17442
rect 5964 17388 6020 17390
rect 6636 17948 6692 18004
rect 5852 16716 5908 16772
rect 6412 17388 6468 17444
rect 5740 15986 5796 15988
rect 5740 15934 5742 15986
rect 5742 15934 5794 15986
rect 5794 15934 5796 15986
rect 5740 15932 5796 15934
rect 5404 15538 5460 15540
rect 5404 15486 5406 15538
rect 5406 15486 5458 15538
rect 5458 15486 5460 15538
rect 5404 15484 5460 15486
rect 5740 14364 5796 14420
rect 5292 13916 5348 13972
rect 5740 13916 5796 13972
rect 5180 13692 5236 13748
rect 5068 12572 5124 12628
rect 5068 12348 5124 12404
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 5292 13468 5348 13524
rect 5628 13244 5684 13300
rect 5292 12236 5348 12292
rect 5404 13132 5460 13188
rect 5068 11564 5124 11620
rect 4284 11340 4340 11396
rect 4956 11394 5012 11396
rect 4956 11342 4958 11394
rect 4958 11342 5010 11394
rect 5010 11342 5012 11394
rect 4956 11340 5012 11342
rect 4396 11116 4452 11172
rect 4284 10834 4340 10836
rect 4284 10782 4286 10834
rect 4286 10782 4338 10834
rect 4338 10782 4340 10834
rect 4284 10780 4340 10782
rect 4620 11004 4676 11060
rect 4508 10668 4564 10724
rect 4732 10332 4788 10388
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4620 9714 4676 9716
rect 4620 9662 4622 9714
rect 4622 9662 4674 9714
rect 4674 9662 4676 9714
rect 4620 9660 4676 9662
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4172 7196 4228 7252
rect 4396 7196 4452 7252
rect 4508 8428 4564 8484
rect 4956 9826 5012 9828
rect 4956 9774 4958 9826
rect 4958 9774 5010 9826
rect 5010 9774 5012 9826
rect 4956 9772 5012 9774
rect 5180 10556 5236 10612
rect 5068 8988 5124 9044
rect 4620 7532 4676 7588
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 5180 6748 5236 6804
rect 4508 6578 4564 6580
rect 4508 6526 4510 6578
rect 4510 6526 4562 6578
rect 4562 6526 4564 6578
rect 4508 6524 4564 6526
rect 4956 6412 5012 6468
rect 3948 6130 4004 6132
rect 3948 6078 3950 6130
rect 3950 6078 4002 6130
rect 4002 6078 4004 6130
rect 3948 6076 4004 6078
rect 3612 4450 3668 4452
rect 3612 4398 3614 4450
rect 3614 4398 3666 4450
rect 3666 4398 3668 4450
rect 3612 4396 3668 4398
rect 3836 3052 3892 3108
rect 4508 6130 4564 6132
rect 4508 6078 4510 6130
rect 4510 6078 4562 6130
rect 4562 6078 4564 6130
rect 4508 6076 4564 6078
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4508 5234 4564 5236
rect 4508 5182 4510 5234
rect 4510 5182 4562 5234
rect 4562 5182 4564 5234
rect 4508 5180 4564 5182
rect 4956 5234 5012 5236
rect 4956 5182 4958 5234
rect 4958 5182 5010 5234
rect 5010 5182 5012 5234
rect 4956 5180 5012 5182
rect 4956 4620 5012 4676
rect 4620 4562 4676 4564
rect 4620 4510 4622 4562
rect 4622 4510 4674 4562
rect 4674 4510 4676 4562
rect 4620 4508 4676 4510
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 5628 12460 5684 12516
rect 5516 10220 5572 10276
rect 5404 9660 5460 9716
rect 6412 16882 6468 16884
rect 6412 16830 6414 16882
rect 6414 16830 6466 16882
rect 6466 16830 6468 16882
rect 6412 16828 6468 16830
rect 6636 17164 6692 17220
rect 6636 15932 6692 15988
rect 6972 17612 7028 17668
rect 7196 21532 7252 21588
rect 7308 23100 7364 23156
rect 7644 23660 7700 23716
rect 7532 23548 7588 23604
rect 7532 23324 7588 23380
rect 7868 23548 7924 23604
rect 7420 22370 7476 22372
rect 7420 22318 7422 22370
rect 7422 22318 7474 22370
rect 7474 22318 7476 22370
rect 7420 22316 7476 22318
rect 7644 22146 7700 22148
rect 7644 22094 7646 22146
rect 7646 22094 7698 22146
rect 7698 22094 7700 22146
rect 7644 22092 7700 22094
rect 8092 21868 8148 21924
rect 7980 21810 8036 21812
rect 7980 21758 7982 21810
rect 7982 21758 8034 21810
rect 8034 21758 8036 21810
rect 7980 21756 8036 21758
rect 7868 21586 7924 21588
rect 7868 21534 7870 21586
rect 7870 21534 7922 21586
rect 7922 21534 7924 21586
rect 7868 21532 7924 21534
rect 7644 21474 7700 21476
rect 7644 21422 7646 21474
rect 7646 21422 7698 21474
rect 7698 21422 7700 21474
rect 7644 21420 7700 21422
rect 7980 21420 8036 21476
rect 7308 20188 7364 20244
rect 7196 20076 7252 20132
rect 7308 20018 7364 20020
rect 7308 19966 7310 20018
rect 7310 19966 7362 20018
rect 7362 19966 7364 20018
rect 7308 19964 7364 19966
rect 7532 20524 7588 20580
rect 8092 21308 8148 21364
rect 7980 20524 8036 20580
rect 7980 20188 8036 20244
rect 7756 19404 7812 19460
rect 7868 18562 7924 18564
rect 7868 18510 7870 18562
rect 7870 18510 7922 18562
rect 7922 18510 7924 18562
rect 7868 18508 7924 18510
rect 7084 17500 7140 17556
rect 6860 16492 6916 16548
rect 7308 16994 7364 16996
rect 7308 16942 7310 16994
rect 7310 16942 7362 16994
rect 7362 16942 7364 16994
rect 7308 16940 7364 16942
rect 7196 16882 7252 16884
rect 7196 16830 7198 16882
rect 7198 16830 7250 16882
rect 7250 16830 7252 16882
rect 7196 16828 7252 16830
rect 7532 18396 7588 18452
rect 7532 18060 7588 18116
rect 7644 17666 7700 17668
rect 7644 17614 7646 17666
rect 7646 17614 7698 17666
rect 7698 17614 7700 17666
rect 7644 17612 7700 17614
rect 7868 17500 7924 17556
rect 7420 16716 7476 16772
rect 7308 16492 7364 16548
rect 7084 16156 7140 16212
rect 7532 17052 7588 17108
rect 7420 15986 7476 15988
rect 7420 15934 7422 15986
rect 7422 15934 7474 15986
rect 7474 15934 7476 15986
rect 7420 15932 7476 15934
rect 6972 15372 7028 15428
rect 7196 15372 7252 15428
rect 6188 13858 6244 13860
rect 6188 13806 6190 13858
rect 6190 13806 6242 13858
rect 6242 13806 6244 13858
rect 6188 13804 6244 13806
rect 5964 13468 6020 13524
rect 5852 12796 5908 12852
rect 6188 12908 6244 12964
rect 5964 12124 6020 12180
rect 6860 15148 6916 15204
rect 7756 16658 7812 16660
rect 7756 16606 7758 16658
rect 7758 16606 7810 16658
rect 7810 16606 7812 16658
rect 7756 16604 7812 16606
rect 8092 20018 8148 20020
rect 8092 19966 8094 20018
rect 8094 19966 8146 20018
rect 8146 19966 8148 20018
rect 8092 19964 8148 19966
rect 8092 19292 8148 19348
rect 8092 19010 8148 19012
rect 8092 18958 8094 19010
rect 8094 18958 8146 19010
rect 8146 18958 8148 19010
rect 8092 18956 8148 18958
rect 8428 25340 8484 25396
rect 8428 24722 8484 24724
rect 8428 24670 8430 24722
rect 8430 24670 8482 24722
rect 8482 24670 8484 24722
rect 8428 24668 8484 24670
rect 8988 26066 9044 26068
rect 8988 26014 8990 26066
rect 8990 26014 9042 26066
rect 9042 26014 9044 26066
rect 8988 26012 9044 26014
rect 8652 25900 8708 25956
rect 9212 26460 9268 26516
rect 9324 26684 9380 26740
rect 9100 25228 9156 25284
rect 9324 25900 9380 25956
rect 9212 24668 9268 24724
rect 8540 24332 8596 24388
rect 9100 24332 9156 24388
rect 9100 24108 9156 24164
rect 8876 24050 8932 24052
rect 8876 23998 8878 24050
rect 8878 23998 8930 24050
rect 8930 23998 8932 24050
rect 8876 23996 8932 23998
rect 8540 23660 8596 23716
rect 8540 22540 8596 22596
rect 8428 22316 8484 22372
rect 9100 22764 9156 22820
rect 9436 24108 9492 24164
rect 8988 21980 9044 22036
rect 9212 21868 9268 21924
rect 8876 21532 8932 21588
rect 8428 19180 8484 19236
rect 8540 20524 8596 20580
rect 8428 18620 8484 18676
rect 8204 18060 8260 18116
rect 8204 17778 8260 17780
rect 8204 17726 8206 17778
rect 8206 17726 8258 17778
rect 8258 17726 8260 17778
rect 8204 17724 8260 17726
rect 8092 17500 8148 17556
rect 7644 15484 7700 15540
rect 7980 15932 8036 15988
rect 7644 15148 7700 15204
rect 6412 14418 6468 14420
rect 6412 14366 6414 14418
rect 6414 14366 6466 14418
rect 6466 14366 6468 14418
rect 6412 14364 6468 14366
rect 6412 12124 6468 12180
rect 6188 11116 6244 11172
rect 6300 10722 6356 10724
rect 6300 10670 6302 10722
rect 6302 10670 6354 10722
rect 6354 10670 6356 10722
rect 6300 10668 6356 10670
rect 6412 10610 6468 10612
rect 6412 10558 6414 10610
rect 6414 10558 6466 10610
rect 6466 10558 6468 10610
rect 6412 10556 6468 10558
rect 6412 10220 6468 10276
rect 5628 8876 5684 8932
rect 5516 8764 5572 8820
rect 5292 6130 5348 6132
rect 5292 6078 5294 6130
rect 5294 6078 5346 6130
rect 5346 6078 5348 6130
rect 5292 6076 5348 6078
rect 5404 7532 5460 7588
rect 5516 7474 5572 7476
rect 5516 7422 5518 7474
rect 5518 7422 5570 7474
rect 5570 7422 5572 7474
rect 5516 7420 5572 7422
rect 5740 6802 5796 6804
rect 5740 6750 5742 6802
rect 5742 6750 5794 6802
rect 5794 6750 5796 6802
rect 5740 6748 5796 6750
rect 5516 6524 5572 6580
rect 5740 6188 5796 6244
rect 6188 9826 6244 9828
rect 6188 9774 6190 9826
rect 6190 9774 6242 9826
rect 6242 9774 6244 9826
rect 6188 9772 6244 9774
rect 6076 7756 6132 7812
rect 6300 9436 6356 9492
rect 6748 15036 6804 15092
rect 7420 14588 7476 14644
rect 6860 14530 6916 14532
rect 6860 14478 6862 14530
rect 6862 14478 6914 14530
rect 6914 14478 6916 14530
rect 6860 14476 6916 14478
rect 7196 14476 7252 14532
rect 6860 14028 6916 14084
rect 6636 13020 6692 13076
rect 6524 9884 6580 9940
rect 6636 11340 6692 11396
rect 6524 9154 6580 9156
rect 6524 9102 6526 9154
rect 6526 9102 6578 9154
rect 6578 9102 6580 9154
rect 6524 9100 6580 9102
rect 6412 9042 6468 9044
rect 6412 8990 6414 9042
rect 6414 8990 6466 9042
rect 6466 8990 6468 9042
rect 6412 8988 6468 8990
rect 6748 10834 6804 10836
rect 6748 10782 6750 10834
rect 6750 10782 6802 10834
rect 6802 10782 6804 10834
rect 6748 10780 6804 10782
rect 6748 10444 6804 10500
rect 7644 14642 7700 14644
rect 7644 14590 7646 14642
rect 7646 14590 7698 14642
rect 7698 14590 7700 14642
rect 7644 14588 7700 14590
rect 7532 14418 7588 14420
rect 7532 14366 7534 14418
rect 7534 14366 7586 14418
rect 7586 14366 7588 14418
rect 7532 14364 7588 14366
rect 7420 14028 7476 14084
rect 7756 13916 7812 13972
rect 7756 13746 7812 13748
rect 7756 13694 7758 13746
rect 7758 13694 7810 13746
rect 7810 13694 7812 13746
rect 7756 13692 7812 13694
rect 7196 12962 7252 12964
rect 7196 12910 7198 12962
rect 7198 12910 7250 12962
rect 7250 12910 7252 12962
rect 7196 12908 7252 12910
rect 6972 12178 7028 12180
rect 6972 12126 6974 12178
rect 6974 12126 7026 12178
rect 7026 12126 7028 12178
rect 6972 12124 7028 12126
rect 7868 13244 7924 13300
rect 7756 13074 7812 13076
rect 7756 13022 7758 13074
rect 7758 13022 7810 13074
rect 7810 13022 7812 13074
rect 7756 13020 7812 13022
rect 8092 15314 8148 15316
rect 8092 15262 8094 15314
rect 8094 15262 8146 15314
rect 8146 15262 8148 15314
rect 8092 15260 8148 15262
rect 8092 13916 8148 13972
rect 8092 12684 8148 12740
rect 7308 12460 7364 12516
rect 7420 11394 7476 11396
rect 7420 11342 7422 11394
rect 7422 11342 7474 11394
rect 7474 11342 7476 11394
rect 7420 11340 7476 11342
rect 7084 10556 7140 10612
rect 7644 12178 7700 12180
rect 7644 12126 7646 12178
rect 7646 12126 7698 12178
rect 7698 12126 7700 12178
rect 7644 12124 7700 12126
rect 7196 9324 7252 9380
rect 7308 9772 7364 9828
rect 6748 7644 6804 7700
rect 6636 7586 6692 7588
rect 6636 7534 6638 7586
rect 6638 7534 6690 7586
rect 6690 7534 6692 7586
rect 6636 7532 6692 7534
rect 6748 7420 6804 7476
rect 6076 6860 6132 6916
rect 6412 5964 6468 6020
rect 6524 6300 6580 6356
rect 5404 4620 5460 4676
rect 5516 5180 5572 5236
rect 7084 7474 7140 7476
rect 7084 7422 7086 7474
rect 7086 7422 7138 7474
rect 7138 7422 7140 7474
rect 7084 7420 7140 7422
rect 7084 6690 7140 6692
rect 7084 6638 7086 6690
rect 7086 6638 7138 6690
rect 7138 6638 7140 6690
rect 7084 6636 7140 6638
rect 6636 5964 6692 6020
rect 5852 5234 5908 5236
rect 5852 5182 5854 5234
rect 5854 5182 5906 5234
rect 5906 5182 5908 5234
rect 5852 5180 5908 5182
rect 6188 5292 6244 5348
rect 5964 5068 6020 5124
rect 5068 4284 5124 4340
rect 4620 3442 4676 3444
rect 4620 3390 4622 3442
rect 4622 3390 4674 3442
rect 4674 3390 4676 3442
rect 4620 3388 4676 3390
rect 5404 3388 5460 3444
rect 4172 2492 4228 2548
rect 3052 1260 3108 1316
rect 5852 3442 5908 3444
rect 5852 3390 5854 3442
rect 5854 3390 5906 3442
rect 5906 3390 5908 3442
rect 5852 3388 5908 3390
rect 7084 5740 7140 5796
rect 6860 5122 6916 5124
rect 6860 5070 6862 5122
rect 6862 5070 6914 5122
rect 6914 5070 6916 5122
rect 6860 5068 6916 5070
rect 7084 4844 7140 4900
rect 6636 4508 6692 4564
rect 7420 8988 7476 9044
rect 7980 11452 8036 11508
rect 8092 12012 8148 12068
rect 8316 17164 8372 17220
rect 8316 16940 8372 16996
rect 8652 19180 8708 19236
rect 8764 18508 8820 18564
rect 8540 18450 8596 18452
rect 8540 18398 8542 18450
rect 8542 18398 8594 18450
rect 8594 18398 8596 18450
rect 8540 18396 8596 18398
rect 8652 18284 8708 18340
rect 8652 17836 8708 17892
rect 8540 17554 8596 17556
rect 8540 17502 8542 17554
rect 8542 17502 8594 17554
rect 8594 17502 8596 17554
rect 8540 17500 8596 17502
rect 8428 16380 8484 16436
rect 8428 16210 8484 16212
rect 8428 16158 8430 16210
rect 8430 16158 8482 16210
rect 8482 16158 8484 16210
rect 8428 16156 8484 16158
rect 8988 20802 9044 20804
rect 8988 20750 8990 20802
rect 8990 20750 9042 20802
rect 9042 20750 9044 20802
rect 8988 20748 9044 20750
rect 9100 20412 9156 20468
rect 8988 19516 9044 19572
rect 8988 19234 9044 19236
rect 8988 19182 8990 19234
rect 8990 19182 9042 19234
rect 9042 19182 9044 19234
rect 8988 19180 9044 19182
rect 8988 18732 9044 18788
rect 9100 18620 9156 18676
rect 9100 18396 9156 18452
rect 9212 18060 9268 18116
rect 9772 28252 9828 28308
rect 9660 27580 9716 27636
rect 9996 29148 10052 29204
rect 9996 28700 10052 28756
rect 10108 28364 10164 28420
rect 10220 28588 10276 28644
rect 10220 28082 10276 28084
rect 10220 28030 10222 28082
rect 10222 28030 10274 28082
rect 10274 28030 10276 28082
rect 10220 28028 10276 28030
rect 9884 27356 9940 27412
rect 10444 31554 10500 31556
rect 10444 31502 10446 31554
rect 10446 31502 10498 31554
rect 10498 31502 10500 31554
rect 10444 31500 10500 31502
rect 10556 30882 10612 30884
rect 10556 30830 10558 30882
rect 10558 30830 10610 30882
rect 10610 30830 10612 30882
rect 10556 30828 10612 30830
rect 10444 29820 10500 29876
rect 10780 31500 10836 31556
rect 10892 31218 10948 31220
rect 10892 31166 10894 31218
rect 10894 31166 10946 31218
rect 10946 31166 10948 31218
rect 10892 31164 10948 31166
rect 10892 30604 10948 30660
rect 11116 31052 11172 31108
rect 10780 30268 10836 30324
rect 10444 29426 10500 29428
rect 10444 29374 10446 29426
rect 10446 29374 10498 29426
rect 10498 29374 10500 29426
rect 10444 29372 10500 29374
rect 10444 29036 10500 29092
rect 10444 27804 10500 27860
rect 10332 26962 10388 26964
rect 10332 26910 10334 26962
rect 10334 26910 10386 26962
rect 10386 26910 10388 26962
rect 10332 26908 10388 26910
rect 9884 26012 9940 26068
rect 9996 25900 10052 25956
rect 10444 26572 10500 26628
rect 10892 29932 10948 29988
rect 10780 29202 10836 29204
rect 10780 29150 10782 29202
rect 10782 29150 10834 29202
rect 10834 29150 10836 29202
rect 10780 29148 10836 29150
rect 11116 30098 11172 30100
rect 11116 30046 11118 30098
rect 11118 30046 11170 30098
rect 11170 30046 11172 30098
rect 11116 30044 11172 30046
rect 11564 34860 11620 34916
rect 11452 30716 11508 30772
rect 11004 29484 11060 29540
rect 11004 29314 11060 29316
rect 11004 29262 11006 29314
rect 11006 29262 11058 29314
rect 11058 29262 11060 29314
rect 11004 29260 11060 29262
rect 10780 28140 10836 28196
rect 10668 28082 10724 28084
rect 10668 28030 10670 28082
rect 10670 28030 10722 28082
rect 10722 28030 10724 28082
rect 10668 28028 10724 28030
rect 10556 26236 10612 26292
rect 10780 26908 10836 26964
rect 9996 25394 10052 25396
rect 9996 25342 9998 25394
rect 9998 25342 10050 25394
rect 10050 25342 10052 25394
rect 9996 25340 10052 25342
rect 9772 25228 9828 25284
rect 9772 25004 9828 25060
rect 10108 25004 10164 25060
rect 9884 24834 9940 24836
rect 9884 24782 9886 24834
rect 9886 24782 9938 24834
rect 9938 24782 9940 24834
rect 9884 24780 9940 24782
rect 10108 24610 10164 24612
rect 10108 24558 10110 24610
rect 10110 24558 10162 24610
rect 10162 24558 10164 24610
rect 10108 24556 10164 24558
rect 9772 23884 9828 23940
rect 9996 23772 10052 23828
rect 9772 21868 9828 21924
rect 9548 17948 9604 18004
rect 10220 23660 10276 23716
rect 10220 22540 10276 22596
rect 10108 22092 10164 22148
rect 10444 25116 10500 25172
rect 10444 24722 10500 24724
rect 10444 24670 10446 24722
rect 10446 24670 10498 24722
rect 10498 24670 10500 24722
rect 10444 24668 10500 24670
rect 11228 29596 11284 29652
rect 11900 36428 11956 36484
rect 12460 37548 12516 37604
rect 11788 35810 11844 35812
rect 11788 35758 11790 35810
rect 11790 35758 11842 35810
rect 11842 35758 11844 35810
rect 11788 35756 11844 35758
rect 12908 37660 12964 37716
rect 12908 36988 12964 37044
rect 12908 36258 12964 36260
rect 12908 36206 12910 36258
rect 12910 36206 12962 36258
rect 12962 36206 12964 36258
rect 12908 36204 12964 36206
rect 14252 43372 14308 43428
rect 14252 43036 14308 43092
rect 14140 42642 14196 42644
rect 14140 42590 14142 42642
rect 14142 42590 14194 42642
rect 14194 42590 14196 42642
rect 14140 42588 14196 42590
rect 13916 42082 13972 42084
rect 13916 42030 13918 42082
rect 13918 42030 13970 42082
rect 13970 42030 13972 42082
rect 13916 42028 13972 42030
rect 13692 40236 13748 40292
rect 13804 40178 13860 40180
rect 13804 40126 13806 40178
rect 13806 40126 13858 40178
rect 13858 40126 13860 40178
rect 13804 40124 13860 40126
rect 13916 39900 13972 39956
rect 14140 40290 14196 40292
rect 14140 40238 14142 40290
rect 14142 40238 14194 40290
rect 14194 40238 14196 40290
rect 14140 40236 14196 40238
rect 14140 39900 14196 39956
rect 14028 39394 14084 39396
rect 14028 39342 14030 39394
rect 14030 39342 14082 39394
rect 14082 39342 14084 39394
rect 14028 39340 14084 39342
rect 13132 37212 13188 37268
rect 13244 36876 13300 36932
rect 13916 38722 13972 38724
rect 13916 38670 13918 38722
rect 13918 38670 13970 38722
rect 13970 38670 13972 38722
rect 13916 38668 13972 38670
rect 14028 38332 14084 38388
rect 13804 37378 13860 37380
rect 13804 37326 13806 37378
rect 13806 37326 13858 37378
rect 13858 37326 13860 37378
rect 13804 37324 13860 37326
rect 13356 36988 13412 37044
rect 13244 35586 13300 35588
rect 13244 35534 13246 35586
rect 13246 35534 13298 35586
rect 13298 35534 13300 35586
rect 13244 35532 13300 35534
rect 12012 34860 12068 34916
rect 12796 34860 12852 34916
rect 12012 34412 12068 34468
rect 11900 34188 11956 34244
rect 11676 32732 11732 32788
rect 11788 33628 11844 33684
rect 13244 34748 13300 34804
rect 12012 33628 12068 33684
rect 11900 33180 11956 33236
rect 12460 33234 12516 33236
rect 12460 33182 12462 33234
rect 12462 33182 12514 33234
rect 12514 33182 12516 33234
rect 12460 33180 12516 33182
rect 12348 33122 12404 33124
rect 12348 33070 12350 33122
rect 12350 33070 12402 33122
rect 12402 33070 12404 33122
rect 12348 33068 12404 33070
rect 12460 32562 12516 32564
rect 12460 32510 12462 32562
rect 12462 32510 12514 32562
rect 12514 32510 12516 32562
rect 12460 32508 12516 32510
rect 12348 31890 12404 31892
rect 12348 31838 12350 31890
rect 12350 31838 12402 31890
rect 12402 31838 12404 31890
rect 12348 31836 12404 31838
rect 12236 30994 12292 30996
rect 12236 30942 12238 30994
rect 12238 30942 12290 30994
rect 12290 30942 12292 30994
rect 12236 30940 12292 30942
rect 11788 30828 11844 30884
rect 11564 29596 11620 29652
rect 12012 30604 12068 30660
rect 11676 30044 11732 30100
rect 11900 29708 11956 29764
rect 11564 29426 11620 29428
rect 11564 29374 11566 29426
rect 11566 29374 11618 29426
rect 11618 29374 11620 29426
rect 11564 29372 11620 29374
rect 11340 28700 11396 28756
rect 11228 28642 11284 28644
rect 11228 28590 11230 28642
rect 11230 28590 11282 28642
rect 11282 28590 11284 28642
rect 11228 28588 11284 28590
rect 11676 28476 11732 28532
rect 11228 27244 11284 27300
rect 11116 26962 11172 26964
rect 11116 26910 11118 26962
rect 11118 26910 11170 26962
rect 11170 26910 11172 26962
rect 11116 26908 11172 26910
rect 11228 26684 11284 26740
rect 10892 26012 10948 26068
rect 10444 23714 10500 23716
rect 10444 23662 10446 23714
rect 10446 23662 10498 23714
rect 10498 23662 10500 23714
rect 10444 23660 10500 23662
rect 10556 23548 10612 23604
rect 10332 22316 10388 22372
rect 10444 22146 10500 22148
rect 10444 22094 10446 22146
rect 10446 22094 10498 22146
rect 10498 22094 10500 22146
rect 10444 22092 10500 22094
rect 10892 24668 10948 24724
rect 10780 22764 10836 22820
rect 9996 21420 10052 21476
rect 10332 20972 10388 21028
rect 10556 20748 10612 20804
rect 10780 21868 10836 21924
rect 10444 20018 10500 20020
rect 10444 19966 10446 20018
rect 10446 19966 10498 20018
rect 10498 19966 10500 20018
rect 10444 19964 10500 19966
rect 10332 19628 10388 19684
rect 9996 18732 10052 18788
rect 10108 19516 10164 19572
rect 9772 18284 9828 18340
rect 9772 17836 9828 17892
rect 10332 19346 10388 19348
rect 10332 19294 10334 19346
rect 10334 19294 10386 19346
rect 10386 19294 10388 19346
rect 10332 19292 10388 19294
rect 10220 19068 10276 19124
rect 10444 19180 10500 19236
rect 10220 18732 10276 18788
rect 10892 19852 10948 19908
rect 10780 19516 10836 19572
rect 10892 19234 10948 19236
rect 10892 19182 10894 19234
rect 10894 19182 10946 19234
rect 10946 19182 10948 19234
rect 10892 19180 10948 19182
rect 10556 18508 10612 18564
rect 9324 17724 9380 17780
rect 9660 17778 9716 17780
rect 9660 17726 9662 17778
rect 9662 17726 9714 17778
rect 9714 17726 9716 17778
rect 9660 17724 9716 17726
rect 8764 16492 8820 16548
rect 8652 15538 8708 15540
rect 8652 15486 8654 15538
rect 8654 15486 8706 15538
rect 8706 15486 8708 15538
rect 8652 15484 8708 15486
rect 8316 13468 8372 13524
rect 8652 14530 8708 14532
rect 8652 14478 8654 14530
rect 8654 14478 8706 14530
rect 8706 14478 8708 14530
rect 8652 14476 8708 14478
rect 8428 12124 8484 12180
rect 8540 14364 8596 14420
rect 9100 16156 9156 16212
rect 8876 15708 8932 15764
rect 8988 15820 9044 15876
rect 8092 11004 8148 11060
rect 7868 10722 7924 10724
rect 7868 10670 7870 10722
rect 7870 10670 7922 10722
rect 7922 10670 7924 10722
rect 7868 10668 7924 10670
rect 7756 10610 7812 10612
rect 7756 10558 7758 10610
rect 7758 10558 7810 10610
rect 7810 10558 7812 10610
rect 7756 10556 7812 10558
rect 7756 8930 7812 8932
rect 7756 8878 7758 8930
rect 7758 8878 7810 8930
rect 7810 8878 7812 8930
rect 7756 8876 7812 8878
rect 7532 8204 7588 8260
rect 7420 7868 7476 7924
rect 7308 7698 7364 7700
rect 7308 7646 7310 7698
rect 7310 7646 7362 7698
rect 7362 7646 7364 7698
rect 7308 7644 7364 7646
rect 8316 10722 8372 10724
rect 8316 10670 8318 10722
rect 8318 10670 8370 10722
rect 8370 10670 8372 10722
rect 8316 10668 8372 10670
rect 8204 10556 8260 10612
rect 8092 9938 8148 9940
rect 8092 9886 8094 9938
rect 8094 9886 8146 9938
rect 8146 9886 8148 9938
rect 8092 9884 8148 9886
rect 7756 7644 7812 7700
rect 7644 6748 7700 6804
rect 7980 7756 8036 7812
rect 7644 5794 7700 5796
rect 7644 5742 7646 5794
rect 7646 5742 7698 5794
rect 7698 5742 7700 5794
rect 7644 5740 7700 5742
rect 7308 5292 7364 5348
rect 7868 5740 7924 5796
rect 7868 4956 7924 5012
rect 7196 4172 7252 4228
rect 8204 9266 8260 9268
rect 8204 9214 8206 9266
rect 8206 9214 8258 9266
rect 8258 9214 8260 9266
rect 8204 9212 8260 9214
rect 9100 15708 9156 15764
rect 8988 15202 9044 15204
rect 8988 15150 8990 15202
rect 8990 15150 9042 15202
rect 9042 15150 9044 15202
rect 8988 15148 9044 15150
rect 8876 13858 8932 13860
rect 8876 13806 8878 13858
rect 8878 13806 8930 13858
rect 8930 13806 8932 13858
rect 8876 13804 8932 13806
rect 8764 13468 8820 13524
rect 10780 18956 10836 19012
rect 10780 18172 10836 18228
rect 10332 17388 10388 17444
rect 9884 17276 9940 17332
rect 10108 17106 10164 17108
rect 10108 17054 10110 17106
rect 10110 17054 10162 17106
rect 10162 17054 10164 17106
rect 10108 17052 10164 17054
rect 10332 17052 10388 17108
rect 9772 16716 9828 16772
rect 9324 16380 9380 16436
rect 9660 16268 9716 16324
rect 11228 25116 11284 25172
rect 11452 28140 11508 28196
rect 11676 27244 11732 27300
rect 11452 26684 11508 26740
rect 11788 26178 11844 26180
rect 11788 26126 11790 26178
rect 11790 26126 11842 26178
rect 11842 26126 11844 26178
rect 11788 26124 11844 26126
rect 11452 25676 11508 25732
rect 11564 25900 11620 25956
rect 11452 25506 11508 25508
rect 11452 25454 11454 25506
rect 11454 25454 11506 25506
rect 11506 25454 11508 25506
rect 11452 25452 11508 25454
rect 11452 24892 11508 24948
rect 11564 23884 11620 23940
rect 11116 22316 11172 22372
rect 11116 21980 11172 22036
rect 11228 22146 11284 22148
rect 11228 22094 11230 22146
rect 11230 22094 11282 22146
rect 11282 22094 11284 22146
rect 11228 22092 11284 22094
rect 11116 19628 11172 19684
rect 10892 17052 10948 17108
rect 11004 17388 11060 17444
rect 11004 16940 11060 16996
rect 10556 16044 10612 16100
rect 10668 15932 10724 15988
rect 10556 15596 10612 15652
rect 9884 15426 9940 15428
rect 9884 15374 9886 15426
rect 9886 15374 9938 15426
rect 9938 15374 9940 15426
rect 9884 15372 9940 15374
rect 11788 24162 11844 24164
rect 11788 24110 11790 24162
rect 11790 24110 11842 24162
rect 11842 24110 11844 24162
rect 11788 24108 11844 24110
rect 11788 23660 11844 23716
rect 11788 22876 11844 22932
rect 11564 20412 11620 20468
rect 11676 20300 11732 20356
rect 11340 19628 11396 19684
rect 11788 19010 11844 19012
rect 11788 18958 11790 19010
rect 11790 18958 11842 19010
rect 11842 18958 11844 19010
rect 11788 18956 11844 18958
rect 11788 18620 11844 18676
rect 11340 18396 11396 18452
rect 11564 18508 11620 18564
rect 11452 18338 11508 18340
rect 11452 18286 11454 18338
rect 11454 18286 11506 18338
rect 11506 18286 11508 18338
rect 11452 18284 11508 18286
rect 11452 17948 11508 18004
rect 11340 16044 11396 16100
rect 10780 15426 10836 15428
rect 10780 15374 10782 15426
rect 10782 15374 10834 15426
rect 10834 15374 10836 15426
rect 10780 15372 10836 15374
rect 9548 14754 9604 14756
rect 9548 14702 9550 14754
rect 9550 14702 9602 14754
rect 9602 14702 9604 14754
rect 9548 14700 9604 14702
rect 9212 13580 9268 13636
rect 9100 12962 9156 12964
rect 9100 12910 9102 12962
rect 9102 12910 9154 12962
rect 9154 12910 9156 12962
rect 9100 12908 9156 12910
rect 8988 11788 9044 11844
rect 8876 11564 8932 11620
rect 8876 11004 8932 11060
rect 8092 6524 8148 6580
rect 8540 8930 8596 8932
rect 8540 8878 8542 8930
rect 8542 8878 8594 8930
rect 8594 8878 8596 8930
rect 8540 8876 8596 8878
rect 8204 7980 8260 8036
rect 8092 6188 8148 6244
rect 8876 8876 8932 8932
rect 8316 7756 8372 7812
rect 8428 8204 8484 8260
rect 8764 8258 8820 8260
rect 8764 8206 8766 8258
rect 8766 8206 8818 8258
rect 8818 8206 8820 8258
rect 8764 8204 8820 8206
rect 8540 7756 8596 7812
rect 8652 7308 8708 7364
rect 8204 5628 8260 5684
rect 8428 5740 8484 5796
rect 8204 4284 8260 4340
rect 7196 2268 7252 2324
rect 6188 1484 6244 1540
rect 8764 5068 8820 5124
rect 8652 4562 8708 4564
rect 8652 4510 8654 4562
rect 8654 4510 8706 4562
rect 8706 4510 8708 4562
rect 8652 4508 8708 4510
rect 9324 11676 9380 11732
rect 8988 8316 9044 8372
rect 9100 8764 9156 8820
rect 8988 8092 9044 8148
rect 8988 6466 9044 6468
rect 8988 6414 8990 6466
rect 8990 6414 9042 6466
rect 9042 6414 9044 6466
rect 8988 6412 9044 6414
rect 9772 14418 9828 14420
rect 9772 14366 9774 14418
rect 9774 14366 9826 14418
rect 9826 14366 9828 14418
rect 9772 14364 9828 14366
rect 9772 13858 9828 13860
rect 9772 13806 9774 13858
rect 9774 13806 9826 13858
rect 9826 13806 9828 13858
rect 9772 13804 9828 13806
rect 9660 12908 9716 12964
rect 10444 14476 10500 14532
rect 10668 14476 10724 14532
rect 10332 14252 10388 14308
rect 10332 13522 10388 13524
rect 10332 13470 10334 13522
rect 10334 13470 10386 13522
rect 10386 13470 10388 13522
rect 10332 13468 10388 13470
rect 10108 13074 10164 13076
rect 10108 13022 10110 13074
rect 10110 13022 10162 13074
rect 10162 13022 10164 13074
rect 10108 13020 10164 13022
rect 10220 12348 10276 12404
rect 9884 12178 9940 12180
rect 9884 12126 9886 12178
rect 9886 12126 9938 12178
rect 9938 12126 9940 12178
rect 9884 12124 9940 12126
rect 10108 11228 10164 11284
rect 10108 10332 10164 10388
rect 10668 12348 10724 12404
rect 11004 14812 11060 14868
rect 10780 14364 10836 14420
rect 10556 12236 10612 12292
rect 10444 11788 10500 11844
rect 10444 11394 10500 11396
rect 10444 11342 10446 11394
rect 10446 11342 10498 11394
rect 10498 11342 10500 11394
rect 10444 11340 10500 11342
rect 9772 9996 9828 10052
rect 10668 11452 10724 11508
rect 11116 14140 11172 14196
rect 11228 13580 11284 13636
rect 12012 28812 12068 28868
rect 12124 30492 12180 30548
rect 12012 27916 12068 27972
rect 12236 29372 12292 29428
rect 12236 27858 12292 27860
rect 12236 27806 12238 27858
rect 12238 27806 12290 27858
rect 12290 27806 12292 27858
rect 12236 27804 12292 27806
rect 12348 28364 12404 28420
rect 12236 27356 12292 27412
rect 12236 26908 12292 26964
rect 12236 26178 12292 26180
rect 12236 26126 12238 26178
rect 12238 26126 12290 26178
rect 12290 26126 12292 26178
rect 12236 26124 12292 26126
rect 13244 34018 13300 34020
rect 13244 33966 13246 34018
rect 13246 33966 13298 34018
rect 13298 33966 13300 34018
rect 13244 33964 13300 33966
rect 12908 33852 12964 33908
rect 13468 36428 13524 36484
rect 13916 36652 13972 36708
rect 14028 36204 14084 36260
rect 14476 40124 14532 40180
rect 16604 45500 16660 45556
rect 14700 44716 14756 44772
rect 14812 44322 14868 44324
rect 14812 44270 14814 44322
rect 14814 44270 14866 44322
rect 14866 44270 14868 44322
rect 14812 44268 14868 44270
rect 15036 43932 15092 43988
rect 15036 43708 15092 43764
rect 15148 43484 15204 43540
rect 19964 49698 20020 49700
rect 19964 49646 19966 49698
rect 19966 49646 20018 49698
rect 20018 49646 20020 49698
rect 19964 49644 20020 49646
rect 20636 49644 20692 49700
rect 20860 48972 20916 49028
rect 17724 48466 17780 48468
rect 17724 48414 17726 48466
rect 17726 48414 17778 48466
rect 17778 48414 17780 48466
rect 17724 48412 17780 48414
rect 17948 48466 18004 48468
rect 17948 48414 17950 48466
rect 17950 48414 18002 48466
rect 18002 48414 18004 48466
rect 17948 48412 18004 48414
rect 18732 48412 18788 48468
rect 17948 48188 18004 48244
rect 18956 48354 19012 48356
rect 18956 48302 18958 48354
rect 18958 48302 19010 48354
rect 19010 48302 19012 48354
rect 18956 48300 19012 48302
rect 19404 47964 19460 48020
rect 18284 47570 18340 47572
rect 18284 47518 18286 47570
rect 18286 47518 18338 47570
rect 18338 47518 18340 47570
rect 18284 47516 18340 47518
rect 18172 47234 18228 47236
rect 18172 47182 18174 47234
rect 18174 47182 18226 47234
rect 18226 47182 18228 47234
rect 18172 47180 18228 47182
rect 17836 46508 17892 46564
rect 18956 47068 19012 47124
rect 16604 43820 16660 43876
rect 15820 43484 15876 43540
rect 15260 42476 15316 42532
rect 14700 42364 14756 42420
rect 15596 42364 15652 42420
rect 14924 42028 14980 42084
rect 14588 40012 14644 40068
rect 14700 40908 14756 40964
rect 14364 39340 14420 39396
rect 14476 39228 14532 39284
rect 14364 37436 14420 37492
rect 14252 37154 14308 37156
rect 14252 37102 14254 37154
rect 14254 37102 14306 37154
rect 14306 37102 14308 37154
rect 14252 37100 14308 37102
rect 14588 37378 14644 37380
rect 14588 37326 14590 37378
rect 14590 37326 14642 37378
rect 14642 37326 14644 37378
rect 14588 37324 14644 37326
rect 14476 36988 14532 37044
rect 13692 34914 13748 34916
rect 13692 34862 13694 34914
rect 13694 34862 13746 34914
rect 13746 34862 13748 34914
rect 13692 34860 13748 34862
rect 13804 34802 13860 34804
rect 13804 34750 13806 34802
rect 13806 34750 13858 34802
rect 13858 34750 13860 34802
rect 13804 34748 13860 34750
rect 13580 34636 13636 34692
rect 14252 35532 14308 35588
rect 15708 41916 15764 41972
rect 15148 40962 15204 40964
rect 15148 40910 15150 40962
rect 15150 40910 15202 40962
rect 15202 40910 15204 40962
rect 15148 40908 15204 40910
rect 15148 40348 15204 40404
rect 14924 39116 14980 39172
rect 14924 38892 14980 38948
rect 14812 38610 14868 38612
rect 14812 38558 14814 38610
rect 14814 38558 14866 38610
rect 14866 38558 14868 38610
rect 14812 38556 14868 38558
rect 15148 38556 15204 38612
rect 15036 38444 15092 38500
rect 15148 38332 15204 38388
rect 14812 37436 14868 37492
rect 14924 37266 14980 37268
rect 14924 37214 14926 37266
rect 14926 37214 14978 37266
rect 14978 37214 14980 37266
rect 14924 37212 14980 37214
rect 15260 37884 15316 37940
rect 15260 37660 15316 37716
rect 15148 37212 15204 37268
rect 15260 36876 15316 36932
rect 14588 36540 14644 36596
rect 14812 36482 14868 36484
rect 14812 36430 14814 36482
rect 14814 36430 14866 36482
rect 14866 36430 14868 36482
rect 14812 36428 14868 36430
rect 14588 36204 14644 36260
rect 14700 36316 14756 36372
rect 14812 34914 14868 34916
rect 14812 34862 14814 34914
rect 14814 34862 14866 34914
rect 14866 34862 14868 34914
rect 14812 34860 14868 34862
rect 13356 33852 13412 33908
rect 13580 33180 13636 33236
rect 12908 33122 12964 33124
rect 12908 33070 12910 33122
rect 12910 33070 12962 33122
rect 12962 33070 12964 33122
rect 12908 33068 12964 33070
rect 13692 33122 13748 33124
rect 13692 33070 13694 33122
rect 13694 33070 13746 33122
rect 13746 33070 13748 33122
rect 13692 33068 13748 33070
rect 12684 32450 12740 32452
rect 12684 32398 12686 32450
rect 12686 32398 12738 32450
rect 12738 32398 12740 32450
rect 12684 32396 12740 32398
rect 12796 31836 12852 31892
rect 12684 31106 12740 31108
rect 12684 31054 12686 31106
rect 12686 31054 12738 31106
rect 12738 31054 12740 31106
rect 12684 31052 12740 31054
rect 12684 29986 12740 29988
rect 12684 29934 12686 29986
rect 12686 29934 12738 29986
rect 12738 29934 12740 29986
rect 12684 29932 12740 29934
rect 13468 32562 13524 32564
rect 13468 32510 13470 32562
rect 13470 32510 13522 32562
rect 13522 32510 13524 32562
rect 13468 32508 13524 32510
rect 13692 32508 13748 32564
rect 14252 33852 14308 33908
rect 14028 32620 14084 32676
rect 13356 31836 13412 31892
rect 14140 32396 14196 32452
rect 12908 29708 12964 29764
rect 13020 30940 13076 30996
rect 12684 29260 12740 29316
rect 12908 29260 12964 29316
rect 12572 28812 12628 28868
rect 12460 26460 12516 26516
rect 12012 24220 12068 24276
rect 12236 22764 12292 22820
rect 12124 21586 12180 21588
rect 12124 21534 12126 21586
rect 12126 21534 12178 21586
rect 12178 21534 12180 21586
rect 12124 21532 12180 21534
rect 13468 29820 13524 29876
rect 14140 32002 14196 32004
rect 14140 31950 14142 32002
rect 14142 31950 14194 32002
rect 14194 31950 14196 32002
rect 14140 31948 14196 31950
rect 13916 31890 13972 31892
rect 13916 31838 13918 31890
rect 13918 31838 13970 31890
rect 13970 31838 13972 31890
rect 13916 31836 13972 31838
rect 15148 36652 15204 36708
rect 15148 36482 15204 36484
rect 15148 36430 15150 36482
rect 15150 36430 15202 36482
rect 15202 36430 15204 36482
rect 15148 36428 15204 36430
rect 15148 34860 15204 34916
rect 15036 34748 15092 34804
rect 15036 34018 15092 34020
rect 15036 33966 15038 34018
rect 15038 33966 15090 34018
rect 15090 33966 15092 34018
rect 15036 33964 15092 33966
rect 14476 32450 14532 32452
rect 14476 32398 14478 32450
rect 14478 32398 14530 32450
rect 14530 32398 14532 32450
rect 14476 32396 14532 32398
rect 15484 38332 15540 38388
rect 15596 38780 15652 38836
rect 15596 37324 15652 37380
rect 15372 36540 15428 36596
rect 15596 36594 15652 36596
rect 15596 36542 15598 36594
rect 15598 36542 15650 36594
rect 15650 36542 15652 36594
rect 15596 36540 15652 36542
rect 15036 32674 15092 32676
rect 15036 32622 15038 32674
rect 15038 32622 15090 32674
rect 15090 32622 15092 32674
rect 15036 32620 15092 32622
rect 13692 30940 13748 30996
rect 14924 32396 14980 32452
rect 13132 28140 13188 28196
rect 13468 28700 13524 28756
rect 12908 27916 12964 27972
rect 12796 27692 12852 27748
rect 13020 27858 13076 27860
rect 13020 27806 13022 27858
rect 13022 27806 13074 27858
rect 13074 27806 13076 27858
rect 13020 27804 13076 27806
rect 13244 27858 13300 27860
rect 13244 27806 13246 27858
rect 13246 27806 13298 27858
rect 13298 27806 13300 27858
rect 13244 27804 13300 27806
rect 13132 27692 13188 27748
rect 12796 27356 12852 27412
rect 12908 27132 12964 27188
rect 13356 27356 13412 27412
rect 14140 30098 14196 30100
rect 14140 30046 14142 30098
rect 14142 30046 14194 30098
rect 14194 30046 14196 30098
rect 14140 30044 14196 30046
rect 14364 29820 14420 29876
rect 14252 29426 14308 29428
rect 14252 29374 14254 29426
rect 14254 29374 14306 29426
rect 14306 29374 14308 29426
rect 14252 29372 14308 29374
rect 14252 28700 14308 28756
rect 14028 28140 14084 28196
rect 14364 28364 14420 28420
rect 14364 28028 14420 28084
rect 14252 27804 14308 27860
rect 13468 27132 13524 27188
rect 12796 26572 12852 26628
rect 12908 26514 12964 26516
rect 12908 26462 12910 26514
rect 12910 26462 12962 26514
rect 12962 26462 12964 26514
rect 12908 26460 12964 26462
rect 12908 25676 12964 25732
rect 13132 26402 13188 26404
rect 13132 26350 13134 26402
rect 13134 26350 13186 26402
rect 13186 26350 13188 26402
rect 13132 26348 13188 26350
rect 13020 25340 13076 25396
rect 12796 25116 12852 25172
rect 12796 24722 12852 24724
rect 12796 24670 12798 24722
rect 12798 24670 12850 24722
rect 12850 24670 12852 24722
rect 12796 24668 12852 24670
rect 13132 23436 13188 23492
rect 12348 20860 12404 20916
rect 12684 22652 12740 22708
rect 12572 22482 12628 22484
rect 12572 22430 12574 22482
rect 12574 22430 12626 22482
rect 12626 22430 12628 22482
rect 12572 22428 12628 22430
rect 12908 21698 12964 21700
rect 12908 21646 12910 21698
rect 12910 21646 12962 21698
rect 12962 21646 12964 21698
rect 12908 21644 12964 21646
rect 12908 21084 12964 21140
rect 13020 21308 13076 21364
rect 12236 20300 12292 20356
rect 12572 20578 12628 20580
rect 12572 20526 12574 20578
rect 12574 20526 12626 20578
rect 12626 20526 12628 20578
rect 12572 20524 12628 20526
rect 12796 20300 12852 20356
rect 12460 19740 12516 19796
rect 12460 19292 12516 19348
rect 12460 18844 12516 18900
rect 12348 18732 12404 18788
rect 11676 17948 11732 18004
rect 11900 17106 11956 17108
rect 11900 17054 11902 17106
rect 11902 17054 11954 17106
rect 11954 17054 11956 17106
rect 11900 17052 11956 17054
rect 12460 18284 12516 18340
rect 12460 17778 12516 17780
rect 12460 17726 12462 17778
rect 12462 17726 12514 17778
rect 12514 17726 12516 17778
rect 12460 17724 12516 17726
rect 12236 16994 12292 16996
rect 12236 16942 12238 16994
rect 12238 16942 12290 16994
rect 12290 16942 12292 16994
rect 12236 16940 12292 16942
rect 12348 16604 12404 16660
rect 12012 16044 12068 16100
rect 12124 15708 12180 15764
rect 12012 15202 12068 15204
rect 12012 15150 12014 15202
rect 12014 15150 12066 15202
rect 12066 15150 12068 15202
rect 12012 15148 12068 15150
rect 11564 13468 11620 13524
rect 11676 14812 11732 14868
rect 11788 14530 11844 14532
rect 11788 14478 11790 14530
rect 11790 14478 11842 14530
rect 11842 14478 11844 14530
rect 11788 14476 11844 14478
rect 9660 9826 9716 9828
rect 9660 9774 9662 9826
rect 9662 9774 9714 9826
rect 9714 9774 9716 9826
rect 9660 9772 9716 9774
rect 9436 8764 9492 8820
rect 9548 9324 9604 9380
rect 9212 6860 9268 6916
rect 9772 9154 9828 9156
rect 9772 9102 9774 9154
rect 9774 9102 9826 9154
rect 9826 9102 9828 9154
rect 9772 9100 9828 9102
rect 9660 7308 9716 7364
rect 9884 8316 9940 8372
rect 9996 8204 10052 8260
rect 9772 6524 9828 6580
rect 9660 5234 9716 5236
rect 9660 5182 9662 5234
rect 9662 5182 9714 5234
rect 9714 5182 9716 5234
rect 9660 5180 9716 5182
rect 9100 4620 9156 4676
rect 8988 4226 9044 4228
rect 8988 4174 8990 4226
rect 8990 4174 9042 4226
rect 9042 4174 9044 4226
rect 8988 4172 9044 4174
rect 8988 3612 9044 3668
rect 10332 8316 10388 8372
rect 10220 7756 10276 7812
rect 10220 7084 10276 7140
rect 10108 6300 10164 6356
rect 9996 5516 10052 5572
rect 10220 6076 10276 6132
rect 10332 6636 10388 6692
rect 10332 6412 10388 6468
rect 10780 10668 10836 10724
rect 10668 9548 10724 9604
rect 10556 7196 10612 7252
rect 11564 12348 11620 12404
rect 11116 12290 11172 12292
rect 11116 12238 11118 12290
rect 11118 12238 11170 12290
rect 11170 12238 11172 12290
rect 11116 12236 11172 12238
rect 11004 12012 11060 12068
rect 11228 12124 11284 12180
rect 11004 11788 11060 11844
rect 10668 6748 10724 6804
rect 10780 8258 10836 8260
rect 10780 8206 10782 8258
rect 10782 8206 10834 8258
rect 10834 8206 10836 8258
rect 10780 8204 10836 8206
rect 10668 6412 10724 6468
rect 10892 7532 10948 7588
rect 10780 6188 10836 6244
rect 11116 11452 11172 11508
rect 10556 5234 10612 5236
rect 10556 5182 10558 5234
rect 10558 5182 10610 5234
rect 10610 5182 10612 5234
rect 10556 5180 10612 5182
rect 11004 6748 11060 6804
rect 10892 4956 10948 5012
rect 10668 4508 10724 4564
rect 10108 3666 10164 3668
rect 10108 3614 10110 3666
rect 10110 3614 10162 3666
rect 10162 3614 10164 3666
rect 10108 3612 10164 3614
rect 11228 10556 11284 10612
rect 11676 12572 11732 12628
rect 11788 11564 11844 11620
rect 11564 10892 11620 10948
rect 11228 9772 11284 9828
rect 11340 6748 11396 6804
rect 12124 15036 12180 15092
rect 12460 16380 12516 16436
rect 12684 19964 12740 20020
rect 12684 19180 12740 19236
rect 12908 19234 12964 19236
rect 12908 19182 12910 19234
rect 12910 19182 12962 19234
rect 12962 19182 12964 19234
rect 12908 19180 12964 19182
rect 13356 25452 13412 25508
rect 13580 27356 13636 27412
rect 14700 31724 14756 31780
rect 16044 41746 16100 41748
rect 16044 41694 16046 41746
rect 16046 41694 16098 41746
rect 16098 41694 16100 41746
rect 16044 41692 16100 41694
rect 16268 43538 16324 43540
rect 16268 43486 16270 43538
rect 16270 43486 16322 43538
rect 16322 43486 16324 43538
rect 16268 43484 16324 43486
rect 17724 44156 17780 44212
rect 17276 43932 17332 43988
rect 16268 42530 16324 42532
rect 16268 42478 16270 42530
rect 16270 42478 16322 42530
rect 16322 42478 16324 42530
rect 16268 42476 16324 42478
rect 16492 42028 16548 42084
rect 16716 41970 16772 41972
rect 16716 41918 16718 41970
rect 16718 41918 16770 41970
rect 16770 41918 16772 41970
rect 16716 41916 16772 41918
rect 17052 42028 17108 42084
rect 17164 42476 17220 42532
rect 16604 41244 16660 41300
rect 15820 40908 15876 40964
rect 16044 40402 16100 40404
rect 16044 40350 16046 40402
rect 16046 40350 16098 40402
rect 16098 40350 16100 40402
rect 16044 40348 16100 40350
rect 16380 40348 16436 40404
rect 16044 40124 16100 40180
rect 16044 39228 16100 39284
rect 16044 38780 16100 38836
rect 16156 38444 16212 38500
rect 16044 37938 16100 37940
rect 16044 37886 16046 37938
rect 16046 37886 16098 37938
rect 16098 37886 16100 37938
rect 16044 37884 16100 37886
rect 15932 37826 15988 37828
rect 15932 37774 15934 37826
rect 15934 37774 15986 37826
rect 15986 37774 15988 37826
rect 15932 37772 15988 37774
rect 16156 37772 16212 37828
rect 16940 40124 16996 40180
rect 16604 38834 16660 38836
rect 16604 38782 16606 38834
rect 16606 38782 16658 38834
rect 16658 38782 16660 38834
rect 16604 38780 16660 38782
rect 16940 39340 16996 39396
rect 16380 37436 16436 37492
rect 16044 37212 16100 37268
rect 15820 36540 15876 36596
rect 16044 36428 16100 36484
rect 15932 34802 15988 34804
rect 15932 34750 15934 34802
rect 15934 34750 15986 34802
rect 15986 34750 15988 34802
rect 15932 34748 15988 34750
rect 15820 34018 15876 34020
rect 15820 33966 15822 34018
rect 15822 33966 15874 34018
rect 15874 33966 15876 34018
rect 15820 33964 15876 33966
rect 15932 33852 15988 33908
rect 15932 33628 15988 33684
rect 15820 33516 15876 33572
rect 14588 29372 14644 29428
rect 15148 30098 15204 30100
rect 15148 30046 15150 30098
rect 15150 30046 15202 30098
rect 15202 30046 15204 30098
rect 15148 30044 15204 30046
rect 15372 30492 15428 30548
rect 15260 29820 15316 29876
rect 15820 29484 15876 29540
rect 15596 29260 15652 29316
rect 15484 28588 15540 28644
rect 14588 27804 14644 27860
rect 14700 28252 14756 28308
rect 15708 29148 15764 29204
rect 15484 28252 15540 28308
rect 15260 27858 15316 27860
rect 15260 27806 15262 27858
rect 15262 27806 15314 27858
rect 15314 27806 15316 27858
rect 15260 27804 15316 27806
rect 15708 27916 15764 27972
rect 15820 28140 15876 28196
rect 14924 27356 14980 27412
rect 15372 27074 15428 27076
rect 15372 27022 15374 27074
rect 15374 27022 15426 27074
rect 15426 27022 15428 27074
rect 15372 27020 15428 27022
rect 13580 26908 13636 26964
rect 13804 26962 13860 26964
rect 13804 26910 13806 26962
rect 13806 26910 13858 26962
rect 13858 26910 13860 26962
rect 13804 26908 13860 26910
rect 14588 26908 14644 26964
rect 15596 26796 15652 26852
rect 14924 26684 14980 26740
rect 14588 26402 14644 26404
rect 14588 26350 14590 26402
rect 14590 26350 14642 26402
rect 14642 26350 14644 26402
rect 14588 26348 14644 26350
rect 14364 26236 14420 26292
rect 14476 26178 14532 26180
rect 14476 26126 14478 26178
rect 14478 26126 14530 26178
rect 14530 26126 14532 26178
rect 14476 26124 14532 26126
rect 14364 25900 14420 25956
rect 14476 25618 14532 25620
rect 14476 25566 14478 25618
rect 14478 25566 14530 25618
rect 14530 25566 14532 25618
rect 14476 25564 14532 25566
rect 14028 25394 14084 25396
rect 14028 25342 14030 25394
rect 14030 25342 14082 25394
rect 14082 25342 14084 25394
rect 14028 25340 14084 25342
rect 13468 24556 13524 24612
rect 13468 24220 13524 24276
rect 13916 25116 13972 25172
rect 14476 25340 14532 25396
rect 13804 24108 13860 24164
rect 13916 23884 13972 23940
rect 13804 23826 13860 23828
rect 13804 23774 13806 23826
rect 13806 23774 13858 23826
rect 13858 23774 13860 23826
rect 13804 23772 13860 23774
rect 13468 23324 13524 23380
rect 13356 21868 13412 21924
rect 13468 22540 13524 22596
rect 13916 22092 13972 22148
rect 13244 20860 13300 20916
rect 13580 21420 13636 21476
rect 13580 21196 13636 21252
rect 13020 18620 13076 18676
rect 13132 19292 13188 19348
rect 12684 18396 12740 18452
rect 12908 17612 12964 17668
rect 12684 17052 12740 17108
rect 12572 15596 12628 15652
rect 12124 14754 12180 14756
rect 12124 14702 12126 14754
rect 12126 14702 12178 14754
rect 12178 14702 12180 14754
rect 12124 14700 12180 14702
rect 12012 14418 12068 14420
rect 12012 14366 12014 14418
rect 12014 14366 12066 14418
rect 12066 14366 12068 14418
rect 12012 14364 12068 14366
rect 12012 13580 12068 13636
rect 12124 13356 12180 13412
rect 13692 20972 13748 21028
rect 13468 19516 13524 19572
rect 13356 18338 13412 18340
rect 13356 18286 13358 18338
rect 13358 18286 13410 18338
rect 13410 18286 13412 18338
rect 13356 18284 13412 18286
rect 13804 19906 13860 19908
rect 13804 19854 13806 19906
rect 13806 19854 13858 19906
rect 13858 19854 13860 19906
rect 13804 19852 13860 19854
rect 14252 22652 14308 22708
rect 14252 22204 14308 22260
rect 14140 21756 14196 21812
rect 14028 20018 14084 20020
rect 14028 19966 14030 20018
rect 14030 19966 14082 20018
rect 14082 19966 14084 20018
rect 14028 19964 14084 19966
rect 15596 26402 15652 26404
rect 15596 26350 15598 26402
rect 15598 26350 15650 26402
rect 15650 26350 15652 26402
rect 15596 26348 15652 26350
rect 15484 26066 15540 26068
rect 15484 26014 15486 26066
rect 15486 26014 15538 26066
rect 15538 26014 15540 26066
rect 15484 26012 15540 26014
rect 15148 25004 15204 25060
rect 15260 25116 15316 25172
rect 15036 24780 15092 24836
rect 14476 24220 14532 24276
rect 14700 23772 14756 23828
rect 14588 23266 14644 23268
rect 14588 23214 14590 23266
rect 14590 23214 14642 23266
rect 14642 23214 14644 23266
rect 14588 23212 14644 23214
rect 14924 23772 14980 23828
rect 14812 23154 14868 23156
rect 14812 23102 14814 23154
rect 14814 23102 14866 23154
rect 14866 23102 14868 23154
rect 14812 23100 14868 23102
rect 14588 22092 14644 22148
rect 14700 21586 14756 21588
rect 14700 21534 14702 21586
rect 14702 21534 14754 21586
rect 14754 21534 14756 21586
rect 14700 21532 14756 21534
rect 15260 24332 15316 24388
rect 15148 24220 15204 24276
rect 15484 25116 15540 25172
rect 15708 25004 15764 25060
rect 15708 24780 15764 24836
rect 15148 23660 15204 23716
rect 15036 22204 15092 22260
rect 15148 23324 15204 23380
rect 15260 23266 15316 23268
rect 15260 23214 15262 23266
rect 15262 23214 15314 23266
rect 15314 23214 15316 23266
rect 15260 23212 15316 23214
rect 15148 23100 15204 23156
rect 14252 20690 14308 20692
rect 14252 20638 14254 20690
rect 14254 20638 14306 20690
rect 14306 20638 14308 20690
rect 14252 20636 14308 20638
rect 13916 19516 13972 19572
rect 14252 19740 14308 19796
rect 13916 19346 13972 19348
rect 13916 19294 13918 19346
rect 13918 19294 13970 19346
rect 13970 19294 13972 19346
rect 13916 19292 13972 19294
rect 13804 19234 13860 19236
rect 13804 19182 13806 19234
rect 13806 19182 13858 19234
rect 13858 19182 13860 19234
rect 13804 19180 13860 19182
rect 13916 18732 13972 18788
rect 13468 17724 13524 17780
rect 13580 18172 13636 18228
rect 14140 19068 14196 19124
rect 14252 18956 14308 19012
rect 14588 20802 14644 20804
rect 14588 20750 14590 20802
rect 14590 20750 14642 20802
rect 14642 20750 14644 20802
rect 14588 20748 14644 20750
rect 14812 20524 14868 20580
rect 14700 20188 14756 20244
rect 14700 19852 14756 19908
rect 14700 19404 14756 19460
rect 14924 19180 14980 19236
rect 13244 16882 13300 16884
rect 13244 16830 13246 16882
rect 13246 16830 13298 16882
rect 13298 16830 13300 16882
rect 13244 16828 13300 16830
rect 12908 16604 12964 16660
rect 12908 16210 12964 16212
rect 12908 16158 12910 16210
rect 12910 16158 12962 16210
rect 12962 16158 12964 16210
rect 12908 16156 12964 16158
rect 13356 16156 13412 16212
rect 13020 16044 13076 16100
rect 13132 15820 13188 15876
rect 12908 15372 12964 15428
rect 13020 15148 13076 15204
rect 12684 14700 12740 14756
rect 13356 15596 13412 15652
rect 12348 13244 12404 13300
rect 12572 14028 12628 14084
rect 12236 12402 12292 12404
rect 12236 12350 12238 12402
rect 12238 12350 12290 12402
rect 12290 12350 12292 12402
rect 12236 12348 12292 12350
rect 12012 11564 12068 11620
rect 11900 9884 11956 9940
rect 12796 14252 12852 14308
rect 13244 14028 13300 14084
rect 12684 12796 12740 12852
rect 12908 12796 12964 12852
rect 12572 12572 12628 12628
rect 13020 12572 13076 12628
rect 12796 12460 12852 12516
rect 12796 12236 12852 12292
rect 11676 9266 11732 9268
rect 11676 9214 11678 9266
rect 11678 9214 11730 9266
rect 11730 9214 11732 9266
rect 11676 9212 11732 9214
rect 11676 8370 11732 8372
rect 11676 8318 11678 8370
rect 11678 8318 11730 8370
rect 11730 8318 11732 8370
rect 11676 8316 11732 8318
rect 11788 8146 11844 8148
rect 11788 8094 11790 8146
rect 11790 8094 11842 8146
rect 11842 8094 11844 8146
rect 11788 8092 11844 8094
rect 11676 7868 11732 7924
rect 11564 7084 11620 7140
rect 11788 7644 11844 7700
rect 11452 6412 11508 6468
rect 11564 5234 11620 5236
rect 11564 5182 11566 5234
rect 11566 5182 11618 5234
rect 11618 5182 11620 5234
rect 11564 5180 11620 5182
rect 11228 4508 11284 4564
rect 11340 5068 11396 5124
rect 11340 4172 11396 4228
rect 12348 11282 12404 11284
rect 12348 11230 12350 11282
rect 12350 11230 12402 11282
rect 12402 11230 12404 11282
rect 12348 11228 12404 11230
rect 12012 7644 12068 7700
rect 12236 9042 12292 9044
rect 12236 8990 12238 9042
rect 12238 8990 12290 9042
rect 12290 8990 12292 9042
rect 12236 8988 12292 8990
rect 12124 7586 12180 7588
rect 12124 7534 12126 7586
rect 12126 7534 12178 7586
rect 12178 7534 12180 7586
rect 12124 7532 12180 7534
rect 12348 8204 12404 8260
rect 12348 7196 12404 7252
rect 12908 11788 12964 11844
rect 12684 9996 12740 10052
rect 12796 9884 12852 9940
rect 12572 8988 12628 9044
rect 13132 12402 13188 12404
rect 13132 12350 13134 12402
rect 13134 12350 13186 12402
rect 13186 12350 13188 12402
rect 13132 12348 13188 12350
rect 12460 7644 12516 7700
rect 12236 6802 12292 6804
rect 12236 6750 12238 6802
rect 12238 6750 12290 6802
rect 12290 6750 12292 6802
rect 12236 6748 12292 6750
rect 12124 6690 12180 6692
rect 12124 6638 12126 6690
rect 12126 6638 12178 6690
rect 12178 6638 12180 6690
rect 12124 6636 12180 6638
rect 12460 5516 12516 5572
rect 12684 7532 12740 7588
rect 11900 5180 11956 5236
rect 12348 5292 12404 5348
rect 13916 17724 13972 17780
rect 13804 17666 13860 17668
rect 13804 17614 13806 17666
rect 13806 17614 13858 17666
rect 13858 17614 13860 17666
rect 13804 17612 13860 17614
rect 13804 17388 13860 17444
rect 13804 15874 13860 15876
rect 13804 15822 13806 15874
rect 13806 15822 13858 15874
rect 13858 15822 13860 15874
rect 13804 15820 13860 15822
rect 13580 15372 13636 15428
rect 13804 15596 13860 15652
rect 13692 14812 13748 14868
rect 13804 15036 13860 15092
rect 14028 14700 14084 14756
rect 13692 14028 13748 14084
rect 13916 14028 13972 14084
rect 13468 13916 13524 13972
rect 13356 13132 13412 13188
rect 13580 13356 13636 13412
rect 13468 12290 13524 12292
rect 13468 12238 13470 12290
rect 13470 12238 13522 12290
rect 13522 12238 13524 12290
rect 13468 12236 13524 12238
rect 13356 10610 13412 10612
rect 13356 10558 13358 10610
rect 13358 10558 13410 10610
rect 13410 10558 13412 10610
rect 13356 10556 13412 10558
rect 12908 6300 12964 6356
rect 13020 6636 13076 6692
rect 13244 6300 13300 6356
rect 13132 6018 13188 6020
rect 13132 5966 13134 6018
rect 13134 5966 13186 6018
rect 13186 5966 13188 6018
rect 13132 5964 13188 5966
rect 13244 5852 13300 5908
rect 13804 12738 13860 12740
rect 13804 12686 13806 12738
rect 13806 12686 13858 12738
rect 13858 12686 13860 12738
rect 13804 12684 13860 12686
rect 14364 17666 14420 17668
rect 14364 17614 14366 17666
rect 14366 17614 14418 17666
rect 14418 17614 14420 17666
rect 14364 17612 14420 17614
rect 14476 17052 14532 17108
rect 14252 15708 14308 15764
rect 14700 18226 14756 18228
rect 14700 18174 14702 18226
rect 14702 18174 14754 18226
rect 14754 18174 14756 18226
rect 14700 18172 14756 18174
rect 15372 21868 15428 21924
rect 15372 21586 15428 21588
rect 15372 21534 15374 21586
rect 15374 21534 15426 21586
rect 15426 21534 15428 21586
rect 15372 21532 15428 21534
rect 15596 23714 15652 23716
rect 15596 23662 15598 23714
rect 15598 23662 15650 23714
rect 15650 23662 15652 23714
rect 15596 23660 15652 23662
rect 15708 23100 15764 23156
rect 15596 22988 15652 23044
rect 15596 22652 15652 22708
rect 16492 38444 16548 38500
rect 16604 37772 16660 37828
rect 16940 38556 16996 38612
rect 16492 36204 16548 36260
rect 16940 36764 16996 36820
rect 17836 43596 17892 43652
rect 17948 44716 18004 44772
rect 17612 42252 17668 42308
rect 17836 41298 17892 41300
rect 17836 41246 17838 41298
rect 17838 41246 17890 41298
rect 17890 41246 17892 41298
rect 17836 41244 17892 41246
rect 17612 40460 17668 40516
rect 17724 40402 17780 40404
rect 17724 40350 17726 40402
rect 17726 40350 17778 40402
rect 17778 40350 17780 40402
rect 17724 40348 17780 40350
rect 17164 39452 17220 39508
rect 17164 38668 17220 38724
rect 17388 38444 17444 38500
rect 17724 38834 17780 38836
rect 17724 38782 17726 38834
rect 17726 38782 17778 38834
rect 17778 38782 17780 38834
rect 17724 38780 17780 38782
rect 17612 38050 17668 38052
rect 17612 37998 17614 38050
rect 17614 37998 17666 38050
rect 17666 37998 17668 38050
rect 17612 37996 17668 37998
rect 17724 38332 17780 38388
rect 17724 37154 17780 37156
rect 17724 37102 17726 37154
rect 17726 37102 17778 37154
rect 17778 37102 17780 37154
rect 17724 37100 17780 37102
rect 17164 36764 17220 36820
rect 17052 36428 17108 36484
rect 17276 36204 17332 36260
rect 17724 36258 17780 36260
rect 17724 36206 17726 36258
rect 17726 36206 17778 36258
rect 17778 36206 17780 36258
rect 17724 36204 17780 36206
rect 16492 34860 16548 34916
rect 18172 44322 18228 44324
rect 18172 44270 18174 44322
rect 18174 44270 18226 44322
rect 18226 44270 18228 44322
rect 18172 44268 18228 44270
rect 18396 46284 18452 46340
rect 18620 46674 18676 46676
rect 18620 46622 18622 46674
rect 18622 46622 18674 46674
rect 18674 46622 18676 46674
rect 18620 46620 18676 46622
rect 18508 45500 18564 45556
rect 18508 45106 18564 45108
rect 18508 45054 18510 45106
rect 18510 45054 18562 45106
rect 18562 45054 18564 45106
rect 18508 45052 18564 45054
rect 18732 45052 18788 45108
rect 18396 44210 18452 44212
rect 18396 44158 18398 44210
rect 18398 44158 18450 44210
rect 18450 44158 18452 44210
rect 18396 44156 18452 44158
rect 18620 43820 18676 43876
rect 18508 43650 18564 43652
rect 18508 43598 18510 43650
rect 18510 43598 18562 43650
rect 18562 43598 18564 43650
rect 18508 43596 18564 43598
rect 18060 42530 18116 42532
rect 18060 42478 18062 42530
rect 18062 42478 18114 42530
rect 18114 42478 18116 42530
rect 18060 42476 18116 42478
rect 18060 41970 18116 41972
rect 18060 41918 18062 41970
rect 18062 41918 18114 41970
rect 18114 41918 18116 41970
rect 18060 41916 18116 41918
rect 18844 44156 18900 44212
rect 19068 46396 19124 46452
rect 19180 46284 19236 46340
rect 19068 45724 19124 45780
rect 19292 45500 19348 45556
rect 19068 44268 19124 44324
rect 18956 43820 19012 43876
rect 18284 41692 18340 41748
rect 18844 42364 18900 42420
rect 18172 40236 18228 40292
rect 18060 39394 18116 39396
rect 18060 39342 18062 39394
rect 18062 39342 18114 39394
rect 18114 39342 18116 39394
rect 18060 39340 18116 39342
rect 17948 38892 18004 38948
rect 19516 47740 19572 47796
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 21196 48466 21252 48468
rect 21196 48414 21198 48466
rect 21198 48414 21250 48466
rect 21250 48414 21252 48466
rect 21196 48412 21252 48414
rect 19516 46620 19572 46676
rect 19740 47516 19796 47572
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19740 46562 19796 46564
rect 19740 46510 19742 46562
rect 19742 46510 19794 46562
rect 19794 46510 19796 46562
rect 19740 46508 19796 46510
rect 20188 46450 20244 46452
rect 20188 46398 20190 46450
rect 20190 46398 20242 46450
rect 20242 46398 20244 46450
rect 20188 46396 20244 46398
rect 19964 45778 20020 45780
rect 19964 45726 19966 45778
rect 19966 45726 20018 45778
rect 20018 45726 20020 45778
rect 19964 45724 20020 45726
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 27020 55916 27076 55972
rect 27580 55970 27636 55972
rect 27580 55918 27582 55970
rect 27582 55918 27634 55970
rect 27634 55918 27636 55970
rect 27580 55916 27636 55918
rect 23660 55804 23716 55860
rect 22876 55074 22932 55076
rect 22876 55022 22878 55074
rect 22878 55022 22930 55074
rect 22930 55022 22932 55074
rect 22876 55020 22932 55022
rect 27132 55244 27188 55300
rect 23324 55020 23380 55076
rect 21532 49810 21588 49812
rect 21532 49758 21534 49810
rect 21534 49758 21586 49810
rect 21586 49758 21588 49810
rect 21532 49756 21588 49758
rect 21756 49138 21812 49140
rect 21756 49086 21758 49138
rect 21758 49086 21810 49138
rect 21810 49086 21812 49138
rect 21756 49084 21812 49086
rect 21644 49026 21700 49028
rect 21644 48974 21646 49026
rect 21646 48974 21698 49026
rect 21698 48974 21700 49026
rect 21644 48972 21700 48974
rect 22764 50594 22820 50596
rect 22764 50542 22766 50594
rect 22766 50542 22818 50594
rect 22818 50542 22820 50594
rect 22764 50540 22820 50542
rect 22204 49810 22260 49812
rect 22204 49758 22206 49810
rect 22206 49758 22258 49810
rect 22258 49758 22260 49810
rect 22204 49756 22260 49758
rect 22428 49810 22484 49812
rect 22428 49758 22430 49810
rect 22430 49758 22482 49810
rect 22482 49758 22484 49810
rect 22428 49756 22484 49758
rect 24108 51378 24164 51380
rect 24108 51326 24110 51378
rect 24110 51326 24162 51378
rect 24162 51326 24164 51378
rect 24108 51324 24164 51326
rect 24220 51100 24276 51156
rect 23660 50316 23716 50372
rect 23436 49756 23492 49812
rect 21868 48466 21924 48468
rect 21868 48414 21870 48466
rect 21870 48414 21922 48466
rect 21922 48414 21924 48466
rect 21868 48412 21924 48414
rect 23436 49586 23492 49588
rect 23436 49534 23438 49586
rect 23438 49534 23490 49586
rect 23490 49534 23492 49586
rect 23436 49532 23492 49534
rect 23996 50316 24052 50372
rect 23660 49084 23716 49140
rect 22428 48412 22484 48468
rect 21980 48354 22036 48356
rect 21980 48302 21982 48354
rect 21982 48302 22034 48354
rect 22034 48302 22036 48354
rect 21980 48300 22036 48302
rect 22316 48300 22372 48356
rect 22428 48076 22484 48132
rect 23436 48242 23492 48244
rect 23436 48190 23438 48242
rect 23438 48190 23490 48242
rect 23490 48190 23492 48242
rect 23436 48188 23492 48190
rect 23212 48076 23268 48132
rect 24668 51324 24724 51380
rect 24668 49532 24724 49588
rect 23996 49084 24052 49140
rect 26124 51154 26180 51156
rect 26124 51102 26126 51154
rect 26126 51102 26178 51154
rect 26178 51102 26180 51154
rect 26124 51100 26180 51102
rect 26124 50876 26180 50932
rect 25004 49868 25060 49924
rect 25228 50428 25284 50484
rect 24892 48748 24948 48804
rect 24332 48354 24388 48356
rect 24332 48302 24334 48354
rect 24334 48302 24386 48354
rect 24386 48302 24388 48354
rect 24332 48300 24388 48302
rect 24108 48242 24164 48244
rect 24108 48190 24110 48242
rect 24110 48190 24162 48242
rect 24162 48190 24164 48242
rect 24108 48188 24164 48190
rect 21868 47404 21924 47460
rect 22988 47292 23044 47348
rect 22652 46898 22708 46900
rect 22652 46846 22654 46898
rect 22654 46846 22706 46898
rect 22706 46846 22708 46898
rect 22652 46844 22708 46846
rect 23436 47458 23492 47460
rect 23436 47406 23438 47458
rect 23438 47406 23490 47458
rect 23490 47406 23492 47458
rect 23436 47404 23492 47406
rect 23772 47458 23828 47460
rect 23772 47406 23774 47458
rect 23774 47406 23826 47458
rect 23826 47406 23828 47458
rect 23772 47404 23828 47406
rect 23548 47346 23604 47348
rect 23548 47294 23550 47346
rect 23550 47294 23602 47346
rect 23602 47294 23604 47346
rect 23548 47292 23604 47294
rect 24892 48130 24948 48132
rect 24892 48078 24894 48130
rect 24894 48078 24946 48130
rect 24946 48078 24948 48130
rect 24892 48076 24948 48078
rect 24444 47292 24500 47348
rect 24892 47740 24948 47796
rect 23212 46898 23268 46900
rect 23212 46846 23214 46898
rect 23214 46846 23266 46898
rect 23266 46846 23268 46898
rect 23212 46844 23268 46846
rect 24108 46844 24164 46900
rect 23324 46620 23380 46676
rect 19964 45106 20020 45108
rect 19964 45054 19966 45106
rect 19966 45054 20018 45106
rect 20018 45054 20020 45106
rect 19964 45052 20020 45054
rect 20300 44994 20356 44996
rect 20300 44942 20302 44994
rect 20302 44942 20354 44994
rect 20354 44942 20356 44994
rect 20300 44940 20356 44942
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19180 42476 19236 42532
rect 21420 45276 21476 45332
rect 20972 45164 21028 45220
rect 20524 44940 20580 44996
rect 20860 44994 20916 44996
rect 20860 44942 20862 44994
rect 20862 44942 20914 44994
rect 20914 44942 20916 44994
rect 20860 44940 20916 44942
rect 20300 43538 20356 43540
rect 20300 43486 20302 43538
rect 20302 43486 20354 43538
rect 20354 43486 20356 43538
rect 20300 43484 20356 43486
rect 18844 40348 18900 40404
rect 18732 40236 18788 40292
rect 19516 42588 19572 42644
rect 19740 42530 19796 42532
rect 19740 42478 19742 42530
rect 19742 42478 19794 42530
rect 19794 42478 19796 42530
rect 19740 42476 19796 42478
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 22428 43708 22484 43764
rect 21420 43538 21476 43540
rect 21420 43486 21422 43538
rect 21422 43486 21474 43538
rect 21474 43486 21476 43538
rect 21420 43484 21476 43486
rect 23212 45836 23268 45892
rect 22988 45218 23044 45220
rect 22988 45166 22990 45218
rect 22990 45166 23042 45218
rect 23042 45166 23044 45218
rect 22988 45164 23044 45166
rect 23100 44322 23156 44324
rect 23100 44270 23102 44322
rect 23102 44270 23154 44322
rect 23154 44270 23156 44322
rect 23100 44268 23156 44270
rect 23660 44322 23716 44324
rect 23660 44270 23662 44322
rect 23662 44270 23714 44322
rect 23714 44270 23716 44322
rect 23660 44268 23716 44270
rect 23100 43708 23156 43764
rect 24668 46674 24724 46676
rect 24668 46622 24670 46674
rect 24670 46622 24722 46674
rect 24722 46622 24724 46674
rect 24668 46620 24724 46622
rect 24780 45948 24836 46004
rect 25004 46172 25060 46228
rect 24220 45836 24276 45892
rect 24892 45890 24948 45892
rect 24892 45838 24894 45890
rect 24894 45838 24946 45890
rect 24946 45838 24948 45890
rect 24892 45836 24948 45838
rect 24220 45388 24276 45444
rect 24668 44380 24724 44436
rect 24332 44322 24388 44324
rect 24332 44270 24334 44322
rect 24334 44270 24386 44322
rect 24386 44270 24388 44322
rect 24332 44268 24388 44270
rect 20860 43314 20916 43316
rect 20860 43262 20862 43314
rect 20862 43262 20914 43314
rect 20914 43262 20916 43314
rect 20860 43260 20916 43262
rect 21196 43148 21252 43204
rect 20188 42194 20244 42196
rect 20188 42142 20190 42194
rect 20190 42142 20242 42194
rect 20242 42142 20244 42194
rect 20188 42140 20244 42142
rect 20748 42476 20804 42532
rect 19404 41804 19460 41860
rect 19628 40962 19684 40964
rect 19628 40910 19630 40962
rect 19630 40910 19682 40962
rect 19682 40910 19684 40962
rect 19628 40908 19684 40910
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19404 40514 19460 40516
rect 19404 40462 19406 40514
rect 19406 40462 19458 40514
rect 19458 40462 19460 40514
rect 19404 40460 19460 40462
rect 19292 40402 19348 40404
rect 19292 40350 19294 40402
rect 19294 40350 19346 40402
rect 19346 40350 19348 40402
rect 19292 40348 19348 40350
rect 18732 38332 18788 38388
rect 20300 40402 20356 40404
rect 20300 40350 20302 40402
rect 20302 40350 20354 40402
rect 20354 40350 20356 40402
rect 20300 40348 20356 40350
rect 20748 41746 20804 41748
rect 20748 41694 20750 41746
rect 20750 41694 20802 41746
rect 20802 41694 20804 41746
rect 20748 41692 20804 41694
rect 20524 40514 20580 40516
rect 20524 40462 20526 40514
rect 20526 40462 20578 40514
rect 20578 40462 20580 40514
rect 20524 40460 20580 40462
rect 18956 39676 19012 39732
rect 20524 39676 20580 39732
rect 19964 39618 20020 39620
rect 19964 39566 19966 39618
rect 19966 39566 20018 39618
rect 20018 39566 20020 39618
rect 19964 39564 20020 39566
rect 19404 39452 19460 39508
rect 20188 39506 20244 39508
rect 20188 39454 20190 39506
rect 20190 39454 20242 39506
rect 20242 39454 20244 39506
rect 20188 39452 20244 39454
rect 19964 39340 20020 39396
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19180 38444 19236 38500
rect 18172 37436 18228 37492
rect 18060 37324 18116 37380
rect 17948 36428 18004 36484
rect 16604 34354 16660 34356
rect 16604 34302 16606 34354
rect 16606 34302 16658 34354
rect 16658 34302 16660 34354
rect 16604 34300 16660 34302
rect 18172 36988 18228 37044
rect 18172 36764 18228 36820
rect 18172 34188 18228 34244
rect 18284 35532 18340 35588
rect 16604 33964 16660 34020
rect 16044 33404 16100 33460
rect 17612 33740 17668 33796
rect 18060 33740 18116 33796
rect 16156 32508 16212 32564
rect 16604 33122 16660 33124
rect 16604 33070 16606 33122
rect 16606 33070 16658 33122
rect 16658 33070 16660 33122
rect 16604 33068 16660 33070
rect 16492 32620 16548 32676
rect 16380 32508 16436 32564
rect 16156 32172 16212 32228
rect 16044 31890 16100 31892
rect 16044 31838 16046 31890
rect 16046 31838 16098 31890
rect 16098 31838 16100 31890
rect 16044 31836 16100 31838
rect 16156 31948 16212 32004
rect 16044 30882 16100 30884
rect 16044 30830 16046 30882
rect 16046 30830 16098 30882
rect 16098 30830 16100 30882
rect 16044 30828 16100 30830
rect 16044 28588 16100 28644
rect 16044 27580 16100 27636
rect 16044 25282 16100 25284
rect 16044 25230 16046 25282
rect 16046 25230 16098 25282
rect 16098 25230 16100 25282
rect 16044 25228 16100 25230
rect 15932 25116 15988 25172
rect 16044 24332 16100 24388
rect 16044 23436 16100 23492
rect 15820 22652 15876 22708
rect 16044 23212 16100 23268
rect 15708 22092 15764 22148
rect 15708 21644 15764 21700
rect 15820 21868 15876 21924
rect 15372 20972 15428 21028
rect 15372 19516 15428 19572
rect 15484 19458 15540 19460
rect 15484 19406 15486 19458
rect 15486 19406 15538 19458
rect 15538 19406 15540 19458
rect 15484 19404 15540 19406
rect 15260 19122 15316 19124
rect 15260 19070 15262 19122
rect 15262 19070 15314 19122
rect 15314 19070 15316 19122
rect 15260 19068 15316 19070
rect 15820 21084 15876 21140
rect 15708 20076 15764 20132
rect 15372 18562 15428 18564
rect 15372 18510 15374 18562
rect 15374 18510 15426 18562
rect 15426 18510 15428 18562
rect 15372 18508 15428 18510
rect 14924 17836 14980 17892
rect 15148 17666 15204 17668
rect 15148 17614 15150 17666
rect 15150 17614 15202 17666
rect 15202 17614 15204 17666
rect 15148 17612 15204 17614
rect 14812 17052 14868 17108
rect 14700 15484 14756 15540
rect 14924 16716 14980 16772
rect 15372 17948 15428 18004
rect 16044 21980 16100 22036
rect 16492 31948 16548 32004
rect 17724 33068 17780 33124
rect 17276 31948 17332 32004
rect 17724 32508 17780 32564
rect 18060 32562 18116 32564
rect 18060 32510 18062 32562
rect 18062 32510 18114 32562
rect 18114 32510 18116 32562
rect 18060 32508 18116 32510
rect 18060 31948 18116 32004
rect 16604 31500 16660 31556
rect 17948 31500 18004 31556
rect 16268 29426 16324 29428
rect 16268 29374 16270 29426
rect 16270 29374 16322 29426
rect 16322 29374 16324 29426
rect 16268 29372 16324 29374
rect 16380 29148 16436 29204
rect 16492 29484 16548 29540
rect 16268 28028 16324 28084
rect 16828 29538 16884 29540
rect 16828 29486 16830 29538
rect 16830 29486 16882 29538
rect 16882 29486 16884 29538
rect 16828 29484 16884 29486
rect 17276 29986 17332 29988
rect 17276 29934 17278 29986
rect 17278 29934 17330 29986
rect 17330 29934 17332 29986
rect 17276 29932 17332 29934
rect 16940 28812 16996 28868
rect 17276 29372 17332 29428
rect 16492 27244 16548 27300
rect 16716 27804 16772 27860
rect 16604 27132 16660 27188
rect 16716 27244 16772 27300
rect 16940 28082 16996 28084
rect 16940 28030 16942 28082
rect 16942 28030 16994 28082
rect 16994 28030 16996 28082
rect 16940 28028 16996 28030
rect 17052 27804 17108 27860
rect 16604 26850 16660 26852
rect 16604 26798 16606 26850
rect 16606 26798 16658 26850
rect 16658 26798 16660 26850
rect 16604 26796 16660 26798
rect 16492 26348 16548 26404
rect 16268 25564 16324 25620
rect 16380 24892 16436 24948
rect 17164 27692 17220 27748
rect 17724 30322 17780 30324
rect 17724 30270 17726 30322
rect 17726 30270 17778 30322
rect 17778 30270 17780 30322
rect 17724 30268 17780 30270
rect 17724 28252 17780 28308
rect 17836 29372 17892 29428
rect 17724 27580 17780 27636
rect 18060 29932 18116 29988
rect 18172 28700 18228 28756
rect 18060 28364 18116 28420
rect 18172 27970 18228 27972
rect 18172 27918 18174 27970
rect 18174 27918 18226 27970
rect 18226 27918 18228 27970
rect 18172 27916 18228 27918
rect 17164 26684 17220 26740
rect 17724 27020 17780 27076
rect 16716 26012 16772 26068
rect 16716 25676 16772 25732
rect 16156 21532 16212 21588
rect 16044 21308 16100 21364
rect 15932 19852 15988 19908
rect 15708 18620 15764 18676
rect 15596 18562 15652 18564
rect 15596 18510 15598 18562
rect 15598 18510 15650 18562
rect 15650 18510 15652 18562
rect 15596 18508 15652 18510
rect 15820 19740 15876 19796
rect 15932 19404 15988 19460
rect 16156 19852 16212 19908
rect 16044 19068 16100 19124
rect 16044 18844 16100 18900
rect 15932 18620 15988 18676
rect 15484 16940 15540 16996
rect 15148 15484 15204 15540
rect 14252 14924 14308 14980
rect 15036 15148 15092 15204
rect 13916 12572 13972 12628
rect 13804 11340 13860 11396
rect 14252 13692 14308 13748
rect 14252 12572 14308 12628
rect 14476 14140 14532 14196
rect 14924 14364 14980 14420
rect 14700 13970 14756 13972
rect 14700 13918 14702 13970
rect 14702 13918 14754 13970
rect 14754 13918 14756 13970
rect 14700 13916 14756 13918
rect 14476 13692 14532 13748
rect 14588 13580 14644 13636
rect 14140 11228 14196 11284
rect 15148 13916 15204 13972
rect 15260 14812 15316 14868
rect 15148 13692 15204 13748
rect 14924 12572 14980 12628
rect 13916 10220 13972 10276
rect 14364 11116 14420 11172
rect 14476 11228 14532 11284
rect 14252 9996 14308 10052
rect 14140 9938 14196 9940
rect 14140 9886 14142 9938
rect 14142 9886 14194 9938
rect 14194 9886 14196 9938
rect 14140 9884 14196 9886
rect 13692 9266 13748 9268
rect 13692 9214 13694 9266
rect 13694 9214 13746 9266
rect 13746 9214 13748 9266
rect 13692 9212 13748 9214
rect 13580 8316 13636 8372
rect 13580 8092 13636 8148
rect 14028 9772 14084 9828
rect 14364 9826 14420 9828
rect 14364 9774 14366 9826
rect 14366 9774 14418 9826
rect 14418 9774 14420 9826
rect 14364 9772 14420 9774
rect 14700 10834 14756 10836
rect 14700 10782 14702 10834
rect 14702 10782 14754 10834
rect 14754 10782 14756 10834
rect 14700 10780 14756 10782
rect 14812 11116 14868 11172
rect 14588 10556 14644 10612
rect 14812 10556 14868 10612
rect 15036 13132 15092 13188
rect 15708 17836 15764 17892
rect 16940 25618 16996 25620
rect 16940 25566 16942 25618
rect 16942 25566 16994 25618
rect 16994 25566 16996 25618
rect 16940 25564 16996 25566
rect 17052 25228 17108 25284
rect 16940 24162 16996 24164
rect 16940 24110 16942 24162
rect 16942 24110 16994 24162
rect 16994 24110 16996 24162
rect 16940 24108 16996 24110
rect 17612 26290 17668 26292
rect 17612 26238 17614 26290
rect 17614 26238 17666 26290
rect 17666 26238 17668 26290
rect 17612 26236 17668 26238
rect 17836 26684 17892 26740
rect 17948 25788 18004 25844
rect 17724 25394 17780 25396
rect 17724 25342 17726 25394
rect 17726 25342 17778 25394
rect 17778 25342 17780 25394
rect 17724 25340 17780 25342
rect 18060 25228 18116 25284
rect 18172 27132 18228 27188
rect 17276 24108 17332 24164
rect 17052 23996 17108 24052
rect 17724 23772 17780 23828
rect 16716 23324 16772 23380
rect 17836 23660 17892 23716
rect 16716 23100 16772 23156
rect 16492 23042 16548 23044
rect 16492 22990 16494 23042
rect 16494 22990 16546 23042
rect 16546 22990 16548 23042
rect 16492 22988 16548 22990
rect 16492 22764 16548 22820
rect 16604 22652 16660 22708
rect 17724 22988 17780 23044
rect 16940 22876 16996 22932
rect 17612 22876 17668 22932
rect 17276 22652 17332 22708
rect 16940 22540 16996 22596
rect 16828 21980 16884 22036
rect 16492 20914 16548 20916
rect 16492 20862 16494 20914
rect 16494 20862 16546 20914
rect 16546 20862 16548 20914
rect 16492 20860 16548 20862
rect 16716 19852 16772 19908
rect 16604 19740 16660 19796
rect 17052 21698 17108 21700
rect 17052 21646 17054 21698
rect 17054 21646 17106 21698
rect 17106 21646 17108 21698
rect 17052 21644 17108 21646
rect 16940 21532 16996 21588
rect 17164 19740 17220 19796
rect 16380 17836 16436 17892
rect 16604 18956 16660 19012
rect 16604 18508 16660 18564
rect 16156 16828 16212 16884
rect 16044 16770 16100 16772
rect 16044 16718 16046 16770
rect 16046 16718 16098 16770
rect 16098 16718 16100 16770
rect 16044 16716 16100 16718
rect 16268 16380 16324 16436
rect 16716 18396 16772 18452
rect 17164 18396 17220 18452
rect 17052 18172 17108 18228
rect 17052 17836 17108 17892
rect 16940 17052 16996 17108
rect 16492 16604 16548 16660
rect 15820 16268 15876 16324
rect 16044 15596 16100 15652
rect 16156 16156 16212 16212
rect 16380 15986 16436 15988
rect 16380 15934 16382 15986
rect 16382 15934 16434 15986
rect 16434 15934 16436 15986
rect 16380 15932 16436 15934
rect 16380 15708 16436 15764
rect 16044 15426 16100 15428
rect 16044 15374 16046 15426
rect 16046 15374 16098 15426
rect 16098 15374 16100 15426
rect 16044 15372 16100 15374
rect 16492 15484 16548 15540
rect 15932 15036 15988 15092
rect 16268 15260 16324 15316
rect 16044 14418 16100 14420
rect 16044 14366 16046 14418
rect 16046 14366 16098 14418
rect 16098 14366 16100 14418
rect 16044 14364 16100 14366
rect 15932 14252 15988 14308
rect 15708 13916 15764 13972
rect 16380 13916 16436 13972
rect 15484 13692 15540 13748
rect 15708 13692 15764 13748
rect 15260 13580 15316 13636
rect 15596 13580 15652 13636
rect 15260 13132 15316 13188
rect 15148 12402 15204 12404
rect 15148 12350 15150 12402
rect 15150 12350 15202 12402
rect 15202 12350 15204 12402
rect 15148 12348 15204 12350
rect 15036 12124 15092 12180
rect 15260 11676 15316 11732
rect 15708 12402 15764 12404
rect 15708 12350 15710 12402
rect 15710 12350 15762 12402
rect 15762 12350 15764 12402
rect 15708 12348 15764 12350
rect 15596 11900 15652 11956
rect 16044 12962 16100 12964
rect 16044 12910 16046 12962
rect 16046 12910 16098 12962
rect 16098 12910 16100 12962
rect 16044 12908 16100 12910
rect 16156 12684 16212 12740
rect 16044 12460 16100 12516
rect 16044 12124 16100 12180
rect 15484 11116 15540 11172
rect 14700 9772 14756 9828
rect 14924 9996 14980 10052
rect 14924 9826 14980 9828
rect 14924 9774 14926 9826
rect 14926 9774 14978 9826
rect 14978 9774 14980 9826
rect 14924 9772 14980 9774
rect 15260 9826 15316 9828
rect 15260 9774 15262 9826
rect 15262 9774 15314 9826
rect 15314 9774 15316 9826
rect 15260 9772 15316 9774
rect 13916 8988 13972 9044
rect 14028 7980 14084 8036
rect 13804 7868 13860 7924
rect 13692 7308 13748 7364
rect 13580 6690 13636 6692
rect 13580 6638 13582 6690
rect 13582 6638 13634 6690
rect 13634 6638 13636 6690
rect 13580 6636 13636 6638
rect 13692 6524 13748 6580
rect 14028 6578 14084 6580
rect 14028 6526 14030 6578
rect 14030 6526 14082 6578
rect 14082 6526 14084 6578
rect 14028 6524 14084 6526
rect 12908 5516 12964 5572
rect 13020 4562 13076 4564
rect 13020 4510 13022 4562
rect 13022 4510 13074 4562
rect 13074 4510 13076 4562
rect 13020 4508 13076 4510
rect 13804 4450 13860 4452
rect 13804 4398 13806 4450
rect 13806 4398 13858 4450
rect 13858 4398 13860 4450
rect 13804 4396 13860 4398
rect 12684 4284 12740 4340
rect 13580 3666 13636 3668
rect 13580 3614 13582 3666
rect 13582 3614 13634 3666
rect 13634 3614 13636 3666
rect 13580 3612 13636 3614
rect 12796 3554 12852 3556
rect 12796 3502 12798 3554
rect 12798 3502 12850 3554
rect 12850 3502 12852 3554
rect 12796 3500 12852 3502
rect 11340 3276 11396 3332
rect 8316 1372 8372 1428
rect 14028 6188 14084 6244
rect 14812 9324 14868 9380
rect 14924 9154 14980 9156
rect 14924 9102 14926 9154
rect 14926 9102 14978 9154
rect 14978 9102 14980 9154
rect 14924 9100 14980 9102
rect 14812 8876 14868 8932
rect 14252 7698 14308 7700
rect 14252 7646 14254 7698
rect 14254 7646 14306 7698
rect 14306 7646 14308 7698
rect 14252 7644 14308 7646
rect 14588 7474 14644 7476
rect 14588 7422 14590 7474
rect 14590 7422 14642 7474
rect 14642 7422 14644 7474
rect 14588 7420 14644 7422
rect 14140 5404 14196 5460
rect 14252 6578 14308 6580
rect 14252 6526 14254 6578
rect 14254 6526 14306 6578
rect 14306 6526 14308 6578
rect 14252 6524 14308 6526
rect 15260 9042 15316 9044
rect 15260 8990 15262 9042
rect 15262 8990 15314 9042
rect 15314 8990 15316 9042
rect 15260 8988 15316 8990
rect 15036 7420 15092 7476
rect 15148 6578 15204 6580
rect 15148 6526 15150 6578
rect 15150 6526 15202 6578
rect 15202 6526 15204 6578
rect 15148 6524 15204 6526
rect 14924 6188 14980 6244
rect 15148 6130 15204 6132
rect 15148 6078 15150 6130
rect 15150 6078 15202 6130
rect 15202 6078 15204 6130
rect 15148 6076 15204 6078
rect 14252 5516 14308 5572
rect 14140 4562 14196 4564
rect 14140 4510 14142 4562
rect 14142 4510 14194 4562
rect 14194 4510 14196 4562
rect 14140 4508 14196 4510
rect 14812 5234 14868 5236
rect 14812 5182 14814 5234
rect 14814 5182 14866 5234
rect 14866 5182 14868 5234
rect 14812 5180 14868 5182
rect 14588 4732 14644 4788
rect 14588 4562 14644 4564
rect 14588 4510 14590 4562
rect 14590 4510 14642 4562
rect 14642 4510 14644 4562
rect 14588 4508 14644 4510
rect 15148 4508 15204 4564
rect 15148 4060 15204 4116
rect 15484 6076 15540 6132
rect 15596 10556 15652 10612
rect 15372 4732 15428 4788
rect 16044 10610 16100 10612
rect 16044 10558 16046 10610
rect 16046 10558 16098 10610
rect 16098 10558 16100 10610
rect 16044 10556 16100 10558
rect 16044 10220 16100 10276
rect 16268 12572 16324 12628
rect 17052 16156 17108 16212
rect 17052 15596 17108 15652
rect 17500 21756 17556 21812
rect 17500 21308 17556 21364
rect 17836 22146 17892 22148
rect 17836 22094 17838 22146
rect 17838 22094 17890 22146
rect 17890 22094 17892 22146
rect 17836 22092 17892 22094
rect 18172 24668 18228 24724
rect 18172 24332 18228 24388
rect 18396 35420 18452 35476
rect 18620 37436 18676 37492
rect 18956 37996 19012 38052
rect 18732 37324 18788 37380
rect 18620 37100 18676 37156
rect 19068 37266 19124 37268
rect 19068 37214 19070 37266
rect 19070 37214 19122 37266
rect 19122 37214 19124 37266
rect 19068 37212 19124 37214
rect 18956 35532 19012 35588
rect 18844 35420 18900 35476
rect 18620 33068 18676 33124
rect 18844 34300 18900 34356
rect 18508 31500 18564 31556
rect 18396 30268 18452 30324
rect 18396 29986 18452 29988
rect 18396 29934 18398 29986
rect 18398 29934 18450 29986
rect 18450 29934 18452 29986
rect 18396 29932 18452 29934
rect 19292 35586 19348 35588
rect 19292 35534 19294 35586
rect 19294 35534 19346 35586
rect 19346 35534 19348 35586
rect 19292 35532 19348 35534
rect 19180 34300 19236 34356
rect 19292 34690 19348 34692
rect 19292 34638 19294 34690
rect 19294 34638 19346 34690
rect 19346 34638 19348 34690
rect 19292 34636 19348 34638
rect 19292 33740 19348 33796
rect 19180 33122 19236 33124
rect 19180 33070 19182 33122
rect 19182 33070 19234 33122
rect 19234 33070 19236 33122
rect 19180 33068 19236 33070
rect 20412 38946 20468 38948
rect 20412 38894 20414 38946
rect 20414 38894 20466 38946
rect 20466 38894 20468 38946
rect 20412 38892 20468 38894
rect 19852 38556 19908 38612
rect 19740 38444 19796 38500
rect 19516 38332 19572 38388
rect 20076 37772 20132 37828
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19964 37266 20020 37268
rect 19964 37214 19966 37266
rect 19966 37214 20018 37266
rect 20018 37214 20020 37266
rect 19964 37212 20020 37214
rect 20524 36540 20580 36596
rect 20412 36370 20468 36372
rect 20412 36318 20414 36370
rect 20414 36318 20466 36370
rect 20466 36318 20468 36370
rect 20412 36316 20468 36318
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20300 35308 20356 35364
rect 20412 35084 20468 35140
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19740 33740 19796 33796
rect 20524 34748 20580 34804
rect 20860 40962 20916 40964
rect 20860 40910 20862 40962
rect 20862 40910 20914 40962
rect 20914 40910 20916 40962
rect 20860 40908 20916 40910
rect 20860 40348 20916 40404
rect 20972 39676 21028 39732
rect 21084 39564 21140 39620
rect 20860 38946 20916 38948
rect 20860 38894 20862 38946
rect 20862 38894 20914 38946
rect 20914 38894 20916 38946
rect 20860 38892 20916 38894
rect 20860 38332 20916 38388
rect 20860 37884 20916 37940
rect 21084 39116 21140 39172
rect 21308 42476 21364 42532
rect 21644 40908 21700 40964
rect 21308 39340 21364 39396
rect 20860 36988 20916 37044
rect 20748 36652 20804 36708
rect 20860 35308 20916 35364
rect 21532 39340 21588 39396
rect 22204 40962 22260 40964
rect 22204 40910 22206 40962
rect 22206 40910 22258 40962
rect 22258 40910 22260 40962
rect 22204 40908 22260 40910
rect 21868 40348 21924 40404
rect 21756 39116 21812 39172
rect 21868 40012 21924 40068
rect 21756 38946 21812 38948
rect 21756 38894 21758 38946
rect 21758 38894 21810 38946
rect 21810 38894 21812 38946
rect 21756 38892 21812 38894
rect 21196 38610 21252 38612
rect 21196 38558 21198 38610
rect 21198 38558 21250 38610
rect 21250 38558 21252 38610
rect 21196 38556 21252 38558
rect 21532 37826 21588 37828
rect 21532 37774 21534 37826
rect 21534 37774 21586 37826
rect 21586 37774 21588 37826
rect 21532 37772 21588 37774
rect 21532 37324 21588 37380
rect 22092 39730 22148 39732
rect 22092 39678 22094 39730
rect 22094 39678 22146 39730
rect 22146 39678 22148 39730
rect 22092 39676 22148 39678
rect 22204 39394 22260 39396
rect 22204 39342 22206 39394
rect 22206 39342 22258 39394
rect 22258 39342 22260 39394
rect 22204 39340 22260 39342
rect 22204 38722 22260 38724
rect 22204 38670 22206 38722
rect 22206 38670 22258 38722
rect 22258 38670 22260 38722
rect 22204 38668 22260 38670
rect 23100 43538 23156 43540
rect 23100 43486 23102 43538
rect 23102 43486 23154 43538
rect 23154 43486 23156 43538
rect 23100 43484 23156 43486
rect 23884 43260 23940 43316
rect 23324 42866 23380 42868
rect 23324 42814 23326 42866
rect 23326 42814 23378 42866
rect 23378 42814 23380 42866
rect 23324 42812 23380 42814
rect 22876 42140 22932 42196
rect 23324 42028 23380 42084
rect 22988 40962 23044 40964
rect 22988 40910 22990 40962
rect 22990 40910 23042 40962
rect 23042 40910 23044 40962
rect 22988 40908 23044 40910
rect 24108 42812 24164 42868
rect 23548 40348 23604 40404
rect 22652 39340 22708 39396
rect 22764 40236 22820 40292
rect 21980 38332 22036 38388
rect 23212 39394 23268 39396
rect 23212 39342 23214 39394
rect 23214 39342 23266 39394
rect 23266 39342 23268 39394
rect 23212 39340 23268 39342
rect 22988 38946 23044 38948
rect 22988 38894 22990 38946
rect 22990 38894 23042 38946
rect 23042 38894 23044 38946
rect 22988 38892 23044 38894
rect 22204 37772 22260 37828
rect 21756 36988 21812 37044
rect 21084 34860 21140 34916
rect 21644 36370 21700 36372
rect 21644 36318 21646 36370
rect 21646 36318 21698 36370
rect 21698 36318 21700 36370
rect 21644 36316 21700 36318
rect 21868 35084 21924 35140
rect 21980 34802 22036 34804
rect 21980 34750 21982 34802
rect 21982 34750 22034 34802
rect 22034 34750 22036 34802
rect 21980 34748 22036 34750
rect 21420 34636 21476 34692
rect 21644 34690 21700 34692
rect 21644 34638 21646 34690
rect 21646 34638 21698 34690
rect 21698 34638 21700 34690
rect 21644 34636 21700 34638
rect 21420 34300 21476 34356
rect 19404 31836 19460 31892
rect 19404 31612 19460 31668
rect 19404 31106 19460 31108
rect 19404 31054 19406 31106
rect 19406 31054 19458 31106
rect 19458 31054 19460 31106
rect 19404 31052 19460 31054
rect 19516 30940 19572 30996
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 20636 32674 20692 32676
rect 20636 32622 20638 32674
rect 20638 32622 20690 32674
rect 20690 32622 20692 32674
rect 20636 32620 20692 32622
rect 20860 32620 20916 32676
rect 20524 32562 20580 32564
rect 20524 32510 20526 32562
rect 20526 32510 20578 32562
rect 20578 32510 20580 32562
rect 20524 32508 20580 32510
rect 19628 31948 19684 32004
rect 20188 31890 20244 31892
rect 20188 31838 20190 31890
rect 20190 31838 20242 31890
rect 20242 31838 20244 31890
rect 20188 31836 20244 31838
rect 20076 31666 20132 31668
rect 20076 31614 20078 31666
rect 20078 31614 20130 31666
rect 20130 31614 20132 31666
rect 20076 31612 20132 31614
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19964 31052 20020 31108
rect 19628 30716 19684 30772
rect 19852 30994 19908 30996
rect 19852 30942 19854 30994
rect 19854 30942 19906 30994
rect 19906 30942 19908 30994
rect 19852 30940 19908 30942
rect 18956 30268 19012 30324
rect 18732 30098 18788 30100
rect 18732 30046 18734 30098
rect 18734 30046 18786 30098
rect 18786 30046 18788 30098
rect 18732 30044 18788 30046
rect 18620 29426 18676 29428
rect 18620 29374 18622 29426
rect 18622 29374 18674 29426
rect 18674 29374 18676 29426
rect 18620 29372 18676 29374
rect 18508 28642 18564 28644
rect 18508 28590 18510 28642
rect 18510 28590 18562 28642
rect 18562 28590 18564 28642
rect 18508 28588 18564 28590
rect 18396 28028 18452 28084
rect 18844 28252 18900 28308
rect 19292 28252 19348 28308
rect 18620 27858 18676 27860
rect 18620 27806 18622 27858
rect 18622 27806 18674 27858
rect 18674 27806 18676 27858
rect 18620 27804 18676 27806
rect 19292 27804 19348 27860
rect 19180 27580 19236 27636
rect 18508 27244 18564 27300
rect 18844 27356 18900 27412
rect 18508 27074 18564 27076
rect 18508 27022 18510 27074
rect 18510 27022 18562 27074
rect 18562 27022 18564 27074
rect 18508 27020 18564 27022
rect 19292 26962 19348 26964
rect 19292 26910 19294 26962
rect 19294 26910 19346 26962
rect 19346 26910 19348 26962
rect 19292 26908 19348 26910
rect 18620 26796 18676 26852
rect 18508 26066 18564 26068
rect 18508 26014 18510 26066
rect 18510 26014 18562 26066
rect 18562 26014 18564 26066
rect 18508 26012 18564 26014
rect 18396 24668 18452 24724
rect 18060 23826 18116 23828
rect 18060 23774 18062 23826
rect 18062 23774 18114 23826
rect 18114 23774 18116 23826
rect 18060 23772 18116 23774
rect 18060 23266 18116 23268
rect 18060 23214 18062 23266
rect 18062 23214 18114 23266
rect 18114 23214 18116 23266
rect 18060 23212 18116 23214
rect 18396 23996 18452 24052
rect 18508 24108 18564 24164
rect 18172 21756 18228 21812
rect 17724 20860 17780 20916
rect 18060 21698 18116 21700
rect 18060 21646 18062 21698
rect 18062 21646 18114 21698
rect 18114 21646 18116 21698
rect 18060 21644 18116 21646
rect 18060 21308 18116 21364
rect 18508 22988 18564 23044
rect 19740 30268 19796 30324
rect 19964 30268 20020 30324
rect 20076 30940 20132 30996
rect 20300 30268 20356 30324
rect 20860 30268 20916 30324
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19628 29426 19684 29428
rect 19628 29374 19630 29426
rect 19630 29374 19682 29426
rect 19682 29374 19684 29426
rect 19628 29372 19684 29374
rect 20972 29650 21028 29652
rect 20972 29598 20974 29650
rect 20974 29598 21026 29650
rect 21026 29598 21028 29650
rect 20972 29596 21028 29598
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19740 27858 19796 27860
rect 19740 27806 19742 27858
rect 19742 27806 19794 27858
rect 19794 27806 19796 27858
rect 19740 27804 19796 27806
rect 20412 29426 20468 29428
rect 20412 29374 20414 29426
rect 20414 29374 20466 29426
rect 20466 29374 20468 29426
rect 20412 29372 20468 29374
rect 20748 29372 20804 29428
rect 20188 27356 20244 27412
rect 20188 27132 20244 27188
rect 20636 28028 20692 28084
rect 20972 28642 21028 28644
rect 20972 28590 20974 28642
rect 20974 28590 21026 28642
rect 21026 28590 21028 28642
rect 20972 28588 21028 28590
rect 21308 32284 21364 32340
rect 21196 29372 21252 29428
rect 21756 34130 21812 34132
rect 21756 34078 21758 34130
rect 21758 34078 21810 34130
rect 21810 34078 21812 34130
rect 21756 34076 21812 34078
rect 21532 32620 21588 32676
rect 22092 33180 22148 33236
rect 21756 32620 21812 32676
rect 21756 31836 21812 31892
rect 21644 31276 21700 31332
rect 21868 31778 21924 31780
rect 21868 31726 21870 31778
rect 21870 31726 21922 31778
rect 21922 31726 21924 31778
rect 21868 31724 21924 31726
rect 22204 32172 22260 32228
rect 23212 38162 23268 38164
rect 23212 38110 23214 38162
rect 23214 38110 23266 38162
rect 23266 38110 23268 38162
rect 23212 38108 23268 38110
rect 22652 37378 22708 37380
rect 22652 37326 22654 37378
rect 22654 37326 22706 37378
rect 22706 37326 22708 37378
rect 22652 37324 22708 37326
rect 23436 37324 23492 37380
rect 23212 34914 23268 34916
rect 23212 34862 23214 34914
rect 23214 34862 23266 34914
rect 23266 34862 23268 34914
rect 23212 34860 23268 34862
rect 22428 34802 22484 34804
rect 22428 34750 22430 34802
rect 22430 34750 22482 34802
rect 22482 34750 22484 34802
rect 22428 34748 22484 34750
rect 23772 38556 23828 38612
rect 23996 38108 24052 38164
rect 24556 43484 24612 43540
rect 24332 42140 24388 42196
rect 25116 44044 25172 44100
rect 25004 42812 25060 42868
rect 26460 50876 26516 50932
rect 26348 50594 26404 50596
rect 26348 50542 26350 50594
rect 26350 50542 26402 50594
rect 26402 50542 26404 50594
rect 26348 50540 26404 50542
rect 26124 50428 26180 50484
rect 28028 53228 28084 53284
rect 31052 55468 31108 55524
rect 43036 57036 43092 57092
rect 43596 57036 43652 57092
rect 29596 53228 29652 53284
rect 26796 50876 26852 50932
rect 27468 50876 27524 50932
rect 26124 49756 26180 49812
rect 25228 42140 25284 42196
rect 25340 48076 25396 48132
rect 25004 41186 25060 41188
rect 25004 41134 25006 41186
rect 25006 41134 25058 41186
rect 25058 41134 25060 41186
rect 25004 41132 25060 41134
rect 26124 47964 26180 48020
rect 25564 47740 25620 47796
rect 25452 46620 25508 46676
rect 26796 49922 26852 49924
rect 26796 49870 26798 49922
rect 26798 49870 26850 49922
rect 26850 49870 26852 49922
rect 26796 49868 26852 49870
rect 26572 49810 26628 49812
rect 26572 49758 26574 49810
rect 26574 49758 26626 49810
rect 26626 49758 26628 49810
rect 26572 49756 26628 49758
rect 26684 49644 26740 49700
rect 26796 49138 26852 49140
rect 26796 49086 26798 49138
rect 26798 49086 26850 49138
rect 26850 49086 26852 49138
rect 26796 49084 26852 49086
rect 27020 49868 27076 49924
rect 29036 51212 29092 51268
rect 28252 51100 28308 51156
rect 28140 49922 28196 49924
rect 28140 49870 28142 49922
rect 28142 49870 28194 49922
rect 28194 49870 28196 49922
rect 28140 49868 28196 49870
rect 29484 50652 29540 50708
rect 27692 49644 27748 49700
rect 26908 48748 26964 48804
rect 27132 48354 27188 48356
rect 27132 48302 27134 48354
rect 27134 48302 27186 48354
rect 27186 48302 27188 48354
rect 27132 48300 27188 48302
rect 27916 49084 27972 49140
rect 26684 47404 26740 47460
rect 27468 48018 27524 48020
rect 27468 47966 27470 48018
rect 27470 47966 27522 48018
rect 27522 47966 27524 48018
rect 27468 47964 27524 47966
rect 28476 47180 28532 47236
rect 27244 46674 27300 46676
rect 27244 46622 27246 46674
rect 27246 46622 27298 46674
rect 27298 46622 27300 46674
rect 27244 46620 27300 46622
rect 26124 46508 26180 46564
rect 26124 46002 26180 46004
rect 26124 45950 26126 46002
rect 26126 45950 26178 46002
rect 26178 45950 26180 46002
rect 26124 45948 26180 45950
rect 27020 46002 27076 46004
rect 27020 45950 27022 46002
rect 27022 45950 27074 46002
rect 27074 45950 27076 46002
rect 27020 45948 27076 45950
rect 25564 44434 25620 44436
rect 25564 44382 25566 44434
rect 25566 44382 25618 44434
rect 25618 44382 25620 44434
rect 25564 44380 25620 44382
rect 28252 46172 28308 46228
rect 28476 45890 28532 45892
rect 28476 45838 28478 45890
rect 28478 45838 28530 45890
rect 28530 45838 28532 45890
rect 28476 45836 28532 45838
rect 27356 45388 27412 45444
rect 25900 44268 25956 44324
rect 25788 44044 25844 44100
rect 26124 44380 26180 44436
rect 28700 45612 28756 45668
rect 25676 43538 25732 43540
rect 25676 43486 25678 43538
rect 25678 43486 25730 43538
rect 25730 43486 25732 43538
rect 25676 43484 25732 43486
rect 26348 42866 26404 42868
rect 26348 42814 26350 42866
rect 26350 42814 26402 42866
rect 26402 42814 26404 42866
rect 26348 42812 26404 42814
rect 26908 42812 26964 42868
rect 28476 42924 28532 42980
rect 28140 42754 28196 42756
rect 28140 42702 28142 42754
rect 28142 42702 28194 42754
rect 28194 42702 28196 42754
rect 28140 42700 28196 42702
rect 27244 42364 27300 42420
rect 26012 42194 26068 42196
rect 26012 42142 26014 42194
rect 26014 42142 26066 42194
rect 26066 42142 26068 42194
rect 26012 42140 26068 42142
rect 25900 41692 25956 41748
rect 26012 41356 26068 41412
rect 25900 40908 25956 40964
rect 24332 40402 24388 40404
rect 24332 40350 24334 40402
rect 24334 40350 24386 40402
rect 24386 40350 24388 40402
rect 24332 40348 24388 40350
rect 24668 39340 24724 39396
rect 24332 38780 24388 38836
rect 24444 38556 24500 38612
rect 24780 38556 24836 38612
rect 26348 41020 26404 41076
rect 27244 41410 27300 41412
rect 27244 41358 27246 41410
rect 27246 41358 27298 41410
rect 27298 41358 27300 41410
rect 27244 41356 27300 41358
rect 26684 41132 26740 41188
rect 25788 39394 25844 39396
rect 25788 39342 25790 39394
rect 25790 39342 25842 39394
rect 25842 39342 25844 39394
rect 25788 39340 25844 39342
rect 25340 38220 25396 38276
rect 25452 38556 25508 38612
rect 24556 36370 24612 36372
rect 24556 36318 24558 36370
rect 24558 36318 24610 36370
rect 24610 36318 24612 36370
rect 24556 36316 24612 36318
rect 24108 36204 24164 36260
rect 24108 34972 24164 35028
rect 23772 34914 23828 34916
rect 23772 34862 23774 34914
rect 23774 34862 23826 34914
rect 23826 34862 23828 34914
rect 23772 34860 23828 34862
rect 23660 34748 23716 34804
rect 22540 33458 22596 33460
rect 22540 33406 22542 33458
rect 22542 33406 22594 33458
rect 22594 33406 22596 33458
rect 22540 33404 22596 33406
rect 22988 33068 23044 33124
rect 22876 32956 22932 33012
rect 22652 32284 22708 32340
rect 22540 31836 22596 31892
rect 22428 31724 22484 31780
rect 22204 31276 22260 31332
rect 22092 30492 22148 30548
rect 21980 30268 22036 30324
rect 21868 29650 21924 29652
rect 21868 29598 21870 29650
rect 21870 29598 21922 29650
rect 21922 29598 21924 29650
rect 21868 29596 21924 29598
rect 21532 29314 21588 29316
rect 21532 29262 21534 29314
rect 21534 29262 21586 29314
rect 21586 29262 21588 29314
rect 21532 29260 21588 29262
rect 21868 29036 21924 29092
rect 23100 32284 23156 32340
rect 23100 32060 23156 32116
rect 24668 37996 24724 38052
rect 24780 37324 24836 37380
rect 24332 35026 24388 35028
rect 24332 34974 24334 35026
rect 24334 34974 24386 35026
rect 24386 34974 24388 35026
rect 24332 34972 24388 34974
rect 24780 34748 24836 34804
rect 24892 36092 24948 36148
rect 24892 35756 24948 35812
rect 24332 33516 24388 33572
rect 24556 33964 24612 34020
rect 23884 32956 23940 33012
rect 23212 31724 23268 31780
rect 23772 32562 23828 32564
rect 23772 32510 23774 32562
rect 23774 32510 23826 32562
rect 23826 32510 23828 32562
rect 23772 32508 23828 32510
rect 23772 32284 23828 32340
rect 23660 31836 23716 31892
rect 22988 31388 23044 31444
rect 23660 31276 23716 31332
rect 21420 28364 21476 28420
rect 21532 28700 21588 28756
rect 20636 27692 20692 27748
rect 20860 27356 20916 27412
rect 18956 26178 19012 26180
rect 18956 26126 18958 26178
rect 18958 26126 19010 26178
rect 19010 26126 19012 26178
rect 18956 26124 19012 26126
rect 18956 25564 19012 25620
rect 18732 25452 18788 25508
rect 19068 25452 19124 25508
rect 18956 24892 19012 24948
rect 18956 24668 19012 24724
rect 18844 24332 18900 24388
rect 18732 22482 18788 22484
rect 18732 22430 18734 22482
rect 18734 22430 18786 22482
rect 18786 22430 18788 22482
rect 18732 22428 18788 22430
rect 18732 22092 18788 22148
rect 18284 20412 18340 20468
rect 18060 20300 18116 20356
rect 17612 19234 17668 19236
rect 17612 19182 17614 19234
rect 17614 19182 17666 19234
rect 17666 19182 17668 19234
rect 17612 19180 17668 19182
rect 17500 18620 17556 18676
rect 17388 17276 17444 17332
rect 17948 19906 18004 19908
rect 17948 19854 17950 19906
rect 17950 19854 18002 19906
rect 18002 19854 18004 19906
rect 17948 19852 18004 19854
rect 17500 17052 17556 17108
rect 17500 15484 17556 15540
rect 18172 20188 18228 20244
rect 17948 18956 18004 19012
rect 18172 18844 18228 18900
rect 17948 18620 18004 18676
rect 18284 18620 18340 18676
rect 18284 18450 18340 18452
rect 18284 18398 18286 18450
rect 18286 18398 18338 18450
rect 18338 18398 18340 18450
rect 18284 18396 18340 18398
rect 18060 18060 18116 18116
rect 17724 17666 17780 17668
rect 17724 17614 17726 17666
rect 17726 17614 17778 17666
rect 17778 17614 17780 17666
rect 17724 17612 17780 17614
rect 18172 17106 18228 17108
rect 18172 17054 18174 17106
rect 18174 17054 18226 17106
rect 18226 17054 18228 17106
rect 18172 17052 18228 17054
rect 17724 16994 17780 16996
rect 17724 16942 17726 16994
rect 17726 16942 17778 16994
rect 17778 16942 17780 16994
rect 17724 16940 17780 16942
rect 18060 16940 18116 16996
rect 17948 16882 18004 16884
rect 17948 16830 17950 16882
rect 17950 16830 18002 16882
rect 18002 16830 18004 16882
rect 17948 16828 18004 16830
rect 17836 15986 17892 15988
rect 17836 15934 17838 15986
rect 17838 15934 17890 15986
rect 17890 15934 17892 15986
rect 17836 15932 17892 15934
rect 17948 15820 18004 15876
rect 16828 13970 16884 13972
rect 16828 13918 16830 13970
rect 16830 13918 16882 13970
rect 16882 13918 16884 13970
rect 16828 13916 16884 13918
rect 16828 13186 16884 13188
rect 16828 13134 16830 13186
rect 16830 13134 16882 13186
rect 16882 13134 16884 13186
rect 16828 13132 16884 13134
rect 16380 11788 16436 11844
rect 15932 9884 15988 9940
rect 16044 9772 16100 9828
rect 15820 9436 15876 9492
rect 16268 9660 16324 9716
rect 16156 9548 16212 9604
rect 16268 9436 16324 9492
rect 16156 9266 16212 9268
rect 16156 9214 16158 9266
rect 16158 9214 16210 9266
rect 16210 9214 16212 9266
rect 16156 9212 16212 9214
rect 15820 9154 15876 9156
rect 15820 9102 15822 9154
rect 15822 9102 15874 9154
rect 15874 9102 15876 9154
rect 15820 9100 15876 9102
rect 16156 8540 16212 8596
rect 15820 8370 15876 8372
rect 15820 8318 15822 8370
rect 15822 8318 15874 8370
rect 15874 8318 15876 8370
rect 15820 8316 15876 8318
rect 15820 7980 15876 8036
rect 15820 6972 15876 7028
rect 15708 6636 15764 6692
rect 15708 6188 15764 6244
rect 15820 6076 15876 6132
rect 15820 5628 15876 5684
rect 15820 5234 15876 5236
rect 15820 5182 15822 5234
rect 15822 5182 15874 5234
rect 15874 5182 15876 5234
rect 15820 5180 15876 5182
rect 15596 4732 15652 4788
rect 16716 12124 16772 12180
rect 16492 9996 16548 10052
rect 16492 8540 16548 8596
rect 16380 7474 16436 7476
rect 16380 7422 16382 7474
rect 16382 7422 16434 7474
rect 16434 7422 16436 7474
rect 16380 7420 16436 7422
rect 16380 7196 16436 7252
rect 16380 6636 16436 6692
rect 15820 4562 15876 4564
rect 15820 4510 15822 4562
rect 15822 4510 15874 4562
rect 15874 4510 15876 4562
rect 15820 4508 15876 4510
rect 15596 4060 15652 4116
rect 16940 11452 16996 11508
rect 16828 11340 16884 11396
rect 16940 10892 16996 10948
rect 17836 15708 17892 15764
rect 17388 13468 17444 13524
rect 17612 13916 17668 13972
rect 17724 13634 17780 13636
rect 17724 13582 17726 13634
rect 17726 13582 17778 13634
rect 17778 13582 17780 13634
rect 17724 13580 17780 13582
rect 17388 12572 17444 12628
rect 17052 10556 17108 10612
rect 17052 9266 17108 9268
rect 17052 9214 17054 9266
rect 17054 9214 17106 9266
rect 17106 9214 17108 9266
rect 17052 9212 17108 9214
rect 16828 8428 16884 8484
rect 16716 6748 16772 6804
rect 16604 6412 16660 6468
rect 16604 5292 16660 5348
rect 16940 6636 16996 6692
rect 16940 5292 16996 5348
rect 16828 5180 16884 5236
rect 17388 8428 17444 8484
rect 18284 16770 18340 16772
rect 18284 16718 18286 16770
rect 18286 16718 18338 16770
rect 18338 16718 18340 16770
rect 18284 16716 18340 16718
rect 18620 20914 18676 20916
rect 18620 20862 18622 20914
rect 18622 20862 18674 20914
rect 18674 20862 18676 20914
rect 18620 20860 18676 20862
rect 18508 20412 18564 20468
rect 18508 19404 18564 19460
rect 18620 18844 18676 18900
rect 18956 23436 19012 23492
rect 19068 24444 19124 24500
rect 19404 26290 19460 26292
rect 19404 26238 19406 26290
rect 19406 26238 19458 26290
rect 19458 26238 19460 26290
rect 19404 26236 19460 26238
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 20412 26402 20468 26404
rect 20412 26350 20414 26402
rect 20414 26350 20466 26402
rect 20466 26350 20468 26402
rect 20412 26348 20468 26350
rect 20188 26012 20244 26068
rect 19852 25788 19908 25844
rect 19740 25564 19796 25620
rect 19292 25004 19348 25060
rect 19180 24108 19236 24164
rect 19068 23212 19124 23268
rect 19292 23938 19348 23940
rect 19292 23886 19294 23938
rect 19294 23886 19346 23938
rect 19346 23886 19348 23938
rect 19292 23884 19348 23886
rect 18956 22540 19012 22596
rect 19068 22428 19124 22484
rect 20076 25228 20132 25284
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19516 24444 19572 24500
rect 19180 22092 19236 22148
rect 19516 23266 19572 23268
rect 19516 23214 19518 23266
rect 19518 23214 19570 23266
rect 19570 23214 19572 23266
rect 19516 23212 19572 23214
rect 19404 22988 19460 23044
rect 20860 27074 20916 27076
rect 20860 27022 20862 27074
rect 20862 27022 20914 27074
rect 20914 27022 20916 27074
rect 20860 27020 20916 27022
rect 20524 26236 20580 26292
rect 20860 25506 20916 25508
rect 20860 25454 20862 25506
rect 20862 25454 20914 25506
rect 20914 25454 20916 25506
rect 20860 25452 20916 25454
rect 20300 24332 20356 24388
rect 20524 25228 20580 25284
rect 20300 24108 20356 24164
rect 20076 23660 20132 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19404 22428 19460 22484
rect 20076 23324 20132 23380
rect 19068 21474 19124 21476
rect 19068 21422 19070 21474
rect 19070 21422 19122 21474
rect 19122 21422 19124 21474
rect 19068 21420 19124 21422
rect 19628 22204 19684 22260
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 21420 27020 21476 27076
rect 20860 24668 20916 24724
rect 20748 23826 20804 23828
rect 20748 23774 20750 23826
rect 20750 23774 20802 23826
rect 20802 23774 20804 23826
rect 20748 23772 20804 23774
rect 20636 23100 20692 23156
rect 20412 22988 20468 23044
rect 20860 22652 20916 22708
rect 20636 22428 20692 22484
rect 20636 22204 20692 22260
rect 20076 21810 20132 21812
rect 20076 21758 20078 21810
rect 20078 21758 20130 21810
rect 20130 21758 20132 21810
rect 20076 21756 20132 21758
rect 19404 21586 19460 21588
rect 19404 21534 19406 21586
rect 19406 21534 19458 21586
rect 19458 21534 19460 21586
rect 19404 21532 19460 21534
rect 19292 20860 19348 20916
rect 19180 20690 19236 20692
rect 19180 20638 19182 20690
rect 19182 20638 19234 20690
rect 19234 20638 19236 20690
rect 19180 20636 19236 20638
rect 19516 20690 19572 20692
rect 19516 20638 19518 20690
rect 19518 20638 19570 20690
rect 19570 20638 19572 20690
rect 19516 20636 19572 20638
rect 19068 20018 19124 20020
rect 19068 19966 19070 20018
rect 19070 19966 19122 20018
rect 19122 19966 19124 20018
rect 19068 19964 19124 19966
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 21308 23996 21364 24052
rect 21196 22764 21252 22820
rect 21084 22428 21140 22484
rect 20524 21586 20580 21588
rect 20524 21534 20526 21586
rect 20526 21534 20578 21586
rect 20578 21534 20580 21586
rect 20524 21532 20580 21534
rect 20748 21196 20804 21252
rect 20636 20914 20692 20916
rect 20636 20862 20638 20914
rect 20638 20862 20690 20914
rect 20690 20862 20692 20914
rect 20636 20860 20692 20862
rect 19740 19628 19796 19684
rect 19404 19516 19460 19572
rect 19404 19292 19460 19348
rect 19628 19346 19684 19348
rect 19628 19294 19630 19346
rect 19630 19294 19682 19346
rect 19682 19294 19684 19346
rect 19628 19292 19684 19294
rect 18844 18060 18900 18116
rect 18844 17052 18900 17108
rect 18844 16882 18900 16884
rect 18844 16830 18846 16882
rect 18846 16830 18898 16882
rect 18898 16830 18900 16882
rect 18844 16828 18900 16830
rect 18284 16156 18340 16212
rect 18396 15932 18452 15988
rect 18284 15708 18340 15764
rect 18172 15538 18228 15540
rect 18172 15486 18174 15538
rect 18174 15486 18226 15538
rect 18226 15486 18228 15538
rect 18172 15484 18228 15486
rect 19404 18450 19460 18452
rect 19404 18398 19406 18450
rect 19406 18398 19458 18450
rect 19458 18398 19460 18450
rect 19404 18396 19460 18398
rect 19292 18284 19348 18340
rect 19180 17554 19236 17556
rect 19180 17502 19182 17554
rect 19182 17502 19234 17554
rect 19234 17502 19236 17554
rect 19180 17500 19236 17502
rect 19292 17052 19348 17108
rect 19628 19068 19684 19124
rect 20524 20300 20580 20356
rect 20748 20412 20804 20468
rect 19852 18956 19908 19012
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19628 18396 19684 18452
rect 19628 17612 19684 17668
rect 19740 17836 19796 17892
rect 20412 18508 20468 18564
rect 20412 17778 20468 17780
rect 20412 17726 20414 17778
rect 20414 17726 20466 17778
rect 20466 17726 20468 17778
rect 20412 17724 20468 17726
rect 20860 19628 20916 19684
rect 21084 19852 21140 19908
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16828 19684 16884
rect 19964 16828 20020 16884
rect 19292 16492 19348 16548
rect 19852 16604 19908 16660
rect 19068 16098 19124 16100
rect 19068 16046 19070 16098
rect 19070 16046 19122 16098
rect 19122 16046 19124 16098
rect 19068 16044 19124 16046
rect 19180 15596 19236 15652
rect 18620 15484 18676 15540
rect 18396 15314 18452 15316
rect 18396 15262 18398 15314
rect 18398 15262 18450 15314
rect 18450 15262 18452 15314
rect 18396 15260 18452 15262
rect 18508 14924 18564 14980
rect 18060 14642 18116 14644
rect 18060 14590 18062 14642
rect 18062 14590 18114 14642
rect 18114 14590 18116 14642
rect 18060 14588 18116 14590
rect 17948 14252 18004 14308
rect 17836 13020 17892 13076
rect 17948 13356 18004 13412
rect 18060 12460 18116 12516
rect 17724 11004 17780 11060
rect 17948 10834 18004 10836
rect 17948 10782 17950 10834
rect 17950 10782 18002 10834
rect 18002 10782 18004 10834
rect 17948 10780 18004 10782
rect 18284 14364 18340 14420
rect 18284 13580 18340 13636
rect 18508 14252 18564 14308
rect 19516 15874 19572 15876
rect 19516 15822 19518 15874
rect 19518 15822 19570 15874
rect 19570 15822 19572 15874
rect 19516 15820 19572 15822
rect 20188 16492 20244 16548
rect 19628 15708 19684 15764
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19516 15372 19572 15428
rect 20188 15372 20244 15428
rect 19292 14924 19348 14980
rect 19068 14642 19124 14644
rect 19068 14590 19070 14642
rect 19070 14590 19122 14642
rect 19122 14590 19124 14642
rect 19068 14588 19124 14590
rect 18956 14306 19012 14308
rect 18956 14254 18958 14306
rect 18958 14254 19010 14306
rect 19010 14254 19012 14306
rect 18956 14252 19012 14254
rect 19180 14306 19236 14308
rect 19180 14254 19182 14306
rect 19182 14254 19234 14306
rect 19234 14254 19236 14306
rect 19180 14252 19236 14254
rect 19068 14140 19124 14196
rect 18732 13858 18788 13860
rect 18732 13806 18734 13858
rect 18734 13806 18786 13858
rect 18786 13806 18788 13858
rect 18732 13804 18788 13806
rect 18732 13132 18788 13188
rect 19852 14700 19908 14756
rect 19740 14476 19796 14532
rect 20636 17276 20692 17332
rect 20748 18172 20804 18228
rect 20860 17442 20916 17444
rect 20860 17390 20862 17442
rect 20862 17390 20914 17442
rect 20914 17390 20916 17442
rect 20860 17388 20916 17390
rect 20524 16098 20580 16100
rect 20524 16046 20526 16098
rect 20526 16046 20578 16098
rect 20578 16046 20580 16098
rect 20524 16044 20580 16046
rect 20524 15484 20580 15540
rect 19964 14476 20020 14532
rect 20300 14418 20356 14420
rect 20300 14366 20302 14418
rect 20302 14366 20354 14418
rect 20354 14366 20356 14418
rect 20300 14364 20356 14366
rect 20076 14252 20132 14308
rect 19628 14140 19684 14196
rect 19836 14138 19892 14140
rect 19516 14028 19572 14084
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19740 13916 19796 13972
rect 19180 13634 19236 13636
rect 19180 13582 19182 13634
rect 19182 13582 19234 13634
rect 19234 13582 19236 13634
rect 19180 13580 19236 13582
rect 18620 12572 18676 12628
rect 18732 12684 18788 12740
rect 18396 11340 18452 11396
rect 18284 10556 18340 10612
rect 17612 8428 17668 8484
rect 17948 8428 18004 8484
rect 17836 8204 17892 8260
rect 17500 7420 17556 7476
rect 17276 6802 17332 6804
rect 17276 6750 17278 6802
rect 17278 6750 17330 6802
rect 17330 6750 17332 6802
rect 17276 6748 17332 6750
rect 16716 4956 16772 5012
rect 17276 4732 17332 4788
rect 16492 4562 16548 4564
rect 16492 4510 16494 4562
rect 16494 4510 16546 4562
rect 16546 4510 16548 4562
rect 16492 4508 16548 4510
rect 16940 4562 16996 4564
rect 16940 4510 16942 4562
rect 16942 4510 16994 4562
rect 16994 4510 16996 4562
rect 16940 4508 16996 4510
rect 16492 4284 16548 4340
rect 16156 4172 16212 4228
rect 15372 3948 15428 4004
rect 17836 7698 17892 7700
rect 17836 7646 17838 7698
rect 17838 7646 17890 7698
rect 17890 7646 17892 7698
rect 17836 7644 17892 7646
rect 18172 7474 18228 7476
rect 18172 7422 18174 7474
rect 18174 7422 18226 7474
rect 18226 7422 18228 7474
rect 18172 7420 18228 7422
rect 18060 6578 18116 6580
rect 18060 6526 18062 6578
rect 18062 6526 18114 6578
rect 18114 6526 18116 6578
rect 18060 6524 18116 6526
rect 18060 6300 18116 6356
rect 17836 5852 17892 5908
rect 17724 4450 17780 4452
rect 17724 4398 17726 4450
rect 17726 4398 17778 4450
rect 17778 4398 17780 4450
rect 17724 4396 17780 4398
rect 18060 5292 18116 5348
rect 19180 12684 19236 12740
rect 20300 13356 20356 13412
rect 20188 13074 20244 13076
rect 20188 13022 20190 13074
rect 20190 13022 20242 13074
rect 20242 13022 20244 13074
rect 20188 13020 20244 13022
rect 19740 12684 19796 12740
rect 19836 12570 19892 12572
rect 19404 12348 19460 12404
rect 19516 12460 19572 12516
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19068 12124 19124 12180
rect 18956 11452 19012 11508
rect 19180 12236 19236 12292
rect 19852 12402 19908 12404
rect 19852 12350 19854 12402
rect 19854 12350 19906 12402
rect 19906 12350 19908 12402
rect 19852 12348 19908 12350
rect 20636 14252 20692 14308
rect 20972 16828 21028 16884
rect 21084 18284 21140 18340
rect 20972 16604 21028 16660
rect 21084 16492 21140 16548
rect 21084 16156 21140 16212
rect 21084 15314 21140 15316
rect 21084 15262 21086 15314
rect 21086 15262 21138 15314
rect 21138 15262 21140 15314
rect 21084 15260 21140 15262
rect 21084 14924 21140 14980
rect 20748 13356 20804 13412
rect 21308 22092 21364 22148
rect 21308 21644 21364 21700
rect 21308 19404 21364 19460
rect 21308 17164 21364 17220
rect 21756 28754 21812 28756
rect 21756 28702 21758 28754
rect 21758 28702 21810 28754
rect 21810 28702 21812 28754
rect 21756 28700 21812 28702
rect 22092 28476 22148 28532
rect 21644 27804 21700 27860
rect 21644 27244 21700 27300
rect 21644 24892 21700 24948
rect 21644 24444 21700 24500
rect 22204 28252 22260 28308
rect 22092 27356 22148 27412
rect 22540 30994 22596 30996
rect 22540 30942 22542 30994
rect 22542 30942 22594 30994
rect 22594 30942 22596 30994
rect 22540 30940 22596 30942
rect 22540 30716 22596 30772
rect 22428 29314 22484 29316
rect 22428 29262 22430 29314
rect 22430 29262 22482 29314
rect 22482 29262 22484 29314
rect 22428 29260 22484 29262
rect 22764 30492 22820 30548
rect 23212 30268 23268 30324
rect 24220 32620 24276 32676
rect 23884 31276 23940 31332
rect 23996 31724 24052 31780
rect 21868 25282 21924 25284
rect 21868 25230 21870 25282
rect 21870 25230 21922 25282
rect 21922 25230 21924 25282
rect 21868 25228 21924 25230
rect 21980 25116 22036 25172
rect 21756 23436 21812 23492
rect 21644 22482 21700 22484
rect 21644 22430 21646 22482
rect 21646 22430 21698 22482
rect 21698 22430 21700 22482
rect 21644 22428 21700 22430
rect 22764 29314 22820 29316
rect 22764 29262 22766 29314
rect 22766 29262 22818 29314
rect 22818 29262 22820 29314
rect 22764 29260 22820 29262
rect 22652 28812 22708 28868
rect 23100 28642 23156 28644
rect 23100 28590 23102 28642
rect 23102 28590 23154 28642
rect 23154 28590 23156 28642
rect 23100 28588 23156 28590
rect 22540 28476 22596 28532
rect 22764 27916 22820 27972
rect 23100 27580 23156 27636
rect 22652 27244 22708 27300
rect 22652 26290 22708 26292
rect 22652 26238 22654 26290
rect 22654 26238 22706 26290
rect 22706 26238 22708 26290
rect 22652 26236 22708 26238
rect 22652 25676 22708 25732
rect 22540 25564 22596 25620
rect 23548 29596 23604 29652
rect 23660 29372 23716 29428
rect 24220 31276 24276 31332
rect 24444 33234 24500 33236
rect 24444 33182 24446 33234
rect 24446 33182 24498 33234
rect 24498 33182 24500 33234
rect 24444 33180 24500 33182
rect 24444 31836 24500 31892
rect 24780 32284 24836 32340
rect 24668 31778 24724 31780
rect 24668 31726 24670 31778
rect 24670 31726 24722 31778
rect 24722 31726 24724 31778
rect 24668 31724 24724 31726
rect 24556 30994 24612 30996
rect 24556 30942 24558 30994
rect 24558 30942 24610 30994
rect 24610 30942 24612 30994
rect 24556 30940 24612 30942
rect 24444 30210 24500 30212
rect 24444 30158 24446 30210
rect 24446 30158 24498 30210
rect 24498 30158 24500 30210
rect 24444 30156 24500 30158
rect 24780 31276 24836 31332
rect 24892 31106 24948 31108
rect 24892 31054 24894 31106
rect 24894 31054 24946 31106
rect 24946 31054 24948 31106
rect 24892 31052 24948 31054
rect 24780 30156 24836 30212
rect 24332 29426 24388 29428
rect 24332 29374 24334 29426
rect 24334 29374 24386 29426
rect 24386 29374 24388 29426
rect 24332 29372 24388 29374
rect 24108 29314 24164 29316
rect 24108 29262 24110 29314
rect 24110 29262 24162 29314
rect 24162 29262 24164 29314
rect 24108 29260 24164 29262
rect 23660 28812 23716 28868
rect 23324 26908 23380 26964
rect 23772 28754 23828 28756
rect 23772 28702 23774 28754
rect 23774 28702 23826 28754
rect 23826 28702 23828 28754
rect 23772 28700 23828 28702
rect 23660 28252 23716 28308
rect 23436 26348 23492 26404
rect 23212 25564 23268 25620
rect 22316 23212 22372 23268
rect 22204 22988 22260 23044
rect 21868 22316 21924 22372
rect 21756 22204 21812 22260
rect 21980 22092 22036 22148
rect 21868 21980 21924 22036
rect 21644 21644 21700 21700
rect 21532 20636 21588 20692
rect 21756 21420 21812 21476
rect 21644 20524 21700 20580
rect 21756 20300 21812 20356
rect 22092 21698 22148 21700
rect 22092 21646 22094 21698
rect 22094 21646 22146 21698
rect 22146 21646 22148 21698
rect 22092 21644 22148 21646
rect 22316 21698 22372 21700
rect 22316 21646 22318 21698
rect 22318 21646 22370 21698
rect 22370 21646 22372 21698
rect 22316 21644 22372 21646
rect 22316 21084 22372 21140
rect 21868 20076 21924 20132
rect 21868 19628 21924 19684
rect 21980 19852 22036 19908
rect 21532 18172 21588 18228
rect 21756 19010 21812 19012
rect 21756 18958 21758 19010
rect 21758 18958 21810 19010
rect 21810 18958 21812 19010
rect 21756 18956 21812 18958
rect 21980 18674 22036 18676
rect 21980 18622 21982 18674
rect 21982 18622 22034 18674
rect 22034 18622 22036 18674
rect 21980 18620 22036 18622
rect 21868 18284 21924 18340
rect 21980 18396 22036 18452
rect 21756 17724 21812 17780
rect 22092 18226 22148 18228
rect 22092 18174 22094 18226
rect 22094 18174 22146 18226
rect 22146 18174 22148 18226
rect 22092 18172 22148 18174
rect 21644 17164 21700 17220
rect 21756 17276 21812 17332
rect 21196 13580 21252 13636
rect 20748 12850 20804 12852
rect 20748 12798 20750 12850
rect 20750 12798 20802 12850
rect 20802 12798 20804 12850
rect 20748 12796 20804 12798
rect 19180 11228 19236 11284
rect 19180 10610 19236 10612
rect 19180 10558 19182 10610
rect 19182 10558 19234 10610
rect 19234 10558 19236 10610
rect 19180 10556 19236 10558
rect 19068 10108 19124 10164
rect 18956 9826 19012 9828
rect 18956 9774 18958 9826
rect 18958 9774 19010 9826
rect 19010 9774 19012 9826
rect 18956 9772 19012 9774
rect 18620 9212 18676 9268
rect 18620 8876 18676 8932
rect 18508 8428 18564 8484
rect 18284 6300 18340 6356
rect 18396 6860 18452 6916
rect 18284 5740 18340 5796
rect 18172 4508 18228 4564
rect 19852 11788 19908 11844
rect 19628 11394 19684 11396
rect 19628 11342 19630 11394
rect 19630 11342 19682 11394
rect 19682 11342 19684 11394
rect 19628 11340 19684 11342
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19852 10332 19908 10388
rect 19964 9884 20020 9940
rect 19964 9548 20020 9604
rect 20412 10722 20468 10724
rect 20412 10670 20414 10722
rect 20414 10670 20466 10722
rect 20466 10670 20468 10722
rect 20412 10668 20468 10670
rect 20300 10610 20356 10612
rect 20300 10558 20302 10610
rect 20302 10558 20354 10610
rect 20354 10558 20356 10610
rect 20300 10556 20356 10558
rect 20188 10498 20244 10500
rect 20188 10446 20190 10498
rect 20190 10446 20242 10498
rect 20242 10446 20244 10498
rect 20188 10444 20244 10446
rect 20860 10668 20916 10724
rect 21420 16770 21476 16772
rect 21420 16718 21422 16770
rect 21422 16718 21474 16770
rect 21474 16718 21476 16770
rect 21420 16716 21476 16718
rect 21420 15484 21476 15540
rect 21868 16492 21924 16548
rect 21756 15986 21812 15988
rect 21756 15934 21758 15986
rect 21758 15934 21810 15986
rect 21810 15934 21812 15986
rect 21756 15932 21812 15934
rect 21644 15484 21700 15540
rect 21868 15260 21924 15316
rect 21644 14700 21700 14756
rect 21532 14588 21588 14644
rect 21532 14252 21588 14308
rect 21308 13020 21364 13076
rect 21532 13244 21588 13300
rect 21644 13020 21700 13076
rect 21420 12684 21476 12740
rect 21196 11676 21252 11732
rect 20972 11564 21028 11620
rect 20636 10556 20692 10612
rect 19628 9436 19684 9492
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19180 8876 19236 8932
rect 19068 8764 19124 8820
rect 19628 8876 19684 8932
rect 18620 7644 18676 7700
rect 18956 8540 19012 8596
rect 18844 7308 18900 7364
rect 18732 7084 18788 7140
rect 18732 6860 18788 6916
rect 19292 8316 19348 8372
rect 18956 6524 19012 6580
rect 17948 3948 18004 4004
rect 16828 3666 16884 3668
rect 16828 3614 16830 3666
rect 16830 3614 16882 3666
rect 16882 3614 16884 3666
rect 16828 3612 16884 3614
rect 18732 3836 18788 3892
rect 19292 7474 19348 7476
rect 19292 7422 19294 7474
rect 19294 7422 19346 7474
rect 19346 7422 19348 7474
rect 19292 7420 19348 7422
rect 19740 8540 19796 8596
rect 19964 9266 20020 9268
rect 19964 9214 19966 9266
rect 19966 9214 20018 9266
rect 20018 9214 20020 9266
rect 19964 9212 20020 9214
rect 19516 8428 19572 8484
rect 19740 8316 19796 8372
rect 20412 8540 20468 8596
rect 19964 8316 20020 8372
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19852 7698 19908 7700
rect 19852 7646 19854 7698
rect 19854 7646 19906 7698
rect 19906 7646 19908 7698
rect 19852 7644 19908 7646
rect 20300 8316 20356 8372
rect 20300 7644 20356 7700
rect 20188 7196 20244 7252
rect 19628 7084 19684 7140
rect 19516 6690 19572 6692
rect 19516 6638 19518 6690
rect 19518 6638 19570 6690
rect 19570 6638 19572 6690
rect 19516 6636 19572 6638
rect 20076 6578 20132 6580
rect 20076 6526 20078 6578
rect 20078 6526 20130 6578
rect 20130 6526 20132 6578
rect 20076 6524 20132 6526
rect 20300 6412 20356 6468
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19628 6076 19684 6132
rect 19628 5516 19684 5572
rect 19292 5068 19348 5124
rect 19964 5234 20020 5236
rect 19964 5182 19966 5234
rect 19966 5182 20018 5234
rect 20018 5182 20020 5234
rect 19964 5180 20020 5182
rect 20300 5068 20356 5124
rect 20748 9884 20804 9940
rect 20748 8930 20804 8932
rect 20748 8878 20750 8930
rect 20750 8878 20802 8930
rect 20802 8878 20804 8930
rect 20748 8876 20804 8878
rect 20860 8316 20916 8372
rect 20860 7196 20916 7252
rect 20636 6130 20692 6132
rect 20636 6078 20638 6130
rect 20638 6078 20690 6130
rect 20690 6078 20692 6130
rect 20636 6076 20692 6078
rect 21308 10444 21364 10500
rect 21532 11340 21588 11396
rect 21532 9324 21588 9380
rect 21084 7644 21140 7700
rect 22092 15932 22148 15988
rect 22316 20188 22372 20244
rect 22764 23042 22820 23044
rect 22764 22990 22766 23042
rect 22766 22990 22818 23042
rect 22818 22990 22820 23042
rect 22764 22988 22820 22990
rect 22876 22370 22932 22372
rect 22876 22318 22878 22370
rect 22878 22318 22930 22370
rect 22930 22318 22932 22370
rect 22876 22316 22932 22318
rect 22652 20860 22708 20916
rect 22764 21532 22820 21588
rect 22876 20524 22932 20580
rect 22428 19516 22484 19572
rect 22316 15596 22372 15652
rect 23324 25900 23380 25956
rect 23212 25394 23268 25396
rect 23212 25342 23214 25394
rect 23214 25342 23266 25394
rect 23266 25342 23268 25394
rect 23212 25340 23268 25342
rect 23100 25116 23156 25172
rect 23100 24780 23156 24836
rect 23212 23938 23268 23940
rect 23212 23886 23214 23938
rect 23214 23886 23266 23938
rect 23266 23886 23268 23938
rect 23212 23884 23268 23886
rect 23212 22988 23268 23044
rect 23100 21026 23156 21028
rect 23100 20974 23102 21026
rect 23102 20974 23154 21026
rect 23154 20974 23156 21026
rect 23100 20972 23156 20974
rect 22652 20076 22708 20132
rect 22764 19794 22820 19796
rect 22764 19742 22766 19794
rect 22766 19742 22818 19794
rect 22818 19742 22820 19794
rect 22764 19740 22820 19742
rect 22988 19516 23044 19572
rect 23100 19010 23156 19012
rect 23100 18958 23102 19010
rect 23102 18958 23154 19010
rect 23154 18958 23156 19010
rect 23100 18956 23156 18958
rect 23436 25506 23492 25508
rect 23436 25454 23438 25506
rect 23438 25454 23490 25506
rect 23490 25454 23492 25506
rect 23436 25452 23492 25454
rect 23548 24668 23604 24724
rect 23660 24444 23716 24500
rect 24108 26796 24164 26852
rect 24108 26460 24164 26516
rect 24332 26348 24388 26404
rect 24556 29372 24612 29428
rect 24780 29372 24836 29428
rect 24892 29260 24948 29316
rect 24668 28588 24724 28644
rect 24556 27858 24612 27860
rect 24556 27806 24558 27858
rect 24558 27806 24610 27858
rect 24610 27806 24612 27858
rect 24556 27804 24612 27806
rect 24220 26012 24276 26068
rect 24220 25282 24276 25284
rect 24220 25230 24222 25282
rect 24222 25230 24274 25282
rect 24274 25230 24276 25282
rect 24220 25228 24276 25230
rect 24332 24834 24388 24836
rect 24332 24782 24334 24834
rect 24334 24782 24386 24834
rect 24386 24782 24388 24834
rect 24332 24780 24388 24782
rect 23548 23772 23604 23828
rect 23324 21868 23380 21924
rect 23436 23212 23492 23268
rect 23772 23826 23828 23828
rect 23772 23774 23774 23826
rect 23774 23774 23826 23826
rect 23826 23774 23828 23826
rect 23772 23772 23828 23774
rect 23660 21980 23716 22036
rect 23324 21586 23380 21588
rect 23324 21534 23326 21586
rect 23326 21534 23378 21586
rect 23378 21534 23380 21586
rect 23324 21532 23380 21534
rect 23324 20636 23380 20692
rect 23660 21698 23716 21700
rect 23660 21646 23662 21698
rect 23662 21646 23714 21698
rect 23714 21646 23716 21698
rect 23660 21644 23716 21646
rect 24332 24444 24388 24500
rect 24108 23884 24164 23940
rect 24220 23042 24276 23044
rect 24220 22990 24222 23042
rect 24222 22990 24274 23042
rect 24274 22990 24276 23042
rect 24220 22988 24276 22990
rect 23884 21756 23940 21812
rect 23884 20300 23940 20356
rect 23772 20130 23828 20132
rect 23772 20078 23774 20130
rect 23774 20078 23826 20130
rect 23826 20078 23828 20130
rect 23772 20076 23828 20078
rect 23548 19740 23604 19796
rect 23324 19234 23380 19236
rect 23324 19182 23326 19234
rect 23326 19182 23378 19234
rect 23378 19182 23380 19234
rect 23324 19180 23380 19182
rect 22988 18284 23044 18340
rect 22764 17836 22820 17892
rect 22540 17442 22596 17444
rect 22540 17390 22542 17442
rect 22542 17390 22594 17442
rect 22594 17390 22596 17442
rect 22540 17388 22596 17390
rect 22652 17724 22708 17780
rect 22428 15538 22484 15540
rect 22428 15486 22430 15538
rect 22430 15486 22482 15538
rect 22482 15486 22484 15538
rect 22428 15484 22484 15486
rect 22204 15148 22260 15204
rect 21980 14812 22036 14868
rect 22092 14252 22148 14308
rect 21980 12908 22036 12964
rect 21868 12290 21924 12292
rect 21868 12238 21870 12290
rect 21870 12238 21922 12290
rect 21922 12238 21924 12290
rect 21868 12236 21924 12238
rect 22428 14364 22484 14420
rect 22652 16940 22708 16996
rect 22428 13692 22484 13748
rect 22540 13356 22596 13412
rect 22428 13244 22484 13300
rect 22204 12290 22260 12292
rect 22204 12238 22206 12290
rect 22206 12238 22258 12290
rect 22258 12238 22260 12290
rect 22204 12236 22260 12238
rect 22092 12124 22148 12180
rect 21980 11900 22036 11956
rect 21756 9772 21812 9828
rect 21868 9212 21924 9268
rect 22092 11676 22148 11732
rect 22092 11170 22148 11172
rect 22092 11118 22094 11170
rect 22094 11118 22146 11170
rect 22146 11118 22148 11170
rect 22092 11116 22148 11118
rect 22204 10780 22260 10836
rect 22092 10610 22148 10612
rect 22092 10558 22094 10610
rect 22094 10558 22146 10610
rect 22146 10558 22148 10610
rect 22092 10556 22148 10558
rect 22316 9436 22372 9492
rect 22652 11116 22708 11172
rect 22540 9826 22596 9828
rect 22540 9774 22542 9826
rect 22542 9774 22594 9826
rect 22594 9774 22596 9826
rect 22540 9772 22596 9774
rect 22540 9266 22596 9268
rect 22540 9214 22542 9266
rect 22542 9214 22594 9266
rect 22594 9214 22596 9266
rect 22540 9212 22596 9214
rect 21980 8540 22036 8596
rect 22092 8316 22148 8372
rect 21420 6076 21476 6132
rect 21532 8204 21588 8260
rect 22204 8092 22260 8148
rect 21868 7420 21924 7476
rect 22204 7420 22260 7476
rect 22316 7084 22372 7140
rect 24108 21868 24164 21924
rect 23548 19346 23604 19348
rect 23548 19294 23550 19346
rect 23550 19294 23602 19346
rect 23602 19294 23604 19346
rect 23548 19292 23604 19294
rect 23436 18620 23492 18676
rect 23996 18732 24052 18788
rect 24444 21756 24500 21812
rect 24444 21586 24500 21588
rect 24444 21534 24446 21586
rect 24446 21534 24498 21586
rect 24498 21534 24500 21586
rect 24444 21532 24500 21534
rect 25116 33516 25172 33572
rect 25340 31948 25396 32004
rect 25116 28924 25172 28980
rect 25004 27692 25060 27748
rect 24780 27244 24836 27300
rect 24892 27132 24948 27188
rect 25116 26460 25172 26516
rect 25228 28364 25284 28420
rect 24892 26236 24948 26292
rect 25340 28140 25396 28196
rect 25340 27692 25396 27748
rect 24892 25676 24948 25732
rect 24892 25228 24948 25284
rect 24780 23938 24836 23940
rect 24780 23886 24782 23938
rect 24782 23886 24834 23938
rect 24834 23886 24836 23938
rect 24780 23884 24836 23886
rect 25228 25228 25284 25284
rect 24892 23100 24948 23156
rect 24892 21474 24948 21476
rect 24892 21422 24894 21474
rect 24894 21422 24946 21474
rect 24946 21422 24948 21474
rect 24892 21420 24948 21422
rect 24668 20636 24724 20692
rect 24444 20188 24500 20244
rect 24332 19964 24388 20020
rect 24332 19516 24388 19572
rect 24332 19180 24388 19236
rect 24220 19010 24276 19012
rect 24220 18958 24222 19010
rect 24222 18958 24274 19010
rect 24274 18958 24276 19010
rect 24220 18956 24276 18958
rect 24220 18562 24276 18564
rect 24220 18510 24222 18562
rect 24222 18510 24274 18562
rect 24274 18510 24276 18562
rect 24220 18508 24276 18510
rect 23772 18396 23828 18452
rect 23436 18284 23492 18340
rect 23324 17836 23380 17892
rect 24892 20300 24948 20356
rect 24556 19740 24612 19796
rect 24668 20076 24724 20132
rect 23436 17724 23492 17780
rect 23884 17836 23940 17892
rect 23324 17666 23380 17668
rect 23324 17614 23326 17666
rect 23326 17614 23378 17666
rect 23378 17614 23380 17666
rect 23324 17612 23380 17614
rect 23212 17554 23268 17556
rect 23212 17502 23214 17554
rect 23214 17502 23266 17554
rect 23266 17502 23268 17554
rect 23212 17500 23268 17502
rect 23324 17388 23380 17444
rect 23212 16380 23268 16436
rect 23660 16828 23716 16884
rect 24444 18172 24500 18228
rect 23436 16658 23492 16660
rect 23436 16606 23438 16658
rect 23438 16606 23490 16658
rect 23490 16606 23492 16658
rect 23436 16604 23492 16606
rect 23996 16492 24052 16548
rect 24556 16492 24612 16548
rect 23324 16044 23380 16100
rect 23548 16044 23604 16100
rect 22988 15932 23044 15988
rect 23324 15708 23380 15764
rect 22988 15538 23044 15540
rect 22988 15486 22990 15538
rect 22990 15486 23042 15538
rect 23042 15486 23044 15538
rect 22988 15484 23044 15486
rect 23324 15148 23380 15204
rect 23884 15372 23940 15428
rect 24220 16268 24276 16324
rect 24556 16098 24612 16100
rect 24556 16046 24558 16098
rect 24558 16046 24610 16098
rect 24610 16046 24612 16098
rect 24556 16044 24612 16046
rect 24220 15708 24276 15764
rect 23660 15148 23716 15204
rect 23100 14642 23156 14644
rect 23100 14590 23102 14642
rect 23102 14590 23154 14642
rect 23154 14590 23156 14642
rect 23100 14588 23156 14590
rect 23212 14306 23268 14308
rect 23212 14254 23214 14306
rect 23214 14254 23266 14306
rect 23266 14254 23268 14306
rect 23212 14252 23268 14254
rect 23324 14140 23380 14196
rect 22988 14028 23044 14084
rect 23436 14028 23492 14084
rect 22876 13244 22932 13300
rect 23436 13244 23492 13300
rect 22988 13132 23044 13188
rect 22876 12236 22932 12292
rect 23100 12684 23156 12740
rect 24556 15538 24612 15540
rect 24556 15486 24558 15538
rect 24558 15486 24610 15538
rect 24610 15486 24612 15538
rect 24556 15484 24612 15486
rect 24780 19292 24836 19348
rect 24892 18732 24948 18788
rect 25116 20636 25172 20692
rect 25004 17500 25060 17556
rect 25116 17612 25172 17668
rect 25116 17388 25172 17444
rect 24780 16716 24836 16772
rect 26348 38668 26404 38724
rect 27804 41186 27860 41188
rect 27804 41134 27806 41186
rect 27806 41134 27858 41186
rect 27858 41134 27860 41186
rect 27804 41132 27860 41134
rect 27356 41074 27412 41076
rect 27356 41022 27358 41074
rect 27358 41022 27410 41074
rect 27410 41022 27412 41074
rect 27356 41020 27412 41022
rect 27244 40962 27300 40964
rect 27244 40910 27246 40962
rect 27246 40910 27298 40962
rect 27298 40910 27300 40962
rect 27244 40908 27300 40910
rect 26796 40572 26852 40628
rect 27468 40402 27524 40404
rect 27468 40350 27470 40402
rect 27470 40350 27522 40402
rect 27522 40350 27524 40402
rect 27468 40348 27524 40350
rect 28364 40402 28420 40404
rect 28364 40350 28366 40402
rect 28366 40350 28418 40402
rect 28418 40350 28420 40402
rect 28364 40348 28420 40350
rect 27692 40290 27748 40292
rect 27692 40238 27694 40290
rect 27694 40238 27746 40290
rect 27746 40238 27748 40290
rect 27692 40236 27748 40238
rect 27916 39340 27972 39396
rect 25900 38220 25956 38276
rect 25900 38050 25956 38052
rect 25900 37998 25902 38050
rect 25902 37998 25954 38050
rect 25954 37998 25956 38050
rect 25900 37996 25956 37998
rect 25788 37378 25844 37380
rect 25788 37326 25790 37378
rect 25790 37326 25842 37378
rect 25842 37326 25844 37378
rect 25788 37324 25844 37326
rect 25676 36258 25732 36260
rect 25676 36206 25678 36258
rect 25678 36206 25730 36258
rect 25730 36206 25732 36258
rect 25676 36204 25732 36206
rect 26012 36258 26068 36260
rect 26012 36206 26014 36258
rect 26014 36206 26066 36258
rect 26066 36206 26068 36258
rect 26012 36204 26068 36206
rect 27020 38722 27076 38724
rect 27020 38670 27022 38722
rect 27022 38670 27074 38722
rect 27074 38670 27076 38722
rect 27020 38668 27076 38670
rect 27804 38556 27860 38612
rect 26908 37996 26964 38052
rect 27356 37490 27412 37492
rect 27356 37438 27358 37490
rect 27358 37438 27410 37490
rect 27410 37438 27412 37490
rect 27356 37436 27412 37438
rect 28140 38892 28196 38948
rect 28028 37378 28084 37380
rect 28028 37326 28030 37378
rect 28030 37326 28082 37378
rect 28082 37326 28084 37378
rect 28028 37324 28084 37326
rect 26684 36204 26740 36260
rect 25564 34860 25620 34916
rect 26348 34242 26404 34244
rect 26348 34190 26350 34242
rect 26350 34190 26402 34242
rect 26402 34190 26404 34242
rect 26348 34188 26404 34190
rect 26124 34076 26180 34132
rect 26012 32956 26068 33012
rect 26124 32562 26180 32564
rect 26124 32510 26126 32562
rect 26126 32510 26178 32562
rect 26178 32510 26180 32562
rect 26124 32508 26180 32510
rect 26012 31948 26068 32004
rect 26572 33292 26628 33348
rect 26572 32956 26628 33012
rect 26796 35868 26852 35924
rect 27356 35756 27412 35812
rect 27468 35644 27524 35700
rect 27020 34242 27076 34244
rect 27020 34190 27022 34242
rect 27022 34190 27074 34242
rect 27074 34190 27076 34242
rect 27020 34188 27076 34190
rect 26908 33570 26964 33572
rect 26908 33518 26910 33570
rect 26910 33518 26962 33570
rect 26962 33518 26964 33570
rect 26908 33516 26964 33518
rect 27020 33404 27076 33460
rect 27356 33458 27412 33460
rect 27356 33406 27358 33458
rect 27358 33406 27410 33458
rect 27410 33406 27412 33458
rect 27356 33404 27412 33406
rect 26236 31106 26292 31108
rect 26236 31054 26238 31106
rect 26238 31054 26290 31106
rect 26290 31054 26292 31106
rect 26236 31052 26292 31054
rect 25564 30994 25620 30996
rect 25564 30942 25566 30994
rect 25566 30942 25618 30994
rect 25618 30942 25620 30994
rect 25564 30940 25620 30942
rect 25900 29596 25956 29652
rect 26236 29650 26292 29652
rect 26236 29598 26238 29650
rect 26238 29598 26290 29650
rect 26290 29598 26292 29650
rect 26236 29596 26292 29598
rect 25564 29426 25620 29428
rect 25564 29374 25566 29426
rect 25566 29374 25618 29426
rect 25618 29374 25620 29426
rect 25564 29372 25620 29374
rect 26012 29426 26068 29428
rect 26012 29374 26014 29426
rect 26014 29374 26066 29426
rect 26066 29374 26068 29426
rect 26012 29372 26068 29374
rect 26348 28530 26404 28532
rect 26348 28478 26350 28530
rect 26350 28478 26402 28530
rect 26402 28478 26404 28530
rect 26348 28476 26404 28478
rect 25900 28418 25956 28420
rect 25900 28366 25902 28418
rect 25902 28366 25954 28418
rect 25954 28366 25956 28418
rect 25900 28364 25956 28366
rect 25900 28140 25956 28196
rect 25452 26908 25508 26964
rect 25676 27356 25732 27412
rect 26460 28364 26516 28420
rect 26460 27580 26516 27636
rect 25900 27020 25956 27076
rect 25788 26796 25844 26852
rect 25676 26290 25732 26292
rect 25676 26238 25678 26290
rect 25678 26238 25730 26290
rect 25730 26238 25732 26290
rect 25676 26236 25732 26238
rect 25564 25394 25620 25396
rect 25564 25342 25566 25394
rect 25566 25342 25618 25394
rect 25618 25342 25620 25394
rect 25564 25340 25620 25342
rect 25340 24220 25396 24276
rect 25564 24780 25620 24836
rect 26124 27132 26180 27188
rect 27356 32620 27412 32676
rect 26796 32562 26852 32564
rect 26796 32510 26798 32562
rect 26798 32510 26850 32562
rect 26850 32510 26852 32562
rect 26796 32508 26852 32510
rect 26684 31948 26740 32004
rect 27020 31388 27076 31444
rect 26796 30828 26852 30884
rect 26684 29426 26740 29428
rect 26684 29374 26686 29426
rect 26686 29374 26738 29426
rect 26738 29374 26740 29426
rect 26684 29372 26740 29374
rect 26684 28642 26740 28644
rect 26684 28590 26686 28642
rect 26686 28590 26738 28642
rect 26738 28590 26740 28642
rect 26684 28588 26740 28590
rect 26460 27020 26516 27076
rect 26572 26962 26628 26964
rect 26572 26910 26574 26962
rect 26574 26910 26626 26962
rect 26626 26910 26628 26962
rect 26572 26908 26628 26910
rect 25900 25676 25956 25732
rect 26012 25394 26068 25396
rect 26012 25342 26014 25394
rect 26014 25342 26066 25394
rect 26066 25342 26068 25394
rect 26012 25340 26068 25342
rect 26012 24834 26068 24836
rect 26012 24782 26014 24834
rect 26014 24782 26066 24834
rect 26066 24782 26068 24834
rect 26012 24780 26068 24782
rect 26236 26348 26292 26404
rect 26236 26124 26292 26180
rect 26348 26236 26404 26292
rect 26124 24444 26180 24500
rect 26236 25564 26292 25620
rect 25788 24220 25844 24276
rect 25788 23884 25844 23940
rect 25340 23772 25396 23828
rect 25676 23436 25732 23492
rect 25788 23324 25844 23380
rect 25788 22930 25844 22932
rect 25788 22878 25790 22930
rect 25790 22878 25842 22930
rect 25842 22878 25844 22930
rect 25788 22876 25844 22878
rect 25564 22764 25620 22820
rect 25340 20914 25396 20916
rect 25340 20862 25342 20914
rect 25342 20862 25394 20914
rect 25394 20862 25396 20914
rect 25340 20860 25396 20862
rect 26124 23772 26180 23828
rect 25900 22204 25956 22260
rect 26012 23548 26068 23604
rect 26236 23660 26292 23716
rect 26124 22540 26180 22596
rect 25676 21980 25732 22036
rect 26012 21810 26068 21812
rect 26012 21758 26014 21810
rect 26014 21758 26066 21810
rect 26066 21758 26068 21810
rect 26012 21756 26068 21758
rect 26012 20412 26068 20468
rect 25900 20300 25956 20356
rect 25788 20188 25844 20244
rect 25564 19964 25620 20020
rect 25452 19740 25508 19796
rect 25340 17948 25396 18004
rect 26012 20188 26068 20244
rect 25900 18732 25956 18788
rect 25676 18338 25732 18340
rect 25676 18286 25678 18338
rect 25678 18286 25730 18338
rect 25730 18286 25732 18338
rect 25676 18284 25732 18286
rect 25564 17106 25620 17108
rect 25564 17054 25566 17106
rect 25566 17054 25618 17106
rect 25618 17054 25620 17106
rect 25564 17052 25620 17054
rect 24780 16492 24836 16548
rect 24780 16044 24836 16100
rect 24780 15820 24836 15876
rect 25004 16492 25060 16548
rect 25116 16098 25172 16100
rect 25116 16046 25118 16098
rect 25118 16046 25170 16098
rect 25170 16046 25172 16098
rect 25116 16044 25172 16046
rect 24892 15314 24948 15316
rect 24892 15262 24894 15314
rect 24894 15262 24946 15314
rect 24946 15262 24948 15314
rect 24892 15260 24948 15262
rect 24332 14306 24388 14308
rect 24332 14254 24334 14306
rect 24334 14254 24386 14306
rect 24386 14254 24388 14306
rect 24332 14252 24388 14254
rect 24332 14028 24388 14084
rect 23212 11394 23268 11396
rect 23212 11342 23214 11394
rect 23214 11342 23266 11394
rect 23266 11342 23268 11394
rect 23212 11340 23268 11342
rect 22764 11004 22820 11060
rect 22428 8876 22484 8932
rect 22764 9996 22820 10052
rect 21756 5964 21812 6020
rect 21644 5794 21700 5796
rect 21644 5742 21646 5794
rect 21646 5742 21698 5794
rect 21698 5742 21700 5794
rect 21644 5740 21700 5742
rect 22316 6748 22372 6804
rect 22092 6636 22148 6692
rect 21868 5180 21924 5236
rect 22092 5404 22148 5460
rect 22764 8428 22820 8484
rect 22540 8034 22596 8036
rect 22540 7982 22542 8034
rect 22542 7982 22594 8034
rect 22594 7982 22596 8034
rect 22540 7980 22596 7982
rect 22540 6636 22596 6692
rect 23100 11004 23156 11060
rect 23212 10892 23268 10948
rect 22988 9100 23044 9156
rect 23324 9996 23380 10052
rect 23100 9884 23156 9940
rect 23660 11676 23716 11732
rect 23548 10332 23604 10388
rect 23100 9436 23156 9492
rect 22988 8540 23044 8596
rect 22876 7532 22932 7588
rect 22764 7308 22820 7364
rect 22876 6748 22932 6804
rect 23212 9100 23268 9156
rect 23100 8146 23156 8148
rect 23100 8094 23102 8146
rect 23102 8094 23154 8146
rect 23154 8094 23156 8146
rect 23100 8092 23156 8094
rect 22764 6524 22820 6580
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 22540 5964 22596 6020
rect 22988 5234 23044 5236
rect 22988 5182 22990 5234
rect 22990 5182 23042 5234
rect 23042 5182 23044 5234
rect 22988 5180 23044 5182
rect 22316 4396 22372 4452
rect 20188 3948 20244 4004
rect 19292 3836 19348 3892
rect 23772 11170 23828 11172
rect 23772 11118 23774 11170
rect 23774 11118 23826 11170
rect 23826 11118 23828 11170
rect 23772 11116 23828 11118
rect 24780 13970 24836 13972
rect 24780 13918 24782 13970
rect 24782 13918 24834 13970
rect 24834 13918 24836 13970
rect 24780 13916 24836 13918
rect 24220 12796 24276 12852
rect 24108 11676 24164 11732
rect 24220 12124 24276 12180
rect 24108 10668 24164 10724
rect 23884 10610 23940 10612
rect 23884 10558 23886 10610
rect 23886 10558 23938 10610
rect 23938 10558 23940 10610
rect 23884 10556 23940 10558
rect 24332 10332 24388 10388
rect 23772 9772 23828 9828
rect 24220 9996 24276 10052
rect 23996 9324 24052 9380
rect 24220 9212 24276 9268
rect 23436 7196 23492 7252
rect 23548 7308 23604 7364
rect 23772 7196 23828 7252
rect 23884 7698 23940 7700
rect 23884 7646 23886 7698
rect 23886 7646 23938 7698
rect 23938 7646 23940 7698
rect 23884 7644 23940 7646
rect 25452 16380 25508 16436
rect 25452 15372 25508 15428
rect 25228 13244 25284 13300
rect 24668 11340 24724 11396
rect 24780 10498 24836 10500
rect 24780 10446 24782 10498
rect 24782 10446 24834 10498
rect 24834 10446 24836 10498
rect 24780 10444 24836 10446
rect 24668 10220 24724 10276
rect 24556 9100 24612 9156
rect 25340 12962 25396 12964
rect 25340 12910 25342 12962
rect 25342 12910 25394 12962
rect 25394 12910 25396 12962
rect 25340 12908 25396 12910
rect 25564 14418 25620 14420
rect 25564 14366 25566 14418
rect 25566 14366 25618 14418
rect 25618 14366 25620 14418
rect 25564 14364 25620 14366
rect 25228 11228 25284 11284
rect 24892 8988 24948 9044
rect 24444 7644 24500 7700
rect 23884 6972 23940 7028
rect 23548 6860 23604 6916
rect 24332 6802 24388 6804
rect 24332 6750 24334 6802
rect 24334 6750 24386 6802
rect 24386 6750 24388 6802
rect 24332 6748 24388 6750
rect 23436 6524 23492 6580
rect 23772 6690 23828 6692
rect 23772 6638 23774 6690
rect 23774 6638 23826 6690
rect 23826 6638 23828 6690
rect 23772 6636 23828 6638
rect 23884 6578 23940 6580
rect 23884 6526 23886 6578
rect 23886 6526 23938 6578
rect 23938 6526 23940 6578
rect 23884 6524 23940 6526
rect 24556 6524 24612 6580
rect 24892 7420 24948 7476
rect 25564 11116 25620 11172
rect 25564 10780 25620 10836
rect 25788 17500 25844 17556
rect 26460 25228 26516 25284
rect 26572 26012 26628 26068
rect 26348 22988 26404 23044
rect 26460 24780 26516 24836
rect 26572 22764 26628 22820
rect 26460 22652 26516 22708
rect 27356 28812 27412 28868
rect 27356 28530 27412 28532
rect 27356 28478 27358 28530
rect 27358 28478 27410 28530
rect 27410 28478 27412 28530
rect 27356 28476 27412 28478
rect 27132 28418 27188 28420
rect 27132 28366 27134 28418
rect 27134 28366 27186 28418
rect 27186 28366 27188 28418
rect 27132 28364 27188 28366
rect 26796 27580 26852 27636
rect 26796 25282 26852 25284
rect 26796 25230 26798 25282
rect 26798 25230 26850 25282
rect 26850 25230 26852 25282
rect 26796 25228 26852 25230
rect 27244 27916 27300 27972
rect 27132 26908 27188 26964
rect 27244 27244 27300 27300
rect 27132 26514 27188 26516
rect 27132 26462 27134 26514
rect 27134 26462 27186 26514
rect 27186 26462 27188 26514
rect 27132 26460 27188 26462
rect 27804 34914 27860 34916
rect 27804 34862 27806 34914
rect 27806 34862 27858 34914
rect 27858 34862 27860 34914
rect 27804 34860 27860 34862
rect 27580 33346 27636 33348
rect 27580 33294 27582 33346
rect 27582 33294 27634 33346
rect 27634 33294 27636 33346
rect 27580 33292 27636 33294
rect 28028 33292 28084 33348
rect 27692 31948 27748 32004
rect 28252 38722 28308 38724
rect 28252 38670 28254 38722
rect 28254 38670 28306 38722
rect 28306 38670 28308 38722
rect 28252 38668 28308 38670
rect 28364 38050 28420 38052
rect 28364 37998 28366 38050
rect 28366 37998 28418 38050
rect 28418 37998 28420 38050
rect 28364 37996 28420 37998
rect 28364 35756 28420 35812
rect 28924 45276 28980 45332
rect 28812 42642 28868 42644
rect 28812 42590 28814 42642
rect 28814 42590 28866 42642
rect 28866 42590 28868 42642
rect 28812 42588 28868 42590
rect 28588 42028 28644 42084
rect 28700 41074 28756 41076
rect 28700 41022 28702 41074
rect 28702 41022 28754 41074
rect 28754 41022 28756 41074
rect 28700 41020 28756 41022
rect 28812 40348 28868 40404
rect 29036 40236 29092 40292
rect 29148 40348 29204 40404
rect 28812 37996 28868 38052
rect 28476 33346 28532 33348
rect 28476 33294 28478 33346
rect 28478 33294 28530 33346
rect 28530 33294 28532 33346
rect 28476 33292 28532 33294
rect 28812 33404 28868 33460
rect 28140 30210 28196 30212
rect 28140 30158 28142 30210
rect 28142 30158 28194 30210
rect 28194 30158 28196 30210
rect 28140 30156 28196 30158
rect 27580 29538 27636 29540
rect 27580 29486 27582 29538
rect 27582 29486 27634 29538
rect 27634 29486 27636 29538
rect 27580 29484 27636 29486
rect 27916 29484 27972 29540
rect 27916 28700 27972 28756
rect 28028 28588 28084 28644
rect 27916 27356 27972 27412
rect 28252 27970 28308 27972
rect 28252 27918 28254 27970
rect 28254 27918 28306 27970
rect 28306 27918 28308 27970
rect 28252 27916 28308 27918
rect 28476 29986 28532 29988
rect 28476 29934 28478 29986
rect 28478 29934 28530 29986
rect 28530 29934 28532 29986
rect 28476 29932 28532 29934
rect 28700 30156 28756 30212
rect 28812 29708 28868 29764
rect 28588 28812 28644 28868
rect 28252 27356 28308 27412
rect 27468 26236 27524 26292
rect 27580 26908 27636 26964
rect 27804 26684 27860 26740
rect 27692 25900 27748 25956
rect 28140 27186 28196 27188
rect 28140 27134 28142 27186
rect 28142 27134 28194 27186
rect 28194 27134 28196 27186
rect 28140 27132 28196 27134
rect 28252 26796 28308 26852
rect 28700 28754 28756 28756
rect 28700 28702 28702 28754
rect 28702 28702 28754 28754
rect 28754 28702 28756 28754
rect 28700 28700 28756 28702
rect 28700 27580 28756 27636
rect 28364 26684 28420 26740
rect 28700 27132 28756 27188
rect 28588 27074 28644 27076
rect 28588 27022 28590 27074
rect 28590 27022 28642 27074
rect 28642 27022 28644 27074
rect 28588 27020 28644 27022
rect 29036 37996 29092 38052
rect 30044 49922 30100 49924
rect 30044 49870 30046 49922
rect 30046 49870 30098 49922
rect 30098 49870 30100 49922
rect 30044 49868 30100 49870
rect 30268 49084 30324 49140
rect 30604 49026 30660 49028
rect 30604 48974 30606 49026
rect 30606 48974 30658 49026
rect 30658 48974 30660 49026
rect 30604 48972 30660 48974
rect 29596 48914 29652 48916
rect 29596 48862 29598 48914
rect 29598 48862 29650 48914
rect 29650 48862 29652 48914
rect 29596 48860 29652 48862
rect 30044 48914 30100 48916
rect 30044 48862 30046 48914
rect 30046 48862 30098 48914
rect 30098 48862 30100 48914
rect 30044 48860 30100 48862
rect 30492 48860 30548 48916
rect 29484 48300 29540 48356
rect 29708 48242 29764 48244
rect 29708 48190 29710 48242
rect 29710 48190 29762 48242
rect 29762 48190 29764 48242
rect 29708 48188 29764 48190
rect 29932 48130 29988 48132
rect 29932 48078 29934 48130
rect 29934 48078 29986 48130
rect 29986 48078 29988 48130
rect 29932 48076 29988 48078
rect 29372 46172 29428 46228
rect 29708 46620 29764 46676
rect 30156 47234 30212 47236
rect 30156 47182 30158 47234
rect 30158 47182 30210 47234
rect 30210 47182 30212 47234
rect 30156 47180 30212 47182
rect 30268 46674 30324 46676
rect 30268 46622 30270 46674
rect 30270 46622 30322 46674
rect 30322 46622 30324 46674
rect 30268 46620 30324 46622
rect 29820 46172 29876 46228
rect 29932 45890 29988 45892
rect 29932 45838 29934 45890
rect 29934 45838 29986 45890
rect 29986 45838 29988 45890
rect 29932 45836 29988 45838
rect 30268 45330 30324 45332
rect 30268 45278 30270 45330
rect 30270 45278 30322 45330
rect 30322 45278 30324 45330
rect 30268 45276 30324 45278
rect 29932 45106 29988 45108
rect 29932 45054 29934 45106
rect 29934 45054 29986 45106
rect 29986 45054 29988 45106
rect 29932 45052 29988 45054
rect 30380 44156 30436 44212
rect 29820 43484 29876 43540
rect 29596 42700 29652 42756
rect 30380 42754 30436 42756
rect 30380 42702 30382 42754
rect 30382 42702 30434 42754
rect 30434 42702 30436 42754
rect 30380 42700 30436 42702
rect 29372 42588 29428 42644
rect 30268 42642 30324 42644
rect 30268 42590 30270 42642
rect 30270 42590 30322 42642
rect 30322 42590 30324 42642
rect 30268 42588 30324 42590
rect 29596 42028 29652 42084
rect 30828 47964 30884 48020
rect 30940 48076 30996 48132
rect 30940 47346 30996 47348
rect 30940 47294 30942 47346
rect 30942 47294 30994 47346
rect 30994 47294 30996 47346
rect 30940 47292 30996 47294
rect 30716 45276 30772 45332
rect 33628 56252 33684 56308
rect 36428 55804 36484 55860
rect 36876 55916 36932 55972
rect 35196 55690 35252 55692
rect 35196 55638 35198 55690
rect 35198 55638 35250 55690
rect 35250 55638 35252 55690
rect 35196 55636 35252 55638
rect 35300 55690 35356 55692
rect 35300 55638 35302 55690
rect 35302 55638 35354 55690
rect 35354 55638 35356 55690
rect 35300 55636 35356 55638
rect 35404 55690 35460 55692
rect 35404 55638 35406 55690
rect 35406 55638 35458 55690
rect 35458 55638 35460 55690
rect 35404 55636 35460 55638
rect 40012 56028 40068 56084
rect 37212 55804 37268 55860
rect 41244 56082 41300 56084
rect 41244 56030 41246 56082
rect 41246 56030 41298 56082
rect 41298 56030 41300 56082
rect 41244 56028 41300 56030
rect 36876 55244 36932 55300
rect 33628 55132 33684 55188
rect 37548 55186 37604 55188
rect 37548 55134 37550 55186
rect 37550 55134 37602 55186
rect 37602 55134 37604 55186
rect 37548 55132 37604 55134
rect 32284 52780 32340 52836
rect 31948 51884 32004 51940
rect 31612 51324 31668 51380
rect 31164 50316 31220 50372
rect 32732 52332 32788 52388
rect 33180 52162 33236 52164
rect 33180 52110 33182 52162
rect 33182 52110 33234 52162
rect 33234 52110 33236 52162
rect 33180 52108 33236 52110
rect 33740 52834 33796 52836
rect 33740 52782 33742 52834
rect 33742 52782 33794 52834
rect 33794 52782 33796 52834
rect 33740 52780 33796 52782
rect 33852 52220 33908 52276
rect 33964 52108 34020 52164
rect 34300 52668 34356 52724
rect 33628 51996 33684 52052
rect 32396 51378 32452 51380
rect 32396 51326 32398 51378
rect 32398 51326 32450 51378
rect 32450 51326 32452 51378
rect 32396 51324 32452 51326
rect 31836 50370 31892 50372
rect 31836 50318 31838 50370
rect 31838 50318 31890 50370
rect 31890 50318 31892 50370
rect 31836 50316 31892 50318
rect 32172 49644 32228 49700
rect 31276 49138 31332 49140
rect 31276 49086 31278 49138
rect 31278 49086 31330 49138
rect 31330 49086 31332 49138
rect 31276 49084 31332 49086
rect 31500 49084 31556 49140
rect 31276 48860 31332 48916
rect 31164 48188 31220 48244
rect 31388 48802 31444 48804
rect 31388 48750 31390 48802
rect 31390 48750 31442 48802
rect 31442 48750 31444 48802
rect 31388 48748 31444 48750
rect 31612 48914 31668 48916
rect 31612 48862 31614 48914
rect 31614 48862 31666 48914
rect 31666 48862 31668 48914
rect 31612 48860 31668 48862
rect 32172 48748 32228 48804
rect 32172 48076 32228 48132
rect 32060 47628 32116 47684
rect 31836 46060 31892 46116
rect 31724 45106 31780 45108
rect 31724 45054 31726 45106
rect 31726 45054 31778 45106
rect 31778 45054 31780 45106
rect 31724 45052 31780 45054
rect 30604 44044 30660 44100
rect 30380 42028 30436 42084
rect 29932 41074 29988 41076
rect 29932 41022 29934 41074
rect 29934 41022 29986 41074
rect 29986 41022 29988 41074
rect 29932 41020 29988 41022
rect 29708 40460 29764 40516
rect 29596 40236 29652 40292
rect 29484 39228 29540 39284
rect 29708 39394 29764 39396
rect 29708 39342 29710 39394
rect 29710 39342 29762 39394
rect 29762 39342 29764 39394
rect 29708 39340 29764 39342
rect 29484 37154 29540 37156
rect 29484 37102 29486 37154
rect 29486 37102 29538 37154
rect 29538 37102 29540 37154
rect 29484 37100 29540 37102
rect 29484 33516 29540 33572
rect 29708 37826 29764 37828
rect 29708 37774 29710 37826
rect 29710 37774 29762 37826
rect 29762 37774 29764 37826
rect 29708 37772 29764 37774
rect 30156 40348 30212 40404
rect 30492 40402 30548 40404
rect 30492 40350 30494 40402
rect 30494 40350 30546 40402
rect 30546 40350 30548 40402
rect 30492 40348 30548 40350
rect 30044 39228 30100 39284
rect 30268 39116 30324 39172
rect 30044 38780 30100 38836
rect 30380 38834 30436 38836
rect 30380 38782 30382 38834
rect 30382 38782 30434 38834
rect 30434 38782 30436 38834
rect 30380 38780 30436 38782
rect 30604 39228 30660 39284
rect 31164 44156 31220 44212
rect 31052 43260 31108 43316
rect 31276 43538 31332 43540
rect 31276 43486 31278 43538
rect 31278 43486 31330 43538
rect 31330 43486 31332 43538
rect 31276 43484 31332 43486
rect 31500 44044 31556 44100
rect 31948 43372 32004 43428
rect 31276 43148 31332 43204
rect 31052 42700 31108 42756
rect 30940 42588 30996 42644
rect 31164 39228 31220 39284
rect 31724 42754 31780 42756
rect 31724 42702 31726 42754
rect 31726 42702 31778 42754
rect 31778 42702 31780 42754
rect 31724 42700 31780 42702
rect 31388 42476 31444 42532
rect 31612 42140 31668 42196
rect 31836 42028 31892 42084
rect 31500 41074 31556 41076
rect 31500 41022 31502 41074
rect 31502 41022 31554 41074
rect 31554 41022 31556 41074
rect 31500 41020 31556 41022
rect 31388 39452 31444 39508
rect 31612 39506 31668 39508
rect 31612 39454 31614 39506
rect 31614 39454 31666 39506
rect 31666 39454 31668 39506
rect 31612 39452 31668 39454
rect 30156 38050 30212 38052
rect 30156 37998 30158 38050
rect 30158 37998 30210 38050
rect 30210 37998 30212 38050
rect 30156 37996 30212 37998
rect 29932 37436 29988 37492
rect 29708 37266 29764 37268
rect 29708 37214 29710 37266
rect 29710 37214 29762 37266
rect 29762 37214 29764 37266
rect 29708 37212 29764 37214
rect 29708 35420 29764 35476
rect 30044 35308 30100 35364
rect 29708 33458 29764 33460
rect 29708 33406 29710 33458
rect 29710 33406 29762 33458
rect 29762 33406 29764 33458
rect 29708 33404 29764 33406
rect 29596 30098 29652 30100
rect 29596 30046 29598 30098
rect 29598 30046 29650 30098
rect 29650 30046 29652 30098
rect 29596 30044 29652 30046
rect 29484 29650 29540 29652
rect 29484 29598 29486 29650
rect 29486 29598 29538 29650
rect 29538 29598 29540 29650
rect 29484 29596 29540 29598
rect 29372 28476 29428 28532
rect 29260 28252 29316 28308
rect 29708 28812 29764 28868
rect 29596 28364 29652 28420
rect 28700 26460 28756 26516
rect 28252 25900 28308 25956
rect 27356 25228 27412 25284
rect 27244 24834 27300 24836
rect 27244 24782 27246 24834
rect 27246 24782 27298 24834
rect 27298 24782 27300 24834
rect 27244 24780 27300 24782
rect 26796 24050 26852 24052
rect 26796 23998 26798 24050
rect 26798 23998 26850 24050
rect 26850 23998 26852 24050
rect 26796 23996 26852 23998
rect 26908 23772 26964 23828
rect 27020 24332 27076 24388
rect 26796 23660 26852 23716
rect 27244 23826 27300 23828
rect 27244 23774 27246 23826
rect 27246 23774 27298 23826
rect 27298 23774 27300 23826
rect 27244 23772 27300 23774
rect 27244 22540 27300 22596
rect 26460 21756 26516 21812
rect 26684 21698 26740 21700
rect 26684 21646 26686 21698
rect 26686 21646 26738 21698
rect 26738 21646 26740 21698
rect 26684 21644 26740 21646
rect 26572 21586 26628 21588
rect 26572 21534 26574 21586
rect 26574 21534 26626 21586
rect 26626 21534 26628 21586
rect 26572 21532 26628 21534
rect 26908 21474 26964 21476
rect 26908 21422 26910 21474
rect 26910 21422 26962 21474
rect 26962 21422 26964 21474
rect 26908 21420 26964 21422
rect 28252 25116 28308 25172
rect 28252 24722 28308 24724
rect 28252 24670 28254 24722
rect 28254 24670 28306 24722
rect 28306 24670 28308 24722
rect 28252 24668 28308 24670
rect 28476 26236 28532 26292
rect 27804 23660 27860 23716
rect 27916 23324 27972 23380
rect 27804 21868 27860 21924
rect 27804 21698 27860 21700
rect 27804 21646 27806 21698
rect 27806 21646 27858 21698
rect 27858 21646 27860 21698
rect 27804 21644 27860 21646
rect 26460 20914 26516 20916
rect 26460 20862 26462 20914
rect 26462 20862 26514 20914
rect 26514 20862 26516 20914
rect 26460 20860 26516 20862
rect 27244 21308 27300 21364
rect 26796 20412 26852 20468
rect 26236 20018 26292 20020
rect 26236 19966 26238 20018
rect 26238 19966 26290 20018
rect 26290 19966 26292 20018
rect 26236 19964 26292 19966
rect 26460 19628 26516 19684
rect 26572 19292 26628 19348
rect 26348 19234 26404 19236
rect 26348 19182 26350 19234
rect 26350 19182 26402 19234
rect 26402 19182 26404 19234
rect 26348 19180 26404 19182
rect 26460 19010 26516 19012
rect 26460 18958 26462 19010
rect 26462 18958 26514 19010
rect 26514 18958 26516 19010
rect 26460 18956 26516 18958
rect 27132 20076 27188 20132
rect 27580 21586 27636 21588
rect 27580 21534 27582 21586
rect 27582 21534 27634 21586
rect 27634 21534 27636 21586
rect 27580 21532 27636 21534
rect 27692 21308 27748 21364
rect 28252 23660 28308 23716
rect 28588 26124 28644 26180
rect 28588 24892 28644 24948
rect 28924 26460 28980 26516
rect 29036 26178 29092 26180
rect 29036 26126 29038 26178
rect 29038 26126 29090 26178
rect 29090 26126 29092 26178
rect 29036 26124 29092 26126
rect 29484 26402 29540 26404
rect 29484 26350 29486 26402
rect 29486 26350 29538 26402
rect 29538 26350 29540 26402
rect 29484 26348 29540 26350
rect 29260 25228 29316 25284
rect 28924 24892 28980 24948
rect 29372 25116 29428 25172
rect 28812 24556 28868 24612
rect 29148 24668 29204 24724
rect 29260 24556 29316 24612
rect 29484 24780 29540 24836
rect 28700 23826 28756 23828
rect 28700 23774 28702 23826
rect 28702 23774 28754 23826
rect 28754 23774 28756 23826
rect 28700 23772 28756 23774
rect 28252 22540 28308 22596
rect 28140 22428 28196 22484
rect 28812 23324 28868 23380
rect 28028 21474 28084 21476
rect 28028 21422 28030 21474
rect 28030 21422 28082 21474
rect 28082 21422 28084 21474
rect 28028 21420 28084 21422
rect 28252 20860 28308 20916
rect 28140 20802 28196 20804
rect 28140 20750 28142 20802
rect 28142 20750 28194 20802
rect 28194 20750 28196 20802
rect 28140 20748 28196 20750
rect 27468 20524 27524 20580
rect 27692 20524 27748 20580
rect 28140 20412 28196 20468
rect 27580 19516 27636 19572
rect 26796 18956 26852 19012
rect 27132 18956 27188 19012
rect 27020 18732 27076 18788
rect 26236 18674 26292 18676
rect 26236 18622 26238 18674
rect 26238 18622 26290 18674
rect 26290 18622 26292 18674
rect 26236 18620 26292 18622
rect 26348 17612 26404 17668
rect 26236 17554 26292 17556
rect 26236 17502 26238 17554
rect 26238 17502 26290 17554
rect 26290 17502 26292 17554
rect 26236 17500 26292 17502
rect 26572 16994 26628 16996
rect 26572 16942 26574 16994
rect 26574 16942 26626 16994
rect 26626 16942 26628 16994
rect 26572 16940 26628 16942
rect 26572 16658 26628 16660
rect 26572 16606 26574 16658
rect 26574 16606 26626 16658
rect 26626 16606 26628 16658
rect 26572 16604 26628 16606
rect 26572 16098 26628 16100
rect 26572 16046 26574 16098
rect 26574 16046 26626 16098
rect 26626 16046 26628 16098
rect 26572 16044 26628 16046
rect 26012 15986 26068 15988
rect 26012 15934 26014 15986
rect 26014 15934 26066 15986
rect 26066 15934 26068 15986
rect 26012 15932 26068 15934
rect 25900 15260 25956 15316
rect 26684 15708 26740 15764
rect 26572 15260 26628 15316
rect 26348 13244 26404 13300
rect 26572 12684 26628 12740
rect 26124 11618 26180 11620
rect 26124 11566 26126 11618
rect 26126 11566 26178 11618
rect 26178 11566 26180 11618
rect 26124 11564 26180 11566
rect 25788 11394 25844 11396
rect 25788 11342 25790 11394
rect 25790 11342 25842 11394
rect 25842 11342 25844 11394
rect 25788 11340 25844 11342
rect 26124 11116 26180 11172
rect 25676 10556 25732 10612
rect 25788 10834 25844 10836
rect 25788 10782 25790 10834
rect 25790 10782 25842 10834
rect 25842 10782 25844 10834
rect 25788 10780 25844 10782
rect 25340 7980 25396 8036
rect 26124 9996 26180 10052
rect 25900 9826 25956 9828
rect 25900 9774 25902 9826
rect 25902 9774 25954 9826
rect 25954 9774 25956 9826
rect 25900 9772 25956 9774
rect 25788 9042 25844 9044
rect 25788 8990 25790 9042
rect 25790 8990 25842 9042
rect 25842 8990 25844 9042
rect 25788 8988 25844 8990
rect 26012 9042 26068 9044
rect 26012 8990 26014 9042
rect 26014 8990 26066 9042
rect 26066 8990 26068 9042
rect 26012 8988 26068 8990
rect 25452 8316 25508 8372
rect 25564 8146 25620 8148
rect 25564 8094 25566 8146
rect 25566 8094 25618 8146
rect 25618 8094 25620 8146
rect 25564 8092 25620 8094
rect 26124 8092 26180 8148
rect 26124 7868 26180 7924
rect 25452 7420 25508 7476
rect 25676 7420 25732 7476
rect 25228 6860 25284 6916
rect 23436 4956 23492 5012
rect 24332 5516 24388 5572
rect 23772 4956 23828 5012
rect 24108 4956 24164 5012
rect 24668 4956 24724 5012
rect 24892 4956 24948 5012
rect 23212 3724 23268 3780
rect 24332 3724 24388 3780
rect 20188 3500 20244 3556
rect 25788 6860 25844 6916
rect 26124 6578 26180 6580
rect 26124 6526 26126 6578
rect 26126 6526 26178 6578
rect 26178 6526 26180 6578
rect 26124 6524 26180 6526
rect 25228 4844 25284 4900
rect 24892 3612 24948 3668
rect 25340 3724 25396 3780
rect 13916 3164 13972 3220
rect 13916 2828 13972 2884
rect 26684 12572 26740 12628
rect 26684 12012 26740 12068
rect 26348 9772 26404 9828
rect 27020 17276 27076 17332
rect 27020 16940 27076 16996
rect 26908 15932 26964 15988
rect 27020 13244 27076 13300
rect 26908 11340 26964 11396
rect 26460 8988 26516 9044
rect 27020 10892 27076 10948
rect 27692 20076 27748 20132
rect 28140 20018 28196 20020
rect 28140 19966 28142 20018
rect 28142 19966 28194 20018
rect 28194 19966 28196 20018
rect 28140 19964 28196 19966
rect 28364 20188 28420 20244
rect 28476 23100 28532 23156
rect 28700 22540 28756 22596
rect 28588 22370 28644 22372
rect 28588 22318 28590 22370
rect 28590 22318 28642 22370
rect 28642 22318 28644 22370
rect 28588 22316 28644 22318
rect 28476 21756 28532 21812
rect 28252 19852 28308 19908
rect 27692 19122 27748 19124
rect 27692 19070 27694 19122
rect 27694 19070 27746 19122
rect 27746 19070 27748 19122
rect 27692 19068 27748 19070
rect 27244 17890 27300 17892
rect 27244 17838 27246 17890
rect 27246 17838 27298 17890
rect 27298 17838 27300 17890
rect 27244 17836 27300 17838
rect 27356 17666 27412 17668
rect 27356 17614 27358 17666
rect 27358 17614 27410 17666
rect 27410 17614 27412 17666
rect 27356 17612 27412 17614
rect 28364 18620 28420 18676
rect 28028 18284 28084 18340
rect 28364 18450 28420 18452
rect 28364 18398 28366 18450
rect 28366 18398 28418 18450
rect 28418 18398 28420 18450
rect 28364 18396 28420 18398
rect 28364 18060 28420 18116
rect 29036 23154 29092 23156
rect 29036 23102 29038 23154
rect 29038 23102 29090 23154
rect 29090 23102 29092 23154
rect 29036 23100 29092 23102
rect 28924 21586 28980 21588
rect 28924 21534 28926 21586
rect 28926 21534 28978 21586
rect 28978 21534 28980 21586
rect 28924 21532 28980 21534
rect 30156 34130 30212 34132
rect 30156 34078 30158 34130
rect 30158 34078 30210 34130
rect 30210 34078 30212 34130
rect 30156 34076 30212 34078
rect 29932 33516 29988 33572
rect 30268 33122 30324 33124
rect 30268 33070 30270 33122
rect 30270 33070 30322 33122
rect 30322 33070 30324 33122
rect 30268 33068 30324 33070
rect 29932 32396 29988 32452
rect 30716 37996 30772 38052
rect 30828 37660 30884 37716
rect 30828 37212 30884 37268
rect 30716 36204 30772 36260
rect 30492 35980 30548 36036
rect 31052 37938 31108 37940
rect 31052 37886 31054 37938
rect 31054 37886 31106 37938
rect 31106 37886 31108 37938
rect 31052 37884 31108 37886
rect 31052 37154 31108 37156
rect 31052 37102 31054 37154
rect 31054 37102 31106 37154
rect 31106 37102 31108 37154
rect 31052 37100 31108 37102
rect 31164 37324 31220 37380
rect 30492 35532 30548 35588
rect 30604 35308 30660 35364
rect 30940 34524 30996 34580
rect 30604 33516 30660 33572
rect 30828 34130 30884 34132
rect 30828 34078 30830 34130
rect 30830 34078 30882 34130
rect 30882 34078 30884 34130
rect 30828 34076 30884 34078
rect 30716 33404 30772 33460
rect 30828 33122 30884 33124
rect 30828 33070 30830 33122
rect 30830 33070 30882 33122
rect 30882 33070 30884 33122
rect 30828 33068 30884 33070
rect 30492 32450 30548 32452
rect 30492 32398 30494 32450
rect 30494 32398 30546 32450
rect 30546 32398 30548 32450
rect 30492 32396 30548 32398
rect 30156 30380 30212 30436
rect 29932 30156 29988 30212
rect 30268 29148 30324 29204
rect 30268 28530 30324 28532
rect 30268 28478 30270 28530
rect 30270 28478 30322 28530
rect 30322 28478 30324 28530
rect 30268 28476 30324 28478
rect 30156 27074 30212 27076
rect 30156 27022 30158 27074
rect 30158 27022 30210 27074
rect 30210 27022 30212 27074
rect 30156 27020 30212 27022
rect 30268 26962 30324 26964
rect 30268 26910 30270 26962
rect 30270 26910 30322 26962
rect 30322 26910 30324 26962
rect 30268 26908 30324 26910
rect 30492 29596 30548 29652
rect 30716 30156 30772 30212
rect 30940 30210 30996 30212
rect 30940 30158 30942 30210
rect 30942 30158 30994 30210
rect 30994 30158 30996 30210
rect 30940 30156 30996 30158
rect 30828 30098 30884 30100
rect 30828 30046 30830 30098
rect 30830 30046 30882 30098
rect 30882 30046 30884 30098
rect 30828 30044 30884 30046
rect 30716 29986 30772 29988
rect 30716 29934 30718 29986
rect 30718 29934 30770 29986
rect 30770 29934 30772 29986
rect 30716 29932 30772 29934
rect 31276 36258 31332 36260
rect 31276 36206 31278 36258
rect 31278 36206 31330 36258
rect 31330 36206 31332 36258
rect 31276 36204 31332 36206
rect 31164 34354 31220 34356
rect 31164 34302 31166 34354
rect 31166 34302 31218 34354
rect 31218 34302 31220 34354
rect 31164 34300 31220 34302
rect 31500 37826 31556 37828
rect 31500 37774 31502 37826
rect 31502 37774 31554 37826
rect 31554 37774 31556 37826
rect 31500 37772 31556 37774
rect 31500 35532 31556 35588
rect 31948 39228 32004 39284
rect 31836 37938 31892 37940
rect 31836 37886 31838 37938
rect 31838 37886 31890 37938
rect 31890 37886 31892 37938
rect 31836 37884 31892 37886
rect 31724 37660 31780 37716
rect 31836 37266 31892 37268
rect 31836 37214 31838 37266
rect 31838 37214 31890 37266
rect 31890 37214 31892 37266
rect 31836 37212 31892 37214
rect 32172 44210 32228 44212
rect 32172 44158 32174 44210
rect 32174 44158 32226 44210
rect 32226 44158 32228 44210
rect 32172 44156 32228 44158
rect 32508 50316 32564 50372
rect 32396 49026 32452 49028
rect 32396 48974 32398 49026
rect 32398 48974 32450 49026
rect 32450 48974 32452 49026
rect 32396 48972 32452 48974
rect 32508 48018 32564 48020
rect 32508 47966 32510 48018
rect 32510 47966 32562 48018
rect 32562 47966 32564 48018
rect 32508 47964 32564 47966
rect 32732 50764 32788 50820
rect 33516 50370 33572 50372
rect 33516 50318 33518 50370
rect 33518 50318 33570 50370
rect 33570 50318 33572 50370
rect 33516 50316 33572 50318
rect 33068 49644 33124 49700
rect 33740 49868 33796 49924
rect 32732 49250 32788 49252
rect 32732 49198 32734 49250
rect 32734 49198 32786 49250
rect 32786 49198 32788 49250
rect 32732 49196 32788 49198
rect 33628 48972 33684 49028
rect 33740 48860 33796 48916
rect 33628 48130 33684 48132
rect 33628 48078 33630 48130
rect 33630 48078 33682 48130
rect 33682 48078 33684 48130
rect 33628 48076 33684 48078
rect 33292 47964 33348 48020
rect 32620 47292 32676 47348
rect 34188 52108 34244 52164
rect 34188 51378 34244 51380
rect 34188 51326 34190 51378
rect 34190 51326 34242 51378
rect 34242 51326 34244 51378
rect 34188 51324 34244 51326
rect 34076 49532 34132 49588
rect 34188 49196 34244 49252
rect 38220 54514 38276 54516
rect 38220 54462 38222 54514
rect 38222 54462 38274 54514
rect 38274 54462 38276 54514
rect 38220 54460 38276 54462
rect 39116 54460 39172 54516
rect 38444 54402 38500 54404
rect 38444 54350 38446 54402
rect 38446 54350 38498 54402
rect 38498 54350 38500 54402
rect 38444 54348 38500 54350
rect 39004 54348 39060 54404
rect 35196 54122 35252 54124
rect 35196 54070 35198 54122
rect 35198 54070 35250 54122
rect 35250 54070 35252 54122
rect 35196 54068 35252 54070
rect 35300 54122 35356 54124
rect 35300 54070 35302 54122
rect 35302 54070 35354 54122
rect 35354 54070 35356 54122
rect 35300 54068 35356 54070
rect 35404 54122 35460 54124
rect 35404 54070 35406 54122
rect 35406 54070 35458 54122
rect 35458 54070 35460 54122
rect 35404 54068 35460 54070
rect 35980 53564 36036 53620
rect 35084 53170 35140 53172
rect 35084 53118 35086 53170
rect 35086 53118 35138 53170
rect 35138 53118 35140 53170
rect 35084 53116 35140 53118
rect 34748 52834 34804 52836
rect 34748 52782 34750 52834
rect 34750 52782 34802 52834
rect 34802 52782 34804 52834
rect 34748 52780 34804 52782
rect 35980 53170 36036 53172
rect 35980 53118 35982 53170
rect 35982 53118 36034 53170
rect 36034 53118 36036 53170
rect 35980 53116 36036 53118
rect 34860 52386 34916 52388
rect 34860 52334 34862 52386
rect 34862 52334 34914 52386
rect 34914 52334 34916 52386
rect 34860 52332 34916 52334
rect 34972 52780 35028 52836
rect 35644 52834 35700 52836
rect 35644 52782 35646 52834
rect 35646 52782 35698 52834
rect 35698 52782 35700 52834
rect 35644 52780 35700 52782
rect 35196 52554 35252 52556
rect 35196 52502 35198 52554
rect 35198 52502 35250 52554
rect 35250 52502 35252 52554
rect 35196 52500 35252 52502
rect 35300 52554 35356 52556
rect 35300 52502 35302 52554
rect 35302 52502 35354 52554
rect 35354 52502 35356 52554
rect 35300 52500 35356 52502
rect 35404 52554 35460 52556
rect 35404 52502 35406 52554
rect 35406 52502 35458 52554
rect 35458 52502 35460 52554
rect 35404 52500 35460 52502
rect 34972 52220 35028 52276
rect 36316 52220 36372 52276
rect 34524 52050 34580 52052
rect 34524 51998 34526 52050
rect 34526 51998 34578 52050
rect 34578 51998 34580 52050
rect 34524 51996 34580 51998
rect 35868 52050 35924 52052
rect 35868 51998 35870 52050
rect 35870 51998 35922 52050
rect 35922 51998 35924 52050
rect 35868 51996 35924 51998
rect 35308 51378 35364 51380
rect 35308 51326 35310 51378
rect 35310 51326 35362 51378
rect 35362 51326 35364 51378
rect 35308 51324 35364 51326
rect 36092 51884 36148 51940
rect 34636 51266 34692 51268
rect 34636 51214 34638 51266
rect 34638 51214 34690 51266
rect 34690 51214 34692 51266
rect 34636 51212 34692 51214
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 36092 50594 36148 50596
rect 36092 50542 36094 50594
rect 36094 50542 36146 50594
rect 36146 50542 36148 50594
rect 36092 50540 36148 50542
rect 34748 50482 34804 50484
rect 34748 50430 34750 50482
rect 34750 50430 34802 50482
rect 34802 50430 34804 50482
rect 34748 50428 34804 50430
rect 35196 50482 35252 50484
rect 35196 50430 35198 50482
rect 35198 50430 35250 50482
rect 35250 50430 35252 50482
rect 35196 50428 35252 50430
rect 37884 52668 37940 52724
rect 36652 52274 36708 52276
rect 36652 52222 36654 52274
rect 36654 52222 36706 52274
rect 36706 52222 36708 52274
rect 36652 52220 36708 52222
rect 36540 51996 36596 52052
rect 37436 51884 37492 51940
rect 36428 51324 36484 51380
rect 34524 48972 34580 49028
rect 33964 48802 34020 48804
rect 33964 48750 33966 48802
rect 33966 48750 34018 48802
rect 34018 48750 34020 48802
rect 33964 48748 34020 48750
rect 33852 47852 33908 47908
rect 34076 48188 34132 48244
rect 33964 47964 34020 48020
rect 33740 47740 33796 47796
rect 33628 47346 33684 47348
rect 33628 47294 33630 47346
rect 33630 47294 33682 47346
rect 33682 47294 33684 47346
rect 33628 47292 33684 47294
rect 34300 47346 34356 47348
rect 34300 47294 34302 47346
rect 34302 47294 34354 47346
rect 34354 47294 34356 47346
rect 34300 47292 34356 47294
rect 36316 50316 36372 50372
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35084 49026 35140 49028
rect 35084 48974 35086 49026
rect 35086 48974 35138 49026
rect 35138 48974 35140 49026
rect 35084 48972 35140 48974
rect 35644 49586 35700 49588
rect 35644 49534 35646 49586
rect 35646 49534 35698 49586
rect 35698 49534 35700 49586
rect 35644 49532 35700 49534
rect 35868 48860 35924 48916
rect 35196 48802 35252 48804
rect 35196 48750 35198 48802
rect 35198 48750 35250 48802
rect 35250 48750 35252 48802
rect 35196 48748 35252 48750
rect 34748 48636 34804 48692
rect 35084 48524 35140 48580
rect 34524 47740 34580 47796
rect 34748 47852 34804 47908
rect 34860 47516 34916 47572
rect 33964 46844 34020 46900
rect 33740 46786 33796 46788
rect 33740 46734 33742 46786
rect 33742 46734 33794 46786
rect 33794 46734 33796 46786
rect 33740 46732 33796 46734
rect 32396 46674 32452 46676
rect 32396 46622 32398 46674
rect 32398 46622 32450 46674
rect 32450 46622 32452 46674
rect 32396 46620 32452 46622
rect 32508 46562 32564 46564
rect 32508 46510 32510 46562
rect 32510 46510 32562 46562
rect 32562 46510 32564 46562
rect 32508 46508 32564 46510
rect 33628 46562 33684 46564
rect 33628 46510 33630 46562
rect 33630 46510 33682 46562
rect 33682 46510 33684 46562
rect 33628 46508 33684 46510
rect 32620 43932 32676 43988
rect 32732 44156 32788 44212
rect 33740 45388 33796 45444
rect 33628 44268 33684 44324
rect 32284 43484 32340 43540
rect 32844 44098 32900 44100
rect 32844 44046 32846 44098
rect 32846 44046 32898 44098
rect 32898 44046 32900 44098
rect 32844 44044 32900 44046
rect 33180 44098 33236 44100
rect 33180 44046 33182 44098
rect 33182 44046 33234 44098
rect 33234 44046 33236 44098
rect 33180 44044 33236 44046
rect 32956 43932 33012 43988
rect 32732 43260 32788 43316
rect 32508 42754 32564 42756
rect 32508 42702 32510 42754
rect 32510 42702 32562 42754
rect 32562 42702 32564 42754
rect 32508 42700 32564 42702
rect 32732 42754 32788 42756
rect 32732 42702 32734 42754
rect 32734 42702 32786 42754
rect 32786 42702 32788 42754
rect 32732 42700 32788 42702
rect 32620 42642 32676 42644
rect 32620 42590 32622 42642
rect 32622 42590 32674 42642
rect 32674 42590 32676 42642
rect 32620 42588 32676 42590
rect 32956 42530 33012 42532
rect 32956 42478 32958 42530
rect 32958 42478 33010 42530
rect 33010 42478 33012 42530
rect 32956 42476 33012 42478
rect 32284 39004 32340 39060
rect 32956 39564 33012 39620
rect 32844 39506 32900 39508
rect 32844 39454 32846 39506
rect 32846 39454 32898 39506
rect 32898 39454 32900 39506
rect 32844 39452 32900 39454
rect 32060 37100 32116 37156
rect 32396 37324 32452 37380
rect 32620 37378 32676 37380
rect 32620 37326 32622 37378
rect 32622 37326 32674 37378
rect 32674 37326 32676 37378
rect 32620 37324 32676 37326
rect 32732 37212 32788 37268
rect 31948 35980 32004 36036
rect 31836 35922 31892 35924
rect 31836 35870 31838 35922
rect 31838 35870 31890 35922
rect 31890 35870 31892 35922
rect 31836 35868 31892 35870
rect 31612 35420 31668 35476
rect 31836 34690 31892 34692
rect 31836 34638 31838 34690
rect 31838 34638 31890 34690
rect 31890 34638 31892 34690
rect 31836 34636 31892 34638
rect 31724 34524 31780 34580
rect 31388 31836 31444 31892
rect 31164 31276 31220 31332
rect 30716 29708 30772 29764
rect 31388 31052 31444 31108
rect 31500 31164 31556 31220
rect 30604 28642 30660 28644
rect 30604 28590 30606 28642
rect 30606 28590 30658 28642
rect 30658 28590 30660 28642
rect 30604 28588 30660 28590
rect 30044 26012 30100 26068
rect 29932 24892 29988 24948
rect 29820 24108 29876 24164
rect 29484 23714 29540 23716
rect 29484 23662 29486 23714
rect 29486 23662 29538 23714
rect 29538 23662 29540 23714
rect 29484 23660 29540 23662
rect 29708 23772 29764 23828
rect 29484 23378 29540 23380
rect 29484 23326 29486 23378
rect 29486 23326 29538 23378
rect 29538 23326 29540 23378
rect 29484 23324 29540 23326
rect 29372 22540 29428 22596
rect 29036 20524 29092 20580
rect 29036 20130 29092 20132
rect 29036 20078 29038 20130
rect 29038 20078 29090 20130
rect 29090 20078 29092 20130
rect 29036 20076 29092 20078
rect 28924 18508 28980 18564
rect 28476 17836 28532 17892
rect 28700 18396 28756 18452
rect 28252 17724 28308 17780
rect 28588 17724 28644 17780
rect 27916 17442 27972 17444
rect 27916 17390 27918 17442
rect 27918 17390 27970 17442
rect 27970 17390 27972 17442
rect 27916 17388 27972 17390
rect 28252 17276 28308 17332
rect 28028 16940 28084 16996
rect 27244 15314 27300 15316
rect 27244 15262 27246 15314
rect 27246 15262 27298 15314
rect 27298 15262 27300 15314
rect 27244 15260 27300 15262
rect 27468 15148 27524 15204
rect 27356 13580 27412 13636
rect 27916 16380 27972 16436
rect 28252 15596 28308 15652
rect 27804 15314 27860 15316
rect 27804 15262 27806 15314
rect 27806 15262 27858 15314
rect 27858 15262 27860 15314
rect 27804 15260 27860 15262
rect 28588 15260 28644 15316
rect 27468 12290 27524 12292
rect 27468 12238 27470 12290
rect 27470 12238 27522 12290
rect 27522 12238 27524 12290
rect 27468 12236 27524 12238
rect 27916 14306 27972 14308
rect 27916 14254 27918 14306
rect 27918 14254 27970 14306
rect 27970 14254 27972 14306
rect 27916 14252 27972 14254
rect 28476 14306 28532 14308
rect 28476 14254 28478 14306
rect 28478 14254 28530 14306
rect 28530 14254 28532 14306
rect 28476 14252 28532 14254
rect 27804 13580 27860 13636
rect 28252 13522 28308 13524
rect 28252 13470 28254 13522
rect 28254 13470 28306 13522
rect 28306 13470 28308 13522
rect 28252 13468 28308 13470
rect 27244 11228 27300 11284
rect 27244 10780 27300 10836
rect 27132 9996 27188 10052
rect 27020 9826 27076 9828
rect 27020 9774 27022 9826
rect 27022 9774 27074 9826
rect 27074 9774 27076 9826
rect 27020 9772 27076 9774
rect 26908 9042 26964 9044
rect 26908 8990 26910 9042
rect 26910 8990 26962 9042
rect 26962 8990 26964 9042
rect 26908 8988 26964 8990
rect 26684 7980 26740 8036
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 26908 7868 26964 7924
rect 26460 7420 26516 7476
rect 26908 7084 26964 7140
rect 26572 6466 26628 6468
rect 26572 6414 26574 6466
rect 26574 6414 26626 6466
rect 26626 6414 26628 6466
rect 26572 6412 26628 6414
rect 26348 2604 26404 2660
rect 26012 2492 26068 2548
rect 27356 9884 27412 9940
rect 27468 8988 27524 9044
rect 27244 8034 27300 8036
rect 27244 7982 27246 8034
rect 27246 7982 27298 8034
rect 27298 7982 27300 8034
rect 27244 7980 27300 7982
rect 27356 5068 27412 5124
rect 27020 3276 27076 3332
rect 26908 2268 26964 2324
rect 28028 11506 28084 11508
rect 28028 11454 28030 11506
rect 28030 11454 28082 11506
rect 28082 11454 28084 11506
rect 28028 11452 28084 11454
rect 28476 12850 28532 12852
rect 28476 12798 28478 12850
rect 28478 12798 28530 12850
rect 28530 12798 28532 12850
rect 28476 12796 28532 12798
rect 28812 16828 28868 16884
rect 28924 17388 28980 17444
rect 28924 16492 28980 16548
rect 28812 16380 28868 16436
rect 28812 15314 28868 15316
rect 28812 15262 28814 15314
rect 28814 15262 28866 15314
rect 28866 15262 28868 15314
rect 28812 15260 28868 15262
rect 28476 12236 28532 12292
rect 28252 11116 28308 11172
rect 28140 10610 28196 10612
rect 28140 10558 28142 10610
rect 28142 10558 28194 10610
rect 28194 10558 28196 10610
rect 28140 10556 28196 10558
rect 27692 7868 27748 7924
rect 28028 6748 28084 6804
rect 28924 12178 28980 12180
rect 28924 12126 28926 12178
rect 28926 12126 28978 12178
rect 28978 12126 28980 12178
rect 28924 12124 28980 12126
rect 29596 22316 29652 22372
rect 29484 21362 29540 21364
rect 29484 21310 29486 21362
rect 29486 21310 29538 21362
rect 29538 21310 29540 21362
rect 29484 21308 29540 21310
rect 29932 23826 29988 23828
rect 29932 23774 29934 23826
rect 29934 23774 29986 23826
rect 29986 23774 29988 23826
rect 29932 23772 29988 23774
rect 29820 23660 29876 23716
rect 29932 23154 29988 23156
rect 29932 23102 29934 23154
rect 29934 23102 29986 23154
rect 29986 23102 29988 23154
rect 29932 23100 29988 23102
rect 29932 22594 29988 22596
rect 29932 22542 29934 22594
rect 29934 22542 29986 22594
rect 29986 22542 29988 22594
rect 29932 22540 29988 22542
rect 30380 24332 30436 24388
rect 30156 22258 30212 22260
rect 30156 22206 30158 22258
rect 30158 22206 30210 22258
rect 30210 22206 30212 22258
rect 30156 22204 30212 22206
rect 30044 21698 30100 21700
rect 30044 21646 30046 21698
rect 30046 21646 30098 21698
rect 30098 21646 30100 21698
rect 30044 21644 30100 21646
rect 29932 20636 29988 20692
rect 30044 20578 30100 20580
rect 30044 20526 30046 20578
rect 30046 20526 30098 20578
rect 30098 20526 30100 20578
rect 30044 20524 30100 20526
rect 29820 20076 29876 20132
rect 29260 17612 29316 17668
rect 29708 20018 29764 20020
rect 29708 19966 29710 20018
rect 29710 19966 29762 20018
rect 29762 19966 29764 20018
rect 29708 19964 29764 19966
rect 30156 19852 30212 19908
rect 29932 19122 29988 19124
rect 29932 19070 29934 19122
rect 29934 19070 29986 19122
rect 29986 19070 29988 19122
rect 29932 19068 29988 19070
rect 30380 20524 30436 20580
rect 30604 23548 30660 23604
rect 31276 30828 31332 30884
rect 31500 30434 31556 30436
rect 31500 30382 31502 30434
rect 31502 30382 31554 30434
rect 31554 30382 31556 30434
rect 31500 30380 31556 30382
rect 31052 28588 31108 28644
rect 31052 28082 31108 28084
rect 31052 28030 31054 28082
rect 31054 28030 31106 28082
rect 31106 28030 31108 28082
rect 31052 28028 31108 28030
rect 31276 28866 31332 28868
rect 31276 28814 31278 28866
rect 31278 28814 31330 28866
rect 31330 28814 31332 28866
rect 31276 28812 31332 28814
rect 31276 28530 31332 28532
rect 31276 28478 31278 28530
rect 31278 28478 31330 28530
rect 31330 28478 31332 28530
rect 31276 28476 31332 28478
rect 31500 28364 31556 28420
rect 30940 27244 30996 27300
rect 30828 26908 30884 26964
rect 31276 27020 31332 27076
rect 31500 27356 31556 27412
rect 31948 31836 32004 31892
rect 31948 31218 32004 31220
rect 31948 31166 31950 31218
rect 31950 31166 32002 31218
rect 32002 31166 32004 31218
rect 31948 31164 32004 31166
rect 31836 29932 31892 29988
rect 31724 29148 31780 29204
rect 32172 36428 32228 36484
rect 32732 36482 32788 36484
rect 32732 36430 32734 36482
rect 32734 36430 32786 36482
rect 32786 36430 32788 36482
rect 32732 36428 32788 36430
rect 32396 35980 32452 36036
rect 32956 37490 33012 37492
rect 32956 37438 32958 37490
rect 32958 37438 33010 37490
rect 33010 37438 33012 37490
rect 32956 37436 33012 37438
rect 33404 43260 33460 43316
rect 33180 36594 33236 36596
rect 33180 36542 33182 36594
rect 33182 36542 33234 36594
rect 33234 36542 33236 36594
rect 33180 36540 33236 36542
rect 33068 35868 33124 35924
rect 32732 35420 32788 35476
rect 33180 36316 33236 36372
rect 32396 34690 32452 34692
rect 32396 34638 32398 34690
rect 32398 34638 32450 34690
rect 32450 34638 32452 34690
rect 32396 34636 32452 34638
rect 32284 34300 32340 34356
rect 32508 33346 32564 33348
rect 32508 33294 32510 33346
rect 32510 33294 32562 33346
rect 32562 33294 32564 33346
rect 32508 33292 32564 33294
rect 32396 33122 32452 33124
rect 32396 33070 32398 33122
rect 32398 33070 32450 33122
rect 32450 33070 32452 33122
rect 32396 33068 32452 33070
rect 32844 32450 32900 32452
rect 32844 32398 32846 32450
rect 32846 32398 32898 32450
rect 32898 32398 32900 32450
rect 32844 32396 32900 32398
rect 32956 31948 33012 32004
rect 32732 31164 32788 31220
rect 32284 30210 32340 30212
rect 32284 30158 32286 30210
rect 32286 30158 32338 30210
rect 32338 30158 32340 30210
rect 32284 30156 32340 30158
rect 32508 28924 32564 28980
rect 32172 28700 32228 28756
rect 32284 28812 32340 28868
rect 32172 28530 32228 28532
rect 32172 28478 32174 28530
rect 32174 28478 32226 28530
rect 32226 28478 32228 28530
rect 32172 28476 32228 28478
rect 31724 28082 31780 28084
rect 31724 28030 31726 28082
rect 31726 28030 31778 28082
rect 31778 28030 31780 28082
rect 31724 28028 31780 28030
rect 32396 28028 32452 28084
rect 31724 27356 31780 27412
rect 31276 25900 31332 25956
rect 31052 25564 31108 25620
rect 31500 26236 31556 26292
rect 31724 26178 31780 26180
rect 31724 26126 31726 26178
rect 31726 26126 31778 26178
rect 31778 26126 31780 26178
rect 31724 26124 31780 26126
rect 31612 25900 31668 25956
rect 32172 26908 32228 26964
rect 32396 26796 32452 26852
rect 32172 26402 32228 26404
rect 32172 26350 32174 26402
rect 32174 26350 32226 26402
rect 32226 26350 32228 26402
rect 32172 26348 32228 26350
rect 32060 26290 32116 26292
rect 32060 26238 32062 26290
rect 32062 26238 32114 26290
rect 32114 26238 32116 26290
rect 32060 26236 32116 26238
rect 31948 26124 32004 26180
rect 32284 25900 32340 25956
rect 32060 25618 32116 25620
rect 32060 25566 32062 25618
rect 32062 25566 32114 25618
rect 32114 25566 32116 25618
rect 32060 25564 32116 25566
rect 30828 24220 30884 24276
rect 31164 24556 31220 24612
rect 32284 25394 32340 25396
rect 32284 25342 32286 25394
rect 32286 25342 32338 25394
rect 32338 25342 32340 25394
rect 32284 25340 32340 25342
rect 31276 25116 31332 25172
rect 31164 24162 31220 24164
rect 31164 24110 31166 24162
rect 31166 24110 31218 24162
rect 31218 24110 31220 24162
rect 31164 24108 31220 24110
rect 30716 22428 30772 22484
rect 30604 22258 30660 22260
rect 30604 22206 30606 22258
rect 30606 22206 30658 22258
rect 30658 22206 30660 22258
rect 30604 22204 30660 22206
rect 30828 21810 30884 21812
rect 30828 21758 30830 21810
rect 30830 21758 30882 21810
rect 30882 21758 30884 21810
rect 30828 21756 30884 21758
rect 31724 25228 31780 25284
rect 31612 24610 31668 24612
rect 31612 24558 31614 24610
rect 31614 24558 31666 24610
rect 31666 24558 31668 24610
rect 31612 24556 31668 24558
rect 32172 24556 32228 24612
rect 32060 24444 32116 24500
rect 31500 23938 31556 23940
rect 31500 23886 31502 23938
rect 31502 23886 31554 23938
rect 31554 23886 31556 23938
rect 31500 23884 31556 23886
rect 31388 22482 31444 22484
rect 31388 22430 31390 22482
rect 31390 22430 31442 22482
rect 31442 22430 31444 22482
rect 31388 22428 31444 22430
rect 31276 21756 31332 21812
rect 31276 21586 31332 21588
rect 31276 21534 31278 21586
rect 31278 21534 31330 21586
rect 31330 21534 31332 21586
rect 31276 21532 31332 21534
rect 30716 21308 30772 21364
rect 30828 20802 30884 20804
rect 30828 20750 30830 20802
rect 30830 20750 30882 20802
rect 30882 20750 30884 20802
rect 30828 20748 30884 20750
rect 31500 20636 31556 20692
rect 30268 19068 30324 19124
rect 30268 18844 30324 18900
rect 29708 18732 29764 18788
rect 30156 18732 30212 18788
rect 29596 18396 29652 18452
rect 29484 17724 29540 17780
rect 29820 17666 29876 17668
rect 29820 17614 29822 17666
rect 29822 17614 29874 17666
rect 29874 17614 29876 17666
rect 29820 17612 29876 17614
rect 29484 17442 29540 17444
rect 29484 17390 29486 17442
rect 29486 17390 29538 17442
rect 29538 17390 29540 17442
rect 29484 17388 29540 17390
rect 29148 16828 29204 16884
rect 29932 16098 29988 16100
rect 29932 16046 29934 16098
rect 29934 16046 29986 16098
rect 29986 16046 29988 16098
rect 29932 16044 29988 16046
rect 29484 15708 29540 15764
rect 29596 15596 29652 15652
rect 29260 15538 29316 15540
rect 29260 15486 29262 15538
rect 29262 15486 29314 15538
rect 29314 15486 29316 15538
rect 29260 15484 29316 15486
rect 29036 11340 29092 11396
rect 28588 10780 28644 10836
rect 28364 9884 28420 9940
rect 28476 10444 28532 10500
rect 28364 9266 28420 9268
rect 28364 9214 28366 9266
rect 28366 9214 28418 9266
rect 28418 9214 28420 9266
rect 28364 9212 28420 9214
rect 28700 10556 28756 10612
rect 28700 9436 28756 9492
rect 28476 5964 28532 6020
rect 28812 5234 28868 5236
rect 28812 5182 28814 5234
rect 28814 5182 28866 5234
rect 28866 5182 28868 5234
rect 28812 5180 28868 5182
rect 28364 5010 28420 5012
rect 28364 4958 28366 5010
rect 28366 4958 28418 5010
rect 28418 4958 28420 5010
rect 28364 4956 28420 4958
rect 28140 4508 28196 4564
rect 28028 3948 28084 4004
rect 27580 1372 27636 1428
rect 28252 3388 28308 3444
rect 29372 15036 29428 15092
rect 29260 10498 29316 10500
rect 29260 10446 29262 10498
rect 29262 10446 29314 10498
rect 29314 10446 29316 10498
rect 29260 10444 29316 10446
rect 29932 15596 29988 15652
rect 30044 15036 30100 15092
rect 30156 15148 30212 15204
rect 29708 14588 29764 14644
rect 29484 14476 29540 14532
rect 30044 14530 30100 14532
rect 30044 14478 30046 14530
rect 30046 14478 30098 14530
rect 30098 14478 30100 14530
rect 30044 14476 30100 14478
rect 30604 18732 30660 18788
rect 31276 19906 31332 19908
rect 31276 19854 31278 19906
rect 31278 19854 31330 19906
rect 31330 19854 31332 19906
rect 31276 19852 31332 19854
rect 31276 18844 31332 18900
rect 31276 18674 31332 18676
rect 31276 18622 31278 18674
rect 31278 18622 31330 18674
rect 31330 18622 31332 18674
rect 31276 18620 31332 18622
rect 31500 18674 31556 18676
rect 31500 18622 31502 18674
rect 31502 18622 31554 18674
rect 31554 18622 31556 18674
rect 31500 18620 31556 18622
rect 31164 18508 31220 18564
rect 30492 17442 30548 17444
rect 30492 17390 30494 17442
rect 30494 17390 30546 17442
rect 30546 17390 30548 17442
rect 30492 17388 30548 17390
rect 30380 17164 30436 17220
rect 30380 16098 30436 16100
rect 30380 16046 30382 16098
rect 30382 16046 30434 16098
rect 30434 16046 30436 16098
rect 30380 16044 30436 16046
rect 31052 17276 31108 17332
rect 30828 16268 30884 16324
rect 30604 15484 30660 15540
rect 30380 15314 30436 15316
rect 30380 15262 30382 15314
rect 30382 15262 30434 15314
rect 30434 15262 30436 15314
rect 30380 15260 30436 15262
rect 30828 15820 30884 15876
rect 30828 15260 30884 15316
rect 30716 15148 30772 15204
rect 30268 14642 30324 14644
rect 30268 14590 30270 14642
rect 30270 14590 30322 14642
rect 30322 14590 30324 14642
rect 30268 14588 30324 14590
rect 30604 14306 30660 14308
rect 30604 14254 30606 14306
rect 30606 14254 30658 14306
rect 30658 14254 30660 14306
rect 30604 14252 30660 14254
rect 30828 14476 30884 14532
rect 30492 14028 30548 14084
rect 30940 13970 30996 13972
rect 30940 13918 30942 13970
rect 30942 13918 30994 13970
rect 30994 13918 30996 13970
rect 30940 13916 30996 13918
rect 30380 13746 30436 13748
rect 30380 13694 30382 13746
rect 30382 13694 30434 13746
rect 30434 13694 30436 13746
rect 30380 13692 30436 13694
rect 29932 13634 29988 13636
rect 29932 13582 29934 13634
rect 29934 13582 29986 13634
rect 29986 13582 29988 13634
rect 29932 13580 29988 13582
rect 29708 12572 29764 12628
rect 29820 13020 29876 13076
rect 29820 12796 29876 12852
rect 29932 12572 29988 12628
rect 30492 13020 30548 13076
rect 29596 11788 29652 11844
rect 30268 11788 30324 11844
rect 29596 11282 29652 11284
rect 29596 11230 29598 11282
rect 29598 11230 29650 11282
rect 29650 11230 29652 11282
rect 29596 11228 29652 11230
rect 29820 10834 29876 10836
rect 29820 10782 29822 10834
rect 29822 10782 29874 10834
rect 29874 10782 29876 10834
rect 29820 10780 29876 10782
rect 30156 10722 30212 10724
rect 30156 10670 30158 10722
rect 30158 10670 30210 10722
rect 30210 10670 30212 10722
rect 30156 10668 30212 10670
rect 29932 10444 29988 10500
rect 29484 9938 29540 9940
rect 29484 9886 29486 9938
rect 29486 9886 29538 9938
rect 29538 9886 29540 9938
rect 29484 9884 29540 9886
rect 29372 8204 29428 8260
rect 30828 13074 30884 13076
rect 30828 13022 30830 13074
rect 30830 13022 30882 13074
rect 30882 13022 30884 13074
rect 30828 13020 30884 13022
rect 30716 12124 30772 12180
rect 30828 11004 30884 11060
rect 30716 10332 30772 10388
rect 30380 6076 30436 6132
rect 31276 17052 31332 17108
rect 31164 14812 31220 14868
rect 31276 15202 31332 15204
rect 31276 15150 31278 15202
rect 31278 15150 31330 15202
rect 31330 15150 31332 15202
rect 31276 15148 31332 15150
rect 31836 23996 31892 24052
rect 32060 22876 32116 22932
rect 31836 22370 31892 22372
rect 31836 22318 31838 22370
rect 31838 22318 31890 22370
rect 31890 22318 31892 22370
rect 31836 22316 31892 22318
rect 32060 21980 32116 22036
rect 32284 23884 32340 23940
rect 32620 28082 32676 28084
rect 32620 28030 32622 28082
rect 32622 28030 32674 28082
rect 32674 28030 32676 28082
rect 32620 28028 32676 28030
rect 32508 26348 32564 26404
rect 32844 30380 32900 30436
rect 32732 26908 32788 26964
rect 33292 33346 33348 33348
rect 33292 33294 33294 33346
rect 33294 33294 33346 33346
rect 33346 33294 33348 33346
rect 33292 33292 33348 33294
rect 33180 31164 33236 31220
rect 33180 29986 33236 29988
rect 33180 29934 33182 29986
rect 33182 29934 33234 29986
rect 33234 29934 33236 29986
rect 33180 29932 33236 29934
rect 33180 29036 33236 29092
rect 33068 28812 33124 28868
rect 32620 26124 32676 26180
rect 32508 25004 32564 25060
rect 32732 23772 32788 23828
rect 32396 23266 32452 23268
rect 32396 23214 32398 23266
rect 32398 23214 32450 23266
rect 32450 23214 32452 23266
rect 32396 23212 32452 23214
rect 32284 22988 32340 23044
rect 32620 23378 32676 23380
rect 32620 23326 32622 23378
rect 32622 23326 32674 23378
rect 32674 23326 32676 23378
rect 32620 23324 32676 23326
rect 32284 20914 32340 20916
rect 32284 20862 32286 20914
rect 32286 20862 32338 20914
rect 32338 20862 32340 20914
rect 32284 20860 32340 20862
rect 31836 20188 31892 20244
rect 31948 20524 32004 20580
rect 31724 19628 31780 19684
rect 31836 18732 31892 18788
rect 32172 18562 32228 18564
rect 32172 18510 32174 18562
rect 32174 18510 32226 18562
rect 32226 18510 32228 18562
rect 32172 18508 32228 18510
rect 32060 17554 32116 17556
rect 32060 17502 32062 17554
rect 32062 17502 32114 17554
rect 32114 17502 32116 17554
rect 32060 17500 32116 17502
rect 31612 17276 31668 17332
rect 32172 17276 32228 17332
rect 31724 17164 31780 17220
rect 32284 17164 32340 17220
rect 32172 17106 32228 17108
rect 32172 17054 32174 17106
rect 32174 17054 32226 17106
rect 32226 17054 32228 17106
rect 32172 17052 32228 17054
rect 31948 16940 32004 16996
rect 32060 16828 32116 16884
rect 31724 15874 31780 15876
rect 31724 15822 31726 15874
rect 31726 15822 31778 15874
rect 31778 15822 31780 15874
rect 31724 15820 31780 15822
rect 32956 24946 33012 24948
rect 32956 24894 32958 24946
rect 32958 24894 33010 24946
rect 33010 24894 33012 24946
rect 32956 24892 33012 24894
rect 34412 46674 34468 46676
rect 34412 46622 34414 46674
rect 34414 46622 34466 46674
rect 34466 46622 34468 46674
rect 34412 46620 34468 46622
rect 34524 45388 34580 45444
rect 34188 44492 34244 44548
rect 34524 43596 34580 43652
rect 34860 46732 34916 46788
rect 35756 48242 35812 48244
rect 35756 48190 35758 48242
rect 35758 48190 35810 48242
rect 35810 48190 35812 48242
rect 35756 48188 35812 48190
rect 35532 48018 35588 48020
rect 35532 47966 35534 48018
rect 35534 47966 35586 48018
rect 35586 47966 35588 48018
rect 35532 47964 35588 47966
rect 35980 47964 36036 48020
rect 37548 51548 37604 51604
rect 37436 51378 37492 51380
rect 37436 51326 37438 51378
rect 37438 51326 37490 51378
rect 37490 51326 37492 51378
rect 37436 51324 37492 51326
rect 37996 52220 38052 52276
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 36092 47740 36148 47796
rect 35084 47292 35140 47348
rect 33852 42700 33908 42756
rect 33516 42530 33572 42532
rect 33516 42478 33518 42530
rect 33518 42478 33570 42530
rect 33570 42478 33572 42530
rect 33516 42476 33572 42478
rect 34076 42082 34132 42084
rect 34076 42030 34078 42082
rect 34078 42030 34130 42082
rect 34130 42030 34132 42082
rect 34076 42028 34132 42030
rect 33628 41970 33684 41972
rect 33628 41918 33630 41970
rect 33630 41918 33682 41970
rect 33682 41918 33684 41970
rect 33628 41916 33684 41918
rect 34300 41692 34356 41748
rect 33852 41074 33908 41076
rect 33852 41022 33854 41074
rect 33854 41022 33906 41074
rect 33906 41022 33908 41074
rect 33852 41020 33908 41022
rect 33628 40348 33684 40404
rect 33628 39058 33684 39060
rect 33628 39006 33630 39058
rect 33630 39006 33682 39058
rect 33682 39006 33684 39058
rect 33628 39004 33684 39006
rect 33852 40514 33908 40516
rect 33852 40462 33854 40514
rect 33854 40462 33906 40514
rect 33906 40462 33908 40514
rect 33852 40460 33908 40462
rect 34076 40962 34132 40964
rect 34076 40910 34078 40962
rect 34078 40910 34130 40962
rect 34130 40910 34132 40962
rect 34076 40908 34132 40910
rect 33740 38668 33796 38724
rect 34076 40460 34132 40516
rect 33740 38108 33796 38164
rect 33516 37436 33572 37492
rect 33628 37266 33684 37268
rect 33628 37214 33630 37266
rect 33630 37214 33682 37266
rect 33682 37214 33684 37266
rect 33628 37212 33684 37214
rect 34300 40348 34356 40404
rect 34188 38668 34244 38724
rect 33964 38556 34020 38612
rect 34076 38108 34132 38164
rect 34300 37996 34356 38052
rect 33628 36482 33684 36484
rect 33628 36430 33630 36482
rect 33630 36430 33682 36482
rect 33682 36430 33684 36482
rect 33628 36428 33684 36430
rect 34188 35980 34244 36036
rect 33516 33346 33572 33348
rect 33516 33294 33518 33346
rect 33518 33294 33570 33346
rect 33570 33294 33572 33346
rect 33516 33292 33572 33294
rect 33740 34690 33796 34692
rect 33740 34638 33742 34690
rect 33742 34638 33794 34690
rect 33794 34638 33796 34690
rect 33740 34636 33796 34638
rect 33628 33068 33684 33124
rect 33740 33516 33796 33572
rect 33740 32396 33796 32452
rect 33852 33068 33908 33124
rect 33740 31778 33796 31780
rect 33740 31726 33742 31778
rect 33742 31726 33794 31778
rect 33794 31726 33796 31778
rect 33740 31724 33796 31726
rect 33628 31106 33684 31108
rect 33628 31054 33630 31106
rect 33630 31054 33682 31106
rect 33682 31054 33684 31106
rect 33628 31052 33684 31054
rect 33516 30380 33572 30436
rect 34188 32396 34244 32452
rect 34412 37212 34468 37268
rect 34412 34690 34468 34692
rect 34412 34638 34414 34690
rect 34414 34638 34466 34690
rect 34466 34638 34468 34690
rect 34412 34636 34468 34638
rect 34748 42252 34804 42308
rect 34748 40908 34804 40964
rect 36652 47740 36708 47796
rect 36764 50594 36820 50596
rect 36764 50542 36766 50594
rect 36766 50542 36818 50594
rect 36818 50542 36820 50594
rect 36764 50540 36820 50542
rect 38332 52274 38388 52276
rect 38332 52222 38334 52274
rect 38334 52222 38386 52274
rect 38386 52222 38388 52274
rect 38332 52220 38388 52222
rect 38108 52108 38164 52164
rect 36764 48412 36820 48468
rect 36988 48242 37044 48244
rect 36988 48190 36990 48242
rect 36990 48190 37042 48242
rect 37042 48190 37044 48242
rect 36988 48188 37044 48190
rect 37660 49644 37716 49700
rect 37324 48466 37380 48468
rect 37324 48414 37326 48466
rect 37326 48414 37378 48466
rect 37378 48414 37380 48466
rect 37324 48412 37380 48414
rect 37548 48188 37604 48244
rect 37100 47964 37156 48020
rect 35644 47068 35700 47124
rect 36988 46844 37044 46900
rect 36316 46620 36372 46676
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 37212 45836 37268 45892
rect 36652 45778 36708 45780
rect 36652 45726 36654 45778
rect 36654 45726 36706 45778
rect 36706 45726 36708 45778
rect 36652 45724 36708 45726
rect 35196 45388 35252 45444
rect 36540 45612 36596 45668
rect 35532 45164 35588 45220
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35084 44380 35140 44436
rect 36428 45218 36484 45220
rect 36428 45166 36430 45218
rect 36430 45166 36482 45218
rect 36482 45166 36484 45218
rect 36428 45164 36484 45166
rect 35420 44322 35476 44324
rect 35420 44270 35422 44322
rect 35422 44270 35474 44322
rect 35474 44270 35476 44322
rect 35420 44268 35476 44270
rect 36204 44828 36260 44884
rect 35084 44210 35140 44212
rect 35084 44158 35086 44210
rect 35086 44158 35138 44210
rect 35138 44158 35140 44210
rect 35084 44156 35140 44158
rect 36428 44604 36484 44660
rect 36316 44546 36372 44548
rect 36316 44494 36318 44546
rect 36318 44494 36370 44546
rect 36370 44494 36372 44546
rect 36316 44492 36372 44494
rect 36652 45500 36708 45556
rect 36204 44156 36260 44212
rect 35868 43596 35924 43652
rect 35084 43426 35140 43428
rect 35084 43374 35086 43426
rect 35086 43374 35138 43426
rect 35138 43374 35140 43426
rect 35084 43372 35140 43374
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 36092 42866 36148 42868
rect 36092 42814 36094 42866
rect 36094 42814 36146 42866
rect 36146 42814 36148 42866
rect 36092 42812 36148 42814
rect 35420 42530 35476 42532
rect 35420 42478 35422 42530
rect 35422 42478 35474 42530
rect 35474 42478 35476 42530
rect 35420 42476 35476 42478
rect 34972 41858 35028 41860
rect 34972 41806 34974 41858
rect 34974 41806 35026 41858
rect 35026 41806 35028 41858
rect 34972 41804 35028 41806
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35420 41186 35476 41188
rect 35420 41134 35422 41186
rect 35422 41134 35474 41186
rect 35474 41134 35476 41186
rect 35420 41132 35476 41134
rect 35868 42476 35924 42532
rect 36092 42252 36148 42308
rect 35756 42028 35812 42084
rect 35980 42028 36036 42084
rect 35644 41970 35700 41972
rect 35644 41918 35646 41970
rect 35646 41918 35698 41970
rect 35698 41918 35700 41970
rect 35644 41916 35700 41918
rect 35756 41692 35812 41748
rect 35532 41020 35588 41076
rect 35308 40572 35364 40628
rect 36204 40626 36260 40628
rect 36204 40574 36206 40626
rect 36206 40574 36258 40626
rect 36258 40574 36260 40626
rect 36204 40572 36260 40574
rect 36428 40684 36484 40740
rect 35644 40348 35700 40404
rect 35532 40236 35588 40292
rect 35084 40178 35140 40180
rect 35084 40126 35086 40178
rect 35086 40126 35138 40178
rect 35138 40126 35140 40178
rect 35084 40124 35140 40126
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35084 39340 35140 39396
rect 37884 49026 37940 49028
rect 37884 48974 37886 49026
rect 37886 48974 37938 49026
rect 37938 48974 37940 49026
rect 37884 48972 37940 48974
rect 37772 48412 37828 48468
rect 38332 51602 38388 51604
rect 38332 51550 38334 51602
rect 38334 51550 38386 51602
rect 38386 51550 38388 51602
rect 38332 51548 38388 51550
rect 38220 51436 38276 51492
rect 41132 55244 41188 55300
rect 41244 55580 41300 55636
rect 40796 54514 40852 54516
rect 40796 54462 40798 54514
rect 40798 54462 40850 54514
rect 40850 54462 40852 54514
rect 40796 54460 40852 54462
rect 39340 54402 39396 54404
rect 39340 54350 39342 54402
rect 39342 54350 39394 54402
rect 39394 54350 39396 54402
rect 39340 54348 39396 54350
rect 40460 54402 40516 54404
rect 40460 54350 40462 54402
rect 40462 54350 40514 54402
rect 40514 54350 40516 54402
rect 40460 54348 40516 54350
rect 39228 53788 39284 53844
rect 39340 53730 39396 53732
rect 39340 53678 39342 53730
rect 39342 53678 39394 53730
rect 39394 53678 39396 53730
rect 39340 53676 39396 53678
rect 40348 53730 40404 53732
rect 40348 53678 40350 53730
rect 40350 53678 40402 53730
rect 40402 53678 40404 53730
rect 40348 53676 40404 53678
rect 40460 53618 40516 53620
rect 40460 53566 40462 53618
rect 40462 53566 40514 53618
rect 40514 53566 40516 53618
rect 40460 53564 40516 53566
rect 40908 53170 40964 53172
rect 40908 53118 40910 53170
rect 40910 53118 40962 53170
rect 40962 53118 40964 53170
rect 40908 53116 40964 53118
rect 38892 51884 38948 51940
rect 38780 51212 38836 51268
rect 38220 50540 38276 50596
rect 38668 50428 38724 50484
rect 38332 48188 38388 48244
rect 38108 47628 38164 47684
rect 37660 47292 37716 47348
rect 37548 46844 37604 46900
rect 37772 47180 37828 47236
rect 37996 46620 38052 46676
rect 38668 47404 38724 47460
rect 37436 45666 37492 45668
rect 37436 45614 37438 45666
rect 37438 45614 37490 45666
rect 37490 45614 37492 45666
rect 37436 45612 37492 45614
rect 37660 46060 37716 46116
rect 38332 46060 38388 46116
rect 37772 45890 37828 45892
rect 37772 45838 37774 45890
rect 37774 45838 37826 45890
rect 37826 45838 37828 45890
rect 37772 45836 37828 45838
rect 39116 52162 39172 52164
rect 39116 52110 39118 52162
rect 39118 52110 39170 52162
rect 39170 52110 39172 52162
rect 39116 52108 39172 52110
rect 39004 51548 39060 51604
rect 39004 50316 39060 50372
rect 38892 49698 38948 49700
rect 38892 49646 38894 49698
rect 38894 49646 38946 49698
rect 38946 49646 38948 49698
rect 38892 49644 38948 49646
rect 39788 52668 39844 52724
rect 39340 51266 39396 51268
rect 39340 51214 39342 51266
rect 39342 51214 39394 51266
rect 39394 51214 39396 51266
rect 39340 51212 39396 51214
rect 39228 50482 39284 50484
rect 39228 50430 39230 50482
rect 39230 50430 39282 50482
rect 39282 50430 39284 50482
rect 39228 50428 39284 50430
rect 40460 52274 40516 52276
rect 40460 52222 40462 52274
rect 40462 52222 40514 52274
rect 40514 52222 40516 52274
rect 40460 52220 40516 52222
rect 40348 51996 40404 52052
rect 40124 51378 40180 51380
rect 40124 51326 40126 51378
rect 40126 51326 40178 51378
rect 40178 51326 40180 51378
rect 40124 51324 40180 51326
rect 39788 50876 39844 50932
rect 40012 51212 40068 51268
rect 39340 49698 39396 49700
rect 39340 49646 39342 49698
rect 39342 49646 39394 49698
rect 39394 49646 39396 49698
rect 39340 49644 39396 49646
rect 39228 49026 39284 49028
rect 39228 48974 39230 49026
rect 39230 48974 39282 49026
rect 39282 48974 39284 49026
rect 39228 48972 39284 48974
rect 38780 45836 38836 45892
rect 39116 45890 39172 45892
rect 39116 45838 39118 45890
rect 39118 45838 39170 45890
rect 39170 45838 39172 45890
rect 39116 45836 39172 45838
rect 39676 50204 39732 50260
rect 39788 50316 39844 50372
rect 40908 52556 40964 52612
rect 39900 50204 39956 50260
rect 39452 48748 39508 48804
rect 39900 49644 39956 49700
rect 40012 49308 40068 49364
rect 40684 49868 40740 49924
rect 40460 49698 40516 49700
rect 40460 49646 40462 49698
rect 40462 49646 40514 49698
rect 40514 49646 40516 49698
rect 40460 49644 40516 49646
rect 39788 48972 39844 49028
rect 40012 48860 40068 48916
rect 40236 48972 40292 49028
rect 40124 48076 40180 48132
rect 39452 47852 39508 47908
rect 40460 49308 40516 49364
rect 40348 48242 40404 48244
rect 40348 48190 40350 48242
rect 40350 48190 40402 48242
rect 40402 48190 40404 48242
rect 40348 48188 40404 48190
rect 40684 49026 40740 49028
rect 40684 48974 40686 49026
rect 40686 48974 40738 49026
rect 40738 48974 40740 49026
rect 40684 48972 40740 48974
rect 41020 51324 41076 51380
rect 41020 50428 41076 50484
rect 41132 50540 41188 50596
rect 42476 55970 42532 55972
rect 42476 55918 42478 55970
rect 42478 55918 42530 55970
rect 42530 55918 42532 55970
rect 42476 55916 42532 55918
rect 42924 55916 42980 55972
rect 46956 56028 47012 56084
rect 41580 54460 41636 54516
rect 41580 53788 41636 53844
rect 42140 54626 42196 54628
rect 42140 54574 42142 54626
rect 42142 54574 42194 54626
rect 42194 54574 42196 54626
rect 42140 54572 42196 54574
rect 42252 54402 42308 54404
rect 42252 54350 42254 54402
rect 42254 54350 42306 54402
rect 42306 54350 42308 54402
rect 42252 54348 42308 54350
rect 42476 54348 42532 54404
rect 42476 53340 42532 53396
rect 43708 55298 43764 55300
rect 43708 55246 43710 55298
rect 43710 55246 43762 55298
rect 43762 55246 43764 55298
rect 43708 55244 43764 55246
rect 44156 55186 44212 55188
rect 44156 55134 44158 55186
rect 44158 55134 44210 55186
rect 44210 55134 44212 55186
rect 44156 55132 44212 55134
rect 46620 55186 46676 55188
rect 46620 55134 46622 55186
rect 46622 55134 46674 55186
rect 46674 55134 46676 55186
rect 46620 55132 46676 55134
rect 50556 56474 50612 56476
rect 50556 56422 50558 56474
rect 50558 56422 50610 56474
rect 50610 56422 50612 56474
rect 50556 56420 50612 56422
rect 50660 56474 50716 56476
rect 50660 56422 50662 56474
rect 50662 56422 50714 56474
rect 50714 56422 50716 56474
rect 50660 56420 50716 56422
rect 50764 56474 50820 56476
rect 50764 56422 50766 56474
rect 50766 56422 50818 56474
rect 50818 56422 50820 56474
rect 50764 56420 50820 56422
rect 54236 56194 54292 56196
rect 54236 56142 54238 56194
rect 54238 56142 54290 56194
rect 54290 56142 54292 56194
rect 54236 56140 54292 56142
rect 48860 56082 48916 56084
rect 48860 56030 48862 56082
rect 48862 56030 48914 56082
rect 48914 56030 48916 56082
rect 48860 56028 48916 56030
rect 48412 55916 48468 55972
rect 49532 55970 49588 55972
rect 49532 55918 49534 55970
rect 49534 55918 49586 55970
rect 49586 55918 49588 55970
rect 49532 55916 49588 55918
rect 54684 56140 54740 56196
rect 57820 56194 57876 56196
rect 57820 56142 57822 56194
rect 57822 56142 57874 56194
rect 57874 56142 57876 56194
rect 57820 56140 57876 56142
rect 59836 56140 59892 56196
rect 54460 55916 54516 55972
rect 55468 55970 55524 55972
rect 55468 55918 55470 55970
rect 55470 55918 55522 55970
rect 55522 55918 55524 55970
rect 55468 55916 55524 55918
rect 49308 55580 49364 55636
rect 43708 54572 43764 54628
rect 42028 52556 42084 52612
rect 42028 52386 42084 52388
rect 42028 52334 42030 52386
rect 42030 52334 42082 52386
rect 42082 52334 42084 52386
rect 42028 52332 42084 52334
rect 41468 51996 41524 52052
rect 42140 52220 42196 52276
rect 41356 51884 41412 51940
rect 41468 51490 41524 51492
rect 41468 51438 41470 51490
rect 41470 51438 41522 51490
rect 41522 51438 41524 51490
rect 41468 51436 41524 51438
rect 42028 51266 42084 51268
rect 42028 51214 42030 51266
rect 42030 51214 42082 51266
rect 42082 51214 42084 51266
rect 42028 51212 42084 51214
rect 39676 47458 39732 47460
rect 39676 47406 39678 47458
rect 39678 47406 39730 47458
rect 39730 47406 39732 47458
rect 39676 47404 39732 47406
rect 40236 47068 40292 47124
rect 39340 45836 39396 45892
rect 37660 45500 37716 45556
rect 38780 45666 38836 45668
rect 38780 45614 38782 45666
rect 38782 45614 38834 45666
rect 38834 45614 38836 45666
rect 38780 45612 38836 45614
rect 38220 45388 38276 45444
rect 36652 43820 36708 43876
rect 37436 43372 37492 43428
rect 36652 42866 36708 42868
rect 36652 42814 36654 42866
rect 36654 42814 36706 42866
rect 36706 42814 36708 42866
rect 36652 42812 36708 42814
rect 36764 42700 36820 42756
rect 36540 40236 36596 40292
rect 36652 42476 36708 42532
rect 36652 42252 36708 42308
rect 36652 40012 36708 40068
rect 36540 39676 36596 39732
rect 35644 39452 35700 39508
rect 35644 39228 35700 39284
rect 34860 38162 34916 38164
rect 34860 38110 34862 38162
rect 34862 38110 34914 38162
rect 34914 38110 34916 38162
rect 34860 38108 34916 38110
rect 34860 37938 34916 37940
rect 34860 37886 34862 37938
rect 34862 37886 34914 37938
rect 34914 37886 34916 37938
rect 34860 37884 34916 37886
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35084 37826 35140 37828
rect 35084 37774 35086 37826
rect 35086 37774 35138 37826
rect 35138 37774 35140 37826
rect 35084 37772 35140 37774
rect 34748 35586 34804 35588
rect 34748 35534 34750 35586
rect 34750 35534 34802 35586
rect 34802 35534 34804 35586
rect 34748 35532 34804 35534
rect 34524 31948 34580 32004
rect 34636 33292 34692 33348
rect 34188 30882 34244 30884
rect 34188 30830 34190 30882
rect 34190 30830 34242 30882
rect 34242 30830 34244 30882
rect 34188 30828 34244 30830
rect 34300 30940 34356 30996
rect 33852 30044 33908 30100
rect 34188 30098 34244 30100
rect 34188 30046 34190 30098
rect 34190 30046 34242 30098
rect 34242 30046 34244 30098
rect 34188 30044 34244 30046
rect 33740 29820 33796 29876
rect 33964 28754 34020 28756
rect 33964 28702 33966 28754
rect 33966 28702 34018 28754
rect 34018 28702 34020 28754
rect 33964 28700 34020 28702
rect 33516 28642 33572 28644
rect 33516 28590 33518 28642
rect 33518 28590 33570 28642
rect 33570 28590 33572 28642
rect 33516 28588 33572 28590
rect 33180 26850 33236 26852
rect 33180 26798 33182 26850
rect 33182 26798 33234 26850
rect 33234 26798 33236 26850
rect 33180 26796 33236 26798
rect 33180 24556 33236 24612
rect 33628 28140 33684 28196
rect 33516 26178 33572 26180
rect 33516 26126 33518 26178
rect 33518 26126 33570 26178
rect 33570 26126 33572 26178
rect 33516 26124 33572 26126
rect 33404 26012 33460 26068
rect 33516 25452 33572 25508
rect 33404 25282 33460 25284
rect 33404 25230 33406 25282
rect 33406 25230 33458 25282
rect 33458 25230 33460 25282
rect 33404 25228 33460 25230
rect 33292 23996 33348 24052
rect 33404 24892 33460 24948
rect 33292 23826 33348 23828
rect 33292 23774 33294 23826
rect 33294 23774 33346 23826
rect 33346 23774 33348 23826
rect 33292 23772 33348 23774
rect 33516 24444 33572 24500
rect 33852 28028 33908 28084
rect 34076 28028 34132 28084
rect 33964 26124 34020 26180
rect 33740 24780 33796 24836
rect 33852 24444 33908 24500
rect 33516 23826 33572 23828
rect 33516 23774 33518 23826
rect 33518 23774 33570 23826
rect 33570 23774 33572 23826
rect 33516 23772 33572 23774
rect 33628 23548 33684 23604
rect 33068 23324 33124 23380
rect 32844 23212 32900 23268
rect 32956 22876 33012 22932
rect 32732 21980 32788 22036
rect 32844 22092 32900 22148
rect 33180 22146 33236 22148
rect 33180 22094 33182 22146
rect 33182 22094 33234 22146
rect 33234 22094 33236 22146
rect 33180 22092 33236 22094
rect 32508 20524 32564 20580
rect 32508 19010 32564 19012
rect 32508 18958 32510 19010
rect 32510 18958 32562 19010
rect 32562 18958 32564 19010
rect 32508 18956 32564 18958
rect 32508 18732 32564 18788
rect 32620 18620 32676 18676
rect 32732 18172 32788 18228
rect 32732 17388 32788 17444
rect 32732 16940 32788 16996
rect 32508 16882 32564 16884
rect 32508 16830 32510 16882
rect 32510 16830 32562 16882
rect 32562 16830 32564 16882
rect 32508 16828 32564 16830
rect 31724 15538 31780 15540
rect 31724 15486 31726 15538
rect 31726 15486 31778 15538
rect 31778 15486 31780 15538
rect 31724 15484 31780 15486
rect 32508 15538 32564 15540
rect 32508 15486 32510 15538
rect 32510 15486 32562 15538
rect 32562 15486 32564 15538
rect 32508 15484 32564 15486
rect 31388 13634 31444 13636
rect 31388 13582 31390 13634
rect 31390 13582 31442 13634
rect 31442 13582 31444 13634
rect 31388 13580 31444 13582
rect 31276 12962 31332 12964
rect 31276 12910 31278 12962
rect 31278 12910 31330 12962
rect 31330 12910 31332 12962
rect 31276 12908 31332 12910
rect 31164 12290 31220 12292
rect 31164 12238 31166 12290
rect 31166 12238 31218 12290
rect 31218 12238 31220 12290
rect 31164 12236 31220 12238
rect 31724 14028 31780 14084
rect 32284 15314 32340 15316
rect 32284 15262 32286 15314
rect 32286 15262 32338 15314
rect 32338 15262 32340 15314
rect 32284 15260 32340 15262
rect 31948 13468 32004 13524
rect 31500 10556 31556 10612
rect 31052 5180 31108 5236
rect 33180 20412 33236 20468
rect 33628 23324 33684 23380
rect 33516 23266 33572 23268
rect 33516 23214 33518 23266
rect 33518 23214 33570 23266
rect 33570 23214 33572 23266
rect 33516 23212 33572 23214
rect 33516 22258 33572 22260
rect 33516 22206 33518 22258
rect 33518 22206 33570 22258
rect 33570 22206 33572 22258
rect 33516 22204 33572 22206
rect 33964 23548 34020 23604
rect 34972 33516 35028 33572
rect 34860 31778 34916 31780
rect 34860 31726 34862 31778
rect 34862 31726 34914 31778
rect 34914 31726 34916 31778
rect 34860 31724 34916 31726
rect 34748 30828 34804 30884
rect 34748 30268 34804 30324
rect 34412 30044 34468 30100
rect 34524 29932 34580 29988
rect 34188 27298 34244 27300
rect 34188 27246 34190 27298
rect 34190 27246 34242 27298
rect 34242 27246 34244 27298
rect 34188 27244 34244 27246
rect 33404 21644 33460 21700
rect 33404 20860 33460 20916
rect 33628 20578 33684 20580
rect 33628 20526 33630 20578
rect 33630 20526 33682 20578
rect 33682 20526 33684 20578
rect 33628 20524 33684 20526
rect 33628 20300 33684 20356
rect 32956 19740 33012 19796
rect 32956 19234 33012 19236
rect 32956 19182 32958 19234
rect 32958 19182 33010 19234
rect 33010 19182 33012 19234
rect 32956 19180 33012 19182
rect 33068 17724 33124 17780
rect 33404 17724 33460 17780
rect 33180 17442 33236 17444
rect 33180 17390 33182 17442
rect 33182 17390 33234 17442
rect 33234 17390 33236 17442
rect 33180 17388 33236 17390
rect 33068 17276 33124 17332
rect 32956 15986 33012 15988
rect 32956 15934 32958 15986
rect 32958 15934 33010 15986
rect 33010 15934 33012 15986
rect 32956 15932 33012 15934
rect 32956 15314 33012 15316
rect 32956 15262 32958 15314
rect 32958 15262 33010 15314
rect 33010 15262 33012 15314
rect 32956 15260 33012 15262
rect 32844 12908 32900 12964
rect 32396 5180 32452 5236
rect 32844 12236 32900 12292
rect 31052 4060 31108 4116
rect 30492 3554 30548 3556
rect 30492 3502 30494 3554
rect 30494 3502 30546 3554
rect 30546 3502 30548 3554
rect 30492 3500 30548 3502
rect 31052 3500 31108 3556
rect 29372 3442 29428 3444
rect 29372 3390 29374 3442
rect 29374 3390 29426 3442
rect 29426 3390 29428 3442
rect 29372 3388 29428 3390
rect 33292 12796 33348 12852
rect 33068 11340 33124 11396
rect 34076 21868 34132 21924
rect 34188 25340 34244 25396
rect 34076 21698 34132 21700
rect 34076 21646 34078 21698
rect 34078 21646 34130 21698
rect 34130 21646 34132 21698
rect 34076 21644 34132 21646
rect 33964 21586 34020 21588
rect 33964 21534 33966 21586
rect 33966 21534 34018 21586
rect 34018 21534 34020 21586
rect 33964 21532 34020 21534
rect 34524 28530 34580 28532
rect 34524 28478 34526 28530
rect 34526 28478 34578 28530
rect 34578 28478 34580 28530
rect 34524 28476 34580 28478
rect 34748 28924 34804 28980
rect 34748 28588 34804 28644
rect 34636 27916 34692 27972
rect 34412 26962 34468 26964
rect 34412 26910 34414 26962
rect 34414 26910 34466 26962
rect 34466 26910 34468 26962
rect 34412 26908 34468 26910
rect 34524 27244 34580 27300
rect 34412 26124 34468 26180
rect 34972 31500 35028 31556
rect 34972 30882 35028 30884
rect 34972 30830 34974 30882
rect 34974 30830 35026 30882
rect 35026 30830 35028 30882
rect 34972 30828 35028 30830
rect 35644 37884 35700 37940
rect 35756 37042 35812 37044
rect 35756 36990 35758 37042
rect 35758 36990 35810 37042
rect 35810 36990 35812 37042
rect 35756 36988 35812 36990
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36204 38220 36260 38276
rect 35980 37660 36036 37716
rect 35308 35698 35364 35700
rect 35308 35646 35310 35698
rect 35310 35646 35362 35698
rect 35362 35646 35364 35698
rect 35308 35644 35364 35646
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35308 33516 35364 33572
rect 36652 39506 36708 39508
rect 36652 39454 36654 39506
rect 36654 39454 36706 39506
rect 36706 39454 36708 39506
rect 36652 39452 36708 39454
rect 37660 42754 37716 42756
rect 37660 42702 37662 42754
rect 37662 42702 37714 42754
rect 37714 42702 37716 42754
rect 37660 42700 37716 42702
rect 37212 42588 37268 42644
rect 36988 42194 37044 42196
rect 36988 42142 36990 42194
rect 36990 42142 37042 42194
rect 37042 42142 37044 42194
rect 36988 42140 37044 42142
rect 37100 41970 37156 41972
rect 37100 41918 37102 41970
rect 37102 41918 37154 41970
rect 37154 41918 37156 41970
rect 37100 41916 37156 41918
rect 36876 41244 36932 41300
rect 36876 40626 36932 40628
rect 36876 40574 36878 40626
rect 36878 40574 36930 40626
rect 36930 40574 36932 40626
rect 36876 40572 36932 40574
rect 36204 37660 36260 37716
rect 36540 37938 36596 37940
rect 36540 37886 36542 37938
rect 36542 37886 36594 37938
rect 36594 37886 36596 37938
rect 36540 37884 36596 37886
rect 36204 36988 36260 37044
rect 36092 34524 36148 34580
rect 35868 33628 35924 33684
rect 35532 32562 35588 32564
rect 35532 32510 35534 32562
rect 35534 32510 35586 32562
rect 35586 32510 35588 32562
rect 35532 32508 35588 32510
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35308 30940 35364 30996
rect 35420 31500 35476 31556
rect 35532 31388 35588 31444
rect 35868 31948 35924 32004
rect 35756 31778 35812 31780
rect 35756 31726 35758 31778
rect 35758 31726 35810 31778
rect 35810 31726 35812 31778
rect 35756 31724 35812 31726
rect 35420 30716 35476 30772
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35084 30044 35140 30100
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35644 30994 35700 30996
rect 35644 30942 35646 30994
rect 35646 30942 35698 30994
rect 35698 30942 35700 30994
rect 35644 30940 35700 30942
rect 35756 30156 35812 30212
rect 35644 30098 35700 30100
rect 35644 30046 35646 30098
rect 35646 30046 35698 30098
rect 35698 30046 35700 30098
rect 35644 30044 35700 30046
rect 35644 29820 35700 29876
rect 35084 28812 35140 28868
rect 35196 28700 35252 28756
rect 35084 28476 35140 28532
rect 34972 27916 35028 27972
rect 35644 28700 35700 28756
rect 35868 28642 35924 28644
rect 35868 28590 35870 28642
rect 35870 28590 35922 28642
rect 35922 28590 35924 28642
rect 35868 28588 35924 28590
rect 35868 28364 35924 28420
rect 35532 27970 35588 27972
rect 35532 27918 35534 27970
rect 35534 27918 35586 27970
rect 35586 27918 35588 27970
rect 35532 27916 35588 27918
rect 35756 27916 35812 27972
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 27020 35252 27076
rect 34412 25506 34468 25508
rect 34412 25454 34414 25506
rect 34414 25454 34466 25506
rect 34466 25454 34468 25506
rect 34412 25452 34468 25454
rect 34300 24892 34356 24948
rect 34412 24834 34468 24836
rect 34412 24782 34414 24834
rect 34414 24782 34466 24834
rect 34466 24782 34468 24834
rect 34412 24780 34468 24782
rect 34636 24780 34692 24836
rect 34860 25340 34916 25396
rect 35420 26796 35476 26852
rect 35644 26684 35700 26740
rect 35420 26572 35476 26628
rect 35532 26348 35588 26404
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35084 25228 35140 25284
rect 34748 24556 34804 24612
rect 34300 23826 34356 23828
rect 34300 23774 34302 23826
rect 34302 23774 34354 23826
rect 34354 23774 34356 23826
rect 34300 23772 34356 23774
rect 34636 23826 34692 23828
rect 34636 23774 34638 23826
rect 34638 23774 34690 23826
rect 34690 23774 34692 23826
rect 34636 23772 34692 23774
rect 34300 23548 34356 23604
rect 34524 23548 34580 23604
rect 34636 23042 34692 23044
rect 34636 22990 34638 23042
rect 34638 22990 34690 23042
rect 34690 22990 34692 23042
rect 34636 22988 34692 22990
rect 34524 22876 34580 22932
rect 34748 22540 34804 22596
rect 35532 25676 35588 25732
rect 35644 26290 35700 26292
rect 35644 26238 35646 26290
rect 35646 26238 35698 26290
rect 35698 26238 35700 26290
rect 35644 26236 35700 26238
rect 36316 35868 36372 35924
rect 36428 35810 36484 35812
rect 36428 35758 36430 35810
rect 36430 35758 36482 35810
rect 36482 35758 36484 35810
rect 36428 35756 36484 35758
rect 36316 33852 36372 33908
rect 36316 33628 36372 33684
rect 36092 32508 36148 32564
rect 36204 32060 36260 32116
rect 36092 29202 36148 29204
rect 36092 29150 36094 29202
rect 36094 29150 36146 29202
rect 36146 29150 36148 29202
rect 36092 29148 36148 29150
rect 36092 28700 36148 28756
rect 36428 32562 36484 32564
rect 36428 32510 36430 32562
rect 36430 32510 36482 32562
rect 36482 32510 36484 32562
rect 36428 32508 36484 32510
rect 36428 31948 36484 32004
rect 36540 31836 36596 31892
rect 38556 45052 38612 45108
rect 37996 43708 38052 43764
rect 37884 42476 37940 42532
rect 37772 41970 37828 41972
rect 37772 41918 37774 41970
rect 37774 41918 37826 41970
rect 37826 41918 37828 41970
rect 37772 41916 37828 41918
rect 37324 40124 37380 40180
rect 37548 39340 37604 39396
rect 36764 38834 36820 38836
rect 36764 38782 36766 38834
rect 36766 38782 36818 38834
rect 36818 38782 36820 38834
rect 36764 38780 36820 38782
rect 36764 38274 36820 38276
rect 36764 38222 36766 38274
rect 36766 38222 36818 38274
rect 36818 38222 36820 38274
rect 36764 38220 36820 38222
rect 38444 43708 38500 43764
rect 38668 44604 38724 44660
rect 38780 43932 38836 43988
rect 38892 43260 38948 43316
rect 38332 42700 38388 42756
rect 38556 42700 38612 42756
rect 38220 42642 38276 42644
rect 38220 42590 38222 42642
rect 38222 42590 38274 42642
rect 38274 42590 38276 42642
rect 38220 42588 38276 42590
rect 38108 42252 38164 42308
rect 39116 44098 39172 44100
rect 39116 44046 39118 44098
rect 39118 44046 39170 44098
rect 39170 44046 39172 44098
rect 39116 44044 39172 44046
rect 39004 42588 39060 42644
rect 38892 42476 38948 42532
rect 38892 42194 38948 42196
rect 38892 42142 38894 42194
rect 38894 42142 38946 42194
rect 38946 42142 38948 42194
rect 38892 42140 38948 42142
rect 38892 41916 38948 41972
rect 37884 41298 37940 41300
rect 37884 41246 37886 41298
rect 37886 41246 37938 41298
rect 37938 41246 37940 41298
rect 37884 41244 37940 41246
rect 38108 41132 38164 41188
rect 37772 39788 37828 39844
rect 37772 39506 37828 39508
rect 37772 39454 37774 39506
rect 37774 39454 37826 39506
rect 37826 39454 37828 39506
rect 37772 39452 37828 39454
rect 37884 39394 37940 39396
rect 37884 39342 37886 39394
rect 37886 39342 37938 39394
rect 37938 39342 37940 39394
rect 37884 39340 37940 39342
rect 37660 38780 37716 38836
rect 37436 38668 37492 38724
rect 39564 46620 39620 46676
rect 40012 46620 40068 46676
rect 40684 48076 40740 48132
rect 40684 47068 40740 47124
rect 40684 46898 40740 46900
rect 40684 46846 40686 46898
rect 40686 46846 40738 46898
rect 40738 46846 40740 46898
rect 40684 46844 40740 46846
rect 40796 46732 40852 46788
rect 40572 46674 40628 46676
rect 40572 46622 40574 46674
rect 40574 46622 40626 46674
rect 40626 46622 40628 46674
rect 40572 46620 40628 46622
rect 40348 46508 40404 46564
rect 39564 45106 39620 45108
rect 39564 45054 39566 45106
rect 39566 45054 39618 45106
rect 39618 45054 39620 45106
rect 39564 45052 39620 45054
rect 39676 44492 39732 44548
rect 39676 43708 39732 43764
rect 39340 43372 39396 43428
rect 39452 43260 39508 43316
rect 39452 42700 39508 42756
rect 39340 42588 39396 42644
rect 38892 41186 38948 41188
rect 38892 41134 38894 41186
rect 38894 41134 38946 41186
rect 38946 41134 38948 41186
rect 38892 41132 38948 41134
rect 39116 41074 39172 41076
rect 39116 41022 39118 41074
rect 39118 41022 39170 41074
rect 39170 41022 39172 41074
rect 39116 41020 39172 41022
rect 38332 40908 38388 40964
rect 38220 40514 38276 40516
rect 38220 40462 38222 40514
rect 38222 40462 38274 40514
rect 38274 40462 38276 40514
rect 38220 40460 38276 40462
rect 39116 40626 39172 40628
rect 39116 40574 39118 40626
rect 39118 40574 39170 40626
rect 39170 40574 39172 40626
rect 39116 40572 39172 40574
rect 38332 39788 38388 39844
rect 38668 39730 38724 39732
rect 38668 39678 38670 39730
rect 38670 39678 38722 39730
rect 38722 39678 38724 39730
rect 38668 39676 38724 39678
rect 39340 39900 39396 39956
rect 39004 39676 39060 39732
rect 38556 39452 38612 39508
rect 38332 39004 38388 39060
rect 38444 39340 38500 39396
rect 39004 39228 39060 39284
rect 40348 46060 40404 46116
rect 40908 48188 40964 48244
rect 40908 47628 40964 47684
rect 41244 48188 41300 48244
rect 41020 46956 41076 47012
rect 41132 46620 41188 46676
rect 40908 46508 40964 46564
rect 40796 46060 40852 46116
rect 40460 45836 40516 45892
rect 40236 44492 40292 44548
rect 39900 42924 39956 42980
rect 39788 42812 39844 42868
rect 39676 42754 39732 42756
rect 39676 42702 39678 42754
rect 39678 42702 39730 42754
rect 39730 42702 39732 42754
rect 39676 42700 39732 42702
rect 40012 42252 40068 42308
rect 39900 41970 39956 41972
rect 39900 41918 39902 41970
rect 39902 41918 39954 41970
rect 39954 41918 39956 41970
rect 39900 41916 39956 41918
rect 40236 43426 40292 43428
rect 40236 43374 40238 43426
rect 40238 43374 40290 43426
rect 40290 43374 40292 43426
rect 40236 43372 40292 43374
rect 40236 42978 40292 42980
rect 40236 42926 40238 42978
rect 40238 42926 40290 42978
rect 40290 42926 40292 42978
rect 40236 42924 40292 42926
rect 39676 41074 39732 41076
rect 39676 41022 39678 41074
rect 39678 41022 39730 41074
rect 39730 41022 39732 41074
rect 39676 41020 39732 41022
rect 39564 40908 39620 40964
rect 40460 42812 40516 42868
rect 40348 41916 40404 41972
rect 41132 45052 41188 45108
rect 40684 44828 40740 44884
rect 40908 44940 40964 44996
rect 40684 44098 40740 44100
rect 40684 44046 40686 44098
rect 40686 44046 40738 44098
rect 40738 44046 40740 44098
rect 40684 44044 40740 44046
rect 40796 43538 40852 43540
rect 40796 43486 40798 43538
rect 40798 43486 40850 43538
rect 40850 43486 40852 43538
rect 40796 43484 40852 43486
rect 40684 43260 40740 43316
rect 40684 42754 40740 42756
rect 40684 42702 40686 42754
rect 40686 42702 40738 42754
rect 40738 42702 40740 42754
rect 40684 42700 40740 42702
rect 40684 42028 40740 42084
rect 40124 41020 40180 41076
rect 40236 41468 40292 41524
rect 40012 40908 40068 40964
rect 37772 38050 37828 38052
rect 37772 37998 37774 38050
rect 37774 37998 37826 38050
rect 37826 37998 37828 38050
rect 37772 37996 37828 37998
rect 37212 37884 37268 37940
rect 36876 37772 36932 37828
rect 36988 37660 37044 37716
rect 36764 36988 36820 37044
rect 36988 36764 37044 36820
rect 37436 36764 37492 36820
rect 36988 35922 37044 35924
rect 36988 35870 36990 35922
rect 36990 35870 37042 35922
rect 37042 35870 37044 35922
rect 36988 35868 37044 35870
rect 37436 35810 37492 35812
rect 37436 35758 37438 35810
rect 37438 35758 37490 35810
rect 37490 35758 37492 35810
rect 37436 35756 37492 35758
rect 37100 35644 37156 35700
rect 36988 34636 37044 34692
rect 36764 33852 36820 33908
rect 36876 33068 36932 33124
rect 36988 32060 37044 32116
rect 36988 31836 37044 31892
rect 36316 31554 36372 31556
rect 36316 31502 36318 31554
rect 36318 31502 36370 31554
rect 36370 31502 36372 31554
rect 36316 31500 36372 31502
rect 36540 31388 36596 31444
rect 36540 29820 36596 29876
rect 36764 29596 36820 29652
rect 36540 28588 36596 28644
rect 36764 28700 36820 28756
rect 36204 27580 36260 27636
rect 36764 27858 36820 27860
rect 36764 27806 36766 27858
rect 36766 27806 36818 27858
rect 36818 27806 36820 27858
rect 36764 27804 36820 27806
rect 36988 29036 37044 29092
rect 36652 27244 36708 27300
rect 36764 27580 36820 27636
rect 36540 27132 36596 27188
rect 36540 26908 36596 26964
rect 35980 26572 36036 26628
rect 36540 26572 36596 26628
rect 35868 25676 35924 25732
rect 35644 24668 35700 24724
rect 34188 21196 34244 21252
rect 35532 24610 35588 24612
rect 35532 24558 35534 24610
rect 35534 24558 35586 24610
rect 35586 24558 35588 24610
rect 35532 24556 35588 24558
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35980 24834 36036 24836
rect 35980 24782 35982 24834
rect 35982 24782 36034 24834
rect 36034 24782 36036 24834
rect 35980 24780 36036 24782
rect 35756 23324 35812 23380
rect 35532 22876 35588 22932
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 34412 21532 34468 21588
rect 34412 20860 34468 20916
rect 34524 21868 34580 21924
rect 33852 19740 33908 19796
rect 33740 18226 33796 18228
rect 33740 18174 33742 18226
rect 33742 18174 33794 18226
rect 33794 18174 33796 18226
rect 33740 18172 33796 18174
rect 33740 17724 33796 17780
rect 33516 16828 33572 16884
rect 33964 17778 34020 17780
rect 33964 17726 33966 17778
rect 33966 17726 34018 17778
rect 34018 17726 34020 17778
rect 33964 17724 34020 17726
rect 33852 17500 33908 17556
rect 33516 16604 33572 16660
rect 33964 17106 34020 17108
rect 33964 17054 33966 17106
rect 33966 17054 34018 17106
rect 34018 17054 34020 17106
rect 33964 17052 34020 17054
rect 34300 18396 34356 18452
rect 34412 18284 34468 18340
rect 34524 19964 34580 20020
rect 34300 18226 34356 18228
rect 34300 18174 34302 18226
rect 34302 18174 34354 18226
rect 34354 18174 34356 18226
rect 34300 18172 34356 18174
rect 34188 17836 34244 17892
rect 34412 16994 34468 16996
rect 34412 16942 34414 16994
rect 34414 16942 34466 16994
rect 34466 16942 34468 16994
rect 34412 16940 34468 16942
rect 33740 15538 33796 15540
rect 33740 15486 33742 15538
rect 33742 15486 33794 15538
rect 33794 15486 33796 15538
rect 33740 15484 33796 15486
rect 33516 15314 33572 15316
rect 33516 15262 33518 15314
rect 33518 15262 33570 15314
rect 33570 15262 33572 15314
rect 33516 15260 33572 15262
rect 33404 8092 33460 8148
rect 33516 14252 33572 14308
rect 33628 13970 33684 13972
rect 33628 13918 33630 13970
rect 33630 13918 33682 13970
rect 33682 13918 33684 13970
rect 33628 13916 33684 13918
rect 34972 21980 35028 22036
rect 34860 20300 34916 20356
rect 34748 19740 34804 19796
rect 34748 19234 34804 19236
rect 34748 19182 34750 19234
rect 34750 19182 34802 19234
rect 34802 19182 34804 19234
rect 34748 19180 34804 19182
rect 34860 19122 34916 19124
rect 34860 19070 34862 19122
rect 34862 19070 34914 19122
rect 34914 19070 34916 19122
rect 34860 19068 34916 19070
rect 35420 21420 35476 21476
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35420 20972 35476 21028
rect 35308 20412 35364 20468
rect 35196 20300 35252 20356
rect 35756 22594 35812 22596
rect 35756 22542 35758 22594
rect 35758 22542 35810 22594
rect 35810 22542 35812 22594
rect 35756 22540 35812 22542
rect 35644 22092 35700 22148
rect 35756 21362 35812 21364
rect 35756 21310 35758 21362
rect 35758 21310 35810 21362
rect 35810 21310 35812 21362
rect 35756 21308 35812 21310
rect 36204 25788 36260 25844
rect 36204 25452 36260 25508
rect 36428 26290 36484 26292
rect 36428 26238 36430 26290
rect 36430 26238 36482 26290
rect 36482 26238 36484 26290
rect 36428 26236 36484 26238
rect 36428 25506 36484 25508
rect 36428 25454 36430 25506
rect 36430 25454 36482 25506
rect 36482 25454 36484 25506
rect 36428 25452 36484 25454
rect 36764 26348 36820 26404
rect 36652 25564 36708 25620
rect 36652 25116 36708 25172
rect 36540 23714 36596 23716
rect 36540 23662 36542 23714
rect 36542 23662 36594 23714
rect 36594 23662 36596 23714
rect 36540 23660 36596 23662
rect 36428 23548 36484 23604
rect 36316 23436 36372 23492
rect 36092 23154 36148 23156
rect 36092 23102 36094 23154
rect 36094 23102 36146 23154
rect 36146 23102 36148 23154
rect 36092 23100 36148 23102
rect 35980 21756 36036 21812
rect 35868 20972 35924 21028
rect 35980 21586 36036 21588
rect 35980 21534 35982 21586
rect 35982 21534 36034 21586
rect 36034 21534 36036 21586
rect 35980 21532 36036 21534
rect 35532 20412 35588 20468
rect 36428 22370 36484 22372
rect 36428 22318 36430 22370
rect 36430 22318 36482 22370
rect 36482 22318 36484 22370
rect 36428 22316 36484 22318
rect 36204 22146 36260 22148
rect 36204 22094 36206 22146
rect 36206 22094 36258 22146
rect 36258 22094 36260 22146
rect 36204 22092 36260 22094
rect 36764 22876 36820 22932
rect 37436 35532 37492 35588
rect 37548 34748 37604 34804
rect 37548 34524 37604 34580
rect 37548 32956 37604 33012
rect 37436 32620 37492 32676
rect 38332 37996 38388 38052
rect 38556 38668 38612 38724
rect 38332 37772 38388 37828
rect 39228 38722 39284 38724
rect 39228 38670 39230 38722
rect 39230 38670 39282 38722
rect 39282 38670 39284 38722
rect 39228 38668 39284 38670
rect 40012 39452 40068 39508
rect 39900 39394 39956 39396
rect 39900 39342 39902 39394
rect 39902 39342 39954 39394
rect 39954 39342 39956 39394
rect 39900 39340 39956 39342
rect 40460 39676 40516 39732
rect 41244 44716 41300 44772
rect 41244 43708 41300 43764
rect 41132 43596 41188 43652
rect 41020 43372 41076 43428
rect 41692 48914 41748 48916
rect 41692 48862 41694 48914
rect 41694 48862 41746 48914
rect 41746 48862 41748 48914
rect 41692 48860 41748 48862
rect 41692 48188 41748 48244
rect 41580 47852 41636 47908
rect 41468 46562 41524 46564
rect 41468 46510 41470 46562
rect 41470 46510 41522 46562
rect 41522 46510 41524 46562
rect 41468 46508 41524 46510
rect 41692 47404 41748 47460
rect 41804 47068 41860 47124
rect 41692 46508 41748 46564
rect 41692 45836 41748 45892
rect 42588 53116 42644 53172
rect 42700 54236 42756 54292
rect 42812 53842 42868 53844
rect 42812 53790 42814 53842
rect 42814 53790 42866 53842
rect 42866 53790 42868 53842
rect 42812 53788 42868 53790
rect 43260 54514 43316 54516
rect 43260 54462 43262 54514
rect 43262 54462 43314 54514
rect 43314 54462 43316 54514
rect 43260 54460 43316 54462
rect 42924 53676 42980 53732
rect 43148 54348 43204 54404
rect 43820 54348 43876 54404
rect 42700 52834 42756 52836
rect 42700 52782 42702 52834
rect 42702 52782 42754 52834
rect 42754 52782 42756 52834
rect 42700 52780 42756 52782
rect 42812 52386 42868 52388
rect 42812 52334 42814 52386
rect 42814 52334 42866 52386
rect 42866 52334 42868 52386
rect 42812 52332 42868 52334
rect 43036 52332 43092 52388
rect 42252 52162 42308 52164
rect 42252 52110 42254 52162
rect 42254 52110 42306 52162
rect 42306 52110 42308 52162
rect 42252 52108 42308 52110
rect 42588 51884 42644 51940
rect 43596 53452 43652 53508
rect 43372 53228 43428 53284
rect 43932 53676 43988 53732
rect 43820 53340 43876 53396
rect 44380 53506 44436 53508
rect 44380 53454 44382 53506
rect 44382 53454 44434 53506
rect 44434 53454 44436 53506
rect 44380 53452 44436 53454
rect 45388 53452 45444 53508
rect 43932 53228 43988 53284
rect 43708 52274 43764 52276
rect 43708 52222 43710 52274
rect 43710 52222 43762 52274
rect 43762 52222 43764 52274
rect 43708 52220 43764 52222
rect 43260 51548 43316 51604
rect 44380 53116 44436 53172
rect 44156 52274 44212 52276
rect 44156 52222 44158 52274
rect 44158 52222 44210 52274
rect 44210 52222 44212 52274
rect 44156 52220 44212 52222
rect 43932 52108 43988 52164
rect 43820 51490 43876 51492
rect 43820 51438 43822 51490
rect 43822 51438 43874 51490
rect 43874 51438 43876 51490
rect 43820 51436 43876 51438
rect 44380 51324 44436 51380
rect 47068 53170 47124 53172
rect 47068 53118 47070 53170
rect 47070 53118 47122 53170
rect 47122 53118 47124 53170
rect 47068 53116 47124 53118
rect 45948 52386 46004 52388
rect 45948 52334 45950 52386
rect 45950 52334 46002 52386
rect 46002 52334 46004 52386
rect 45948 52332 46004 52334
rect 46060 51938 46116 51940
rect 46060 51886 46062 51938
rect 46062 51886 46114 51938
rect 46114 51886 46116 51938
rect 46060 51884 46116 51886
rect 45052 51660 45108 51716
rect 42252 51212 42308 51268
rect 42700 50988 42756 51044
rect 42476 50876 42532 50932
rect 42700 50594 42756 50596
rect 42700 50542 42702 50594
rect 42702 50542 42754 50594
rect 42754 50542 42756 50594
rect 42700 50540 42756 50542
rect 42476 48748 42532 48804
rect 43260 50428 43316 50484
rect 42364 48130 42420 48132
rect 42364 48078 42366 48130
rect 42366 48078 42418 48130
rect 42418 48078 42420 48130
rect 42364 48076 42420 48078
rect 42700 47964 42756 48020
rect 42028 47628 42084 47684
rect 41916 46956 41972 47012
rect 41804 45052 41860 45108
rect 42252 46396 42308 46452
rect 41580 44380 41636 44436
rect 41468 43596 41524 43652
rect 41580 43260 41636 43316
rect 41132 42530 41188 42532
rect 41132 42478 41134 42530
rect 41134 42478 41186 42530
rect 41186 42478 41188 42530
rect 41132 42476 41188 42478
rect 41356 42530 41412 42532
rect 41356 42478 41358 42530
rect 41358 42478 41410 42530
rect 41410 42478 41412 42530
rect 41356 42476 41412 42478
rect 41244 42140 41300 42196
rect 41020 41298 41076 41300
rect 41020 41246 41022 41298
rect 41022 41246 41074 41298
rect 41074 41246 41076 41298
rect 41020 41244 41076 41246
rect 40908 39564 40964 39620
rect 39004 37938 39060 37940
rect 39004 37886 39006 37938
rect 39006 37886 39058 37938
rect 39058 37886 39060 37938
rect 39004 37884 39060 37886
rect 37996 36370 38052 36372
rect 37996 36318 37998 36370
rect 37998 36318 38050 36370
rect 38050 36318 38052 36370
rect 37996 36316 38052 36318
rect 37772 35756 37828 35812
rect 39564 37490 39620 37492
rect 39564 37438 39566 37490
rect 39566 37438 39618 37490
rect 39618 37438 39620 37490
rect 39564 37436 39620 37438
rect 39900 37212 39956 37268
rect 38780 36988 38836 37044
rect 39676 37100 39732 37156
rect 39004 36876 39060 36932
rect 38780 36428 38836 36484
rect 38108 35644 38164 35700
rect 38220 36316 38276 36372
rect 38668 36258 38724 36260
rect 38668 36206 38670 36258
rect 38670 36206 38722 36258
rect 38722 36206 38724 36258
rect 38668 36204 38724 36206
rect 38556 35980 38612 36036
rect 38220 35810 38276 35812
rect 38220 35758 38222 35810
rect 38222 35758 38274 35810
rect 38274 35758 38276 35810
rect 38220 35756 38276 35758
rect 38444 35698 38500 35700
rect 38444 35646 38446 35698
rect 38446 35646 38498 35698
rect 38498 35646 38500 35698
rect 38444 35644 38500 35646
rect 38668 35532 38724 35588
rect 38892 35698 38948 35700
rect 38892 35646 38894 35698
rect 38894 35646 38946 35698
rect 38946 35646 38948 35698
rect 38892 35644 38948 35646
rect 39676 36482 39732 36484
rect 39676 36430 39678 36482
rect 39678 36430 39730 36482
rect 39730 36430 39732 36482
rect 39676 36428 39732 36430
rect 39116 36204 39172 36260
rect 37212 29708 37268 29764
rect 37772 33628 37828 33684
rect 37436 31778 37492 31780
rect 37436 31726 37438 31778
rect 37438 31726 37490 31778
rect 37490 31726 37492 31778
rect 37436 31724 37492 31726
rect 38108 33628 38164 33684
rect 38444 33516 38500 33572
rect 38108 32450 38164 32452
rect 38108 32398 38110 32450
rect 38110 32398 38162 32450
rect 38162 32398 38164 32450
rect 38108 32396 38164 32398
rect 37660 31554 37716 31556
rect 37660 31502 37662 31554
rect 37662 31502 37714 31554
rect 37714 31502 37716 31554
rect 37660 31500 37716 31502
rect 37996 31388 38052 31444
rect 38556 32956 38612 33012
rect 38444 32620 38500 32676
rect 38444 31724 38500 31780
rect 37548 28754 37604 28756
rect 37548 28702 37550 28754
rect 37550 28702 37602 28754
rect 37602 28702 37604 28754
rect 37548 28700 37604 28702
rect 37212 27580 37268 27636
rect 37436 27804 37492 27860
rect 37772 29596 37828 29652
rect 37884 29484 37940 29540
rect 38556 31836 38612 31892
rect 39004 34748 39060 34804
rect 39004 34524 39060 34580
rect 38892 32508 38948 32564
rect 39228 34914 39284 34916
rect 39228 34862 39230 34914
rect 39230 34862 39282 34914
rect 39282 34862 39284 34914
rect 39228 34860 39284 34862
rect 39564 35698 39620 35700
rect 39564 35646 39566 35698
rect 39566 35646 39618 35698
rect 39618 35646 39620 35698
rect 39564 35644 39620 35646
rect 39340 34524 39396 34580
rect 39788 35532 39844 35588
rect 39900 35196 39956 35252
rect 40572 39228 40628 39284
rect 41692 43148 41748 43204
rect 41916 43762 41972 43764
rect 41916 43710 41918 43762
rect 41918 43710 41970 43762
rect 41970 43710 41972 43762
rect 41916 43708 41972 43710
rect 41804 42866 41860 42868
rect 41804 42814 41806 42866
rect 41806 42814 41858 42866
rect 41858 42814 41860 42866
rect 41804 42812 41860 42814
rect 41580 42476 41636 42532
rect 41692 41804 41748 41860
rect 41580 40962 41636 40964
rect 41580 40910 41582 40962
rect 41582 40910 41634 40962
rect 41634 40910 41636 40962
rect 41580 40908 41636 40910
rect 44044 50540 44100 50596
rect 43596 50034 43652 50036
rect 43596 49982 43598 50034
rect 43598 49982 43650 50034
rect 43650 49982 43652 50034
rect 43596 49980 43652 49982
rect 43372 49644 43428 49700
rect 44716 50428 44772 50484
rect 43932 49420 43988 49476
rect 42924 48076 42980 48132
rect 43820 48802 43876 48804
rect 43820 48750 43822 48802
rect 43822 48750 43874 48802
rect 43874 48750 43876 48802
rect 43820 48748 43876 48750
rect 44380 48748 44436 48804
rect 43596 48636 43652 48692
rect 43036 47852 43092 47908
rect 42812 47068 42868 47124
rect 42924 47404 42980 47460
rect 43036 46674 43092 46676
rect 43036 46622 43038 46674
rect 43038 46622 43090 46674
rect 43090 46622 43092 46674
rect 43036 46620 43092 46622
rect 42252 44044 42308 44100
rect 42364 43820 42420 43876
rect 42140 43372 42196 43428
rect 42476 43372 42532 43428
rect 42812 43708 42868 43764
rect 43036 43372 43092 43428
rect 42812 42754 42868 42756
rect 42812 42702 42814 42754
rect 42814 42702 42866 42754
rect 42866 42702 42868 42754
rect 42812 42700 42868 42702
rect 43260 44380 43316 44436
rect 42476 42028 42532 42084
rect 42812 42252 42868 42308
rect 42252 41804 42308 41860
rect 41916 40908 41972 40964
rect 41580 40402 41636 40404
rect 41580 40350 41582 40402
rect 41582 40350 41634 40402
rect 41634 40350 41636 40402
rect 41580 40348 41636 40350
rect 42700 41186 42756 41188
rect 42700 41134 42702 41186
rect 42702 41134 42754 41186
rect 42754 41134 42756 41186
rect 42700 41132 42756 41134
rect 42252 40348 42308 40404
rect 41692 39730 41748 39732
rect 41692 39678 41694 39730
rect 41694 39678 41746 39730
rect 41746 39678 41748 39730
rect 41692 39676 41748 39678
rect 42924 40572 42980 40628
rect 43036 41356 43092 41412
rect 40124 37436 40180 37492
rect 40460 37212 40516 37268
rect 40796 38274 40852 38276
rect 40796 38222 40798 38274
rect 40798 38222 40850 38274
rect 40850 38222 40852 38274
rect 40796 38220 40852 38222
rect 40908 37324 40964 37380
rect 40796 37154 40852 37156
rect 40796 37102 40798 37154
rect 40798 37102 40850 37154
rect 40850 37102 40852 37154
rect 40796 37100 40852 37102
rect 40572 36540 40628 36596
rect 40572 36370 40628 36372
rect 40572 36318 40574 36370
rect 40574 36318 40626 36370
rect 40626 36318 40628 36370
rect 40572 36316 40628 36318
rect 40348 36204 40404 36260
rect 41020 35532 41076 35588
rect 40236 34860 40292 34916
rect 40348 34524 40404 34580
rect 40012 34242 40068 34244
rect 40012 34190 40014 34242
rect 40014 34190 40066 34242
rect 40066 34190 40068 34242
rect 40012 34188 40068 34190
rect 39900 33852 39956 33908
rect 39228 33122 39284 33124
rect 39228 33070 39230 33122
rect 39230 33070 39282 33122
rect 39282 33070 39284 33122
rect 39228 33068 39284 33070
rect 39788 33180 39844 33236
rect 40012 33346 40068 33348
rect 40012 33294 40014 33346
rect 40014 33294 40066 33346
rect 40066 33294 40068 33346
rect 40012 33292 40068 33294
rect 39676 32844 39732 32900
rect 39452 32786 39508 32788
rect 39452 32734 39454 32786
rect 39454 32734 39506 32786
rect 39506 32734 39508 32786
rect 39452 32732 39508 32734
rect 38668 31500 38724 31556
rect 38556 31276 38612 31332
rect 38444 30492 38500 30548
rect 38668 30716 38724 30772
rect 38108 29932 38164 29988
rect 38444 29932 38500 29988
rect 38332 29650 38388 29652
rect 38332 29598 38334 29650
rect 38334 29598 38386 29650
rect 38386 29598 38388 29650
rect 38332 29596 38388 29598
rect 38220 29538 38276 29540
rect 38220 29486 38222 29538
rect 38222 29486 38274 29538
rect 38274 29486 38276 29538
rect 38220 29484 38276 29486
rect 37996 28924 38052 28980
rect 38556 28924 38612 28980
rect 38556 28588 38612 28644
rect 37884 28028 37940 28084
rect 37548 27692 37604 27748
rect 37772 27580 37828 27636
rect 37324 27132 37380 27188
rect 36988 25564 37044 25620
rect 37436 26124 37492 26180
rect 37100 25228 37156 25284
rect 36988 25004 37044 25060
rect 37212 25116 37268 25172
rect 37324 25004 37380 25060
rect 37212 23884 37268 23940
rect 38556 28364 38612 28420
rect 37996 27356 38052 27412
rect 38444 28028 38500 28084
rect 38668 28028 38724 28084
rect 38556 27580 38612 27636
rect 38668 27804 38724 27860
rect 37884 26962 37940 26964
rect 37884 26910 37886 26962
rect 37886 26910 37938 26962
rect 37938 26910 37940 26962
rect 37884 26908 37940 26910
rect 37996 26402 38052 26404
rect 37996 26350 37998 26402
rect 37998 26350 38050 26402
rect 38050 26350 38052 26402
rect 37996 26348 38052 26350
rect 37996 26124 38052 26180
rect 37772 26012 37828 26068
rect 37660 25900 37716 25956
rect 37660 25676 37716 25732
rect 37772 25506 37828 25508
rect 37772 25454 37774 25506
rect 37774 25454 37826 25506
rect 37826 25454 37828 25506
rect 37772 25452 37828 25454
rect 37660 25228 37716 25284
rect 37548 24722 37604 24724
rect 37548 24670 37550 24722
rect 37550 24670 37602 24722
rect 37602 24670 37604 24722
rect 37548 24668 37604 24670
rect 37772 24220 37828 24276
rect 36988 23042 37044 23044
rect 36988 22990 36990 23042
rect 36990 22990 37042 23042
rect 37042 22990 37044 23042
rect 36988 22988 37044 22990
rect 36876 22764 36932 22820
rect 36652 22258 36708 22260
rect 36652 22206 36654 22258
rect 36654 22206 36706 22258
rect 36706 22206 36708 22258
rect 36652 22204 36708 22206
rect 36988 22652 37044 22708
rect 36652 21810 36708 21812
rect 36652 21758 36654 21810
rect 36654 21758 36706 21810
rect 36706 21758 36708 21810
rect 36652 21756 36708 21758
rect 36652 21420 36708 21476
rect 36764 21308 36820 21364
rect 36652 20914 36708 20916
rect 36652 20862 36654 20914
rect 36654 20862 36706 20914
rect 36706 20862 36708 20914
rect 36652 20860 36708 20862
rect 35756 20300 35812 20356
rect 36204 20578 36260 20580
rect 36204 20526 36206 20578
rect 36206 20526 36258 20578
rect 36258 20526 36260 20578
rect 36204 20524 36260 20526
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35084 18956 35140 19012
rect 34748 18172 34804 18228
rect 34636 17836 34692 17892
rect 35532 18396 35588 18452
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 34524 16210 34580 16212
rect 34524 16158 34526 16210
rect 34526 16158 34578 16210
rect 34578 16158 34580 16210
rect 34524 16156 34580 16158
rect 34076 15986 34132 15988
rect 34076 15934 34078 15986
rect 34078 15934 34130 15986
rect 34130 15934 34132 15986
rect 34076 15932 34132 15934
rect 34300 15538 34356 15540
rect 34300 15486 34302 15538
rect 34302 15486 34354 15538
rect 34354 15486 34356 15538
rect 34300 15484 34356 15486
rect 34636 16044 34692 16100
rect 36092 19852 36148 19908
rect 35868 19122 35924 19124
rect 35868 19070 35870 19122
rect 35870 19070 35922 19122
rect 35922 19070 35924 19122
rect 35868 19068 35924 19070
rect 36092 18956 36148 19012
rect 36428 19458 36484 19460
rect 36428 19406 36430 19458
rect 36430 19406 36482 19458
rect 36482 19406 36484 19458
rect 36428 19404 36484 19406
rect 36204 18620 36260 18676
rect 36428 18956 36484 19012
rect 35980 18562 36036 18564
rect 35980 18510 35982 18562
rect 35982 18510 36034 18562
rect 36034 18510 36036 18562
rect 35980 18508 36036 18510
rect 36428 17778 36484 17780
rect 36428 17726 36430 17778
rect 36430 17726 36482 17778
rect 36482 17726 36484 17778
rect 36428 17724 36484 17726
rect 34860 15932 34916 15988
rect 35196 16940 35252 16996
rect 35420 17442 35476 17444
rect 35420 17390 35422 17442
rect 35422 17390 35474 17442
rect 35474 17390 35476 17442
rect 35420 17388 35476 17390
rect 36092 17276 36148 17332
rect 35532 17052 35588 17108
rect 35868 17052 35924 17108
rect 35644 16882 35700 16884
rect 35644 16830 35646 16882
rect 35646 16830 35698 16882
rect 35698 16830 35700 16882
rect 35644 16828 35700 16830
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 35308 16156 35364 16212
rect 35084 16098 35140 16100
rect 35084 16046 35086 16098
rect 35086 16046 35138 16098
rect 35138 16046 35140 16098
rect 35084 16044 35140 16046
rect 34972 15596 35028 15652
rect 34300 14306 34356 14308
rect 34300 14254 34302 14306
rect 34302 14254 34354 14306
rect 34354 14254 34356 14306
rect 34300 14252 34356 14254
rect 34412 13970 34468 13972
rect 34412 13918 34414 13970
rect 34414 13918 34466 13970
rect 34466 13918 34468 13970
rect 34412 13916 34468 13918
rect 33852 13468 33908 13524
rect 33628 12962 33684 12964
rect 33628 12910 33630 12962
rect 33630 12910 33682 12962
rect 33682 12910 33684 12962
rect 33628 12908 33684 12910
rect 33740 12796 33796 12852
rect 33964 12290 34020 12292
rect 33964 12238 33966 12290
rect 33966 12238 34018 12290
rect 34018 12238 34020 12290
rect 33964 12236 34020 12238
rect 34636 13020 34692 13076
rect 34524 12850 34580 12852
rect 34524 12798 34526 12850
rect 34526 12798 34578 12850
rect 34578 12798 34580 12850
rect 34524 12796 34580 12798
rect 35756 16098 35812 16100
rect 35756 16046 35758 16098
rect 35758 16046 35810 16098
rect 35810 16046 35812 16098
rect 35756 16044 35812 16046
rect 35084 15036 35140 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 36428 16940 36484 16996
rect 35980 16044 36036 16100
rect 36316 15986 36372 15988
rect 36316 15934 36318 15986
rect 36318 15934 36370 15986
rect 36370 15934 36372 15986
rect 36316 15932 36372 15934
rect 36652 20636 36708 20692
rect 36764 20524 36820 20580
rect 37100 21644 37156 21700
rect 37212 21420 37268 21476
rect 37884 23826 37940 23828
rect 37884 23774 37886 23826
rect 37886 23774 37938 23826
rect 37938 23774 37940 23826
rect 37884 23772 37940 23774
rect 37772 23436 37828 23492
rect 37436 22092 37492 22148
rect 37660 22316 37716 22372
rect 37548 21756 37604 21812
rect 37884 23324 37940 23380
rect 37884 22988 37940 23044
rect 38220 27132 38276 27188
rect 38444 27074 38500 27076
rect 38444 27022 38446 27074
rect 38446 27022 38498 27074
rect 38498 27022 38500 27074
rect 38444 27020 38500 27022
rect 38668 27356 38724 27412
rect 39676 32562 39732 32564
rect 39676 32510 39678 32562
rect 39678 32510 39730 32562
rect 39730 32510 39732 32562
rect 39676 32508 39732 32510
rect 38892 30268 38948 30324
rect 39004 29596 39060 29652
rect 39340 29708 39396 29764
rect 39340 28812 39396 28868
rect 39228 28754 39284 28756
rect 39228 28702 39230 28754
rect 39230 28702 39282 28754
rect 39282 28702 39284 28754
rect 39228 28700 39284 28702
rect 39116 27916 39172 27972
rect 39228 28028 39284 28084
rect 39788 31106 39844 31108
rect 39788 31054 39790 31106
rect 39790 31054 39842 31106
rect 39842 31054 39844 31106
rect 39788 31052 39844 31054
rect 40124 31724 40180 31780
rect 40236 33628 40292 33684
rect 39900 30604 39956 30660
rect 41580 38834 41636 38836
rect 41580 38782 41582 38834
rect 41582 38782 41634 38834
rect 41634 38782 41636 38834
rect 41580 38780 41636 38782
rect 41244 37212 41300 37268
rect 40460 33852 40516 33908
rect 40572 33516 40628 33572
rect 41020 33180 41076 33236
rect 40796 33068 40852 33124
rect 40908 32844 40964 32900
rect 40908 31554 40964 31556
rect 40908 31502 40910 31554
rect 40910 31502 40962 31554
rect 40962 31502 40964 31554
rect 40908 31500 40964 31502
rect 40908 31218 40964 31220
rect 40908 31166 40910 31218
rect 40910 31166 40962 31218
rect 40962 31166 40964 31218
rect 40908 31164 40964 31166
rect 40796 31106 40852 31108
rect 40796 31054 40798 31106
rect 40798 31054 40850 31106
rect 40850 31054 40852 31106
rect 40796 31052 40852 31054
rect 40460 30210 40516 30212
rect 40460 30158 40462 30210
rect 40462 30158 40514 30210
rect 40514 30158 40516 30210
rect 40460 30156 40516 30158
rect 40012 29820 40068 29876
rect 39564 28700 39620 28756
rect 39116 27468 39172 27524
rect 39116 27244 39172 27300
rect 39004 27132 39060 27188
rect 38332 26684 38388 26740
rect 38556 26850 38612 26852
rect 38556 26798 38558 26850
rect 38558 26798 38610 26850
rect 38610 26798 38612 26850
rect 38556 26796 38612 26798
rect 38332 26348 38388 26404
rect 38108 24668 38164 24724
rect 38668 26348 38724 26404
rect 38444 25900 38500 25956
rect 38332 25116 38388 25172
rect 38108 23660 38164 23716
rect 38220 24220 38276 24276
rect 38108 22652 38164 22708
rect 37884 22316 37940 22372
rect 37996 22092 38052 22148
rect 37772 21532 37828 21588
rect 37660 21026 37716 21028
rect 37660 20974 37662 21026
rect 37662 20974 37714 21026
rect 37714 20974 37716 21026
rect 37660 20972 37716 20974
rect 38108 21644 38164 21700
rect 37996 21532 38052 21588
rect 38108 21474 38164 21476
rect 38108 21422 38110 21474
rect 38110 21422 38162 21474
rect 38162 21422 38164 21474
rect 38108 21420 38164 21422
rect 37100 20300 37156 20356
rect 36652 18732 36708 18788
rect 36652 16380 36708 16436
rect 36540 16156 36596 16212
rect 36652 15986 36708 15988
rect 36652 15934 36654 15986
rect 36654 15934 36706 15986
rect 36706 15934 36708 15986
rect 36652 15932 36708 15934
rect 36092 15036 36148 15092
rect 36540 15314 36596 15316
rect 36540 15262 36542 15314
rect 36542 15262 36594 15314
rect 36594 15262 36596 15314
rect 36540 15260 36596 15262
rect 35308 13746 35364 13748
rect 35308 13694 35310 13746
rect 35310 13694 35362 13746
rect 35362 13694 35364 13746
rect 35308 13692 35364 13694
rect 36876 19852 36932 19908
rect 36876 18284 36932 18340
rect 37548 20018 37604 20020
rect 37548 19966 37550 20018
rect 37550 19966 37602 20018
rect 37602 19966 37604 20018
rect 37548 19964 37604 19966
rect 37212 19292 37268 19348
rect 37100 18956 37156 19012
rect 38332 23714 38388 23716
rect 38332 23662 38334 23714
rect 38334 23662 38386 23714
rect 38386 23662 38388 23714
rect 38332 23660 38388 23662
rect 38556 25564 38612 25620
rect 38892 26460 38948 26516
rect 38892 25228 38948 25284
rect 39228 27020 39284 27076
rect 39676 28642 39732 28644
rect 39676 28590 39678 28642
rect 39678 28590 39730 28642
rect 39730 28590 39732 28642
rect 39676 28588 39732 28590
rect 39788 27580 39844 27636
rect 40572 29820 40628 29876
rect 40124 28252 40180 28308
rect 39116 26236 39172 26292
rect 38780 24556 38836 24612
rect 38892 23938 38948 23940
rect 38892 23886 38894 23938
rect 38894 23886 38946 23938
rect 38946 23886 38948 23938
rect 38892 23884 38948 23886
rect 38444 23548 38500 23604
rect 38556 22876 38612 22932
rect 38556 22204 38612 22260
rect 38668 22428 38724 22484
rect 38220 21196 38276 21252
rect 38332 21980 38388 22036
rect 38556 21084 38612 21140
rect 38108 20802 38164 20804
rect 38108 20750 38110 20802
rect 38110 20750 38162 20802
rect 38162 20750 38164 20802
rect 38108 20748 38164 20750
rect 37884 19292 37940 19348
rect 37996 19906 38052 19908
rect 37996 19854 37998 19906
rect 37998 19854 38050 19906
rect 38050 19854 38052 19906
rect 37996 19852 38052 19854
rect 37548 18732 37604 18788
rect 37324 18562 37380 18564
rect 37324 18510 37326 18562
rect 37326 18510 37378 18562
rect 37378 18510 37380 18562
rect 37324 18508 37380 18510
rect 37548 18508 37604 18564
rect 36988 18060 37044 18116
rect 36876 17778 36932 17780
rect 36876 17726 36878 17778
rect 36878 17726 36930 17778
rect 36930 17726 36932 17778
rect 36876 17724 36932 17726
rect 36876 17164 36932 17220
rect 36988 17052 37044 17108
rect 37100 18172 37156 18228
rect 36988 16044 37044 16100
rect 37100 15708 37156 15764
rect 37100 15484 37156 15540
rect 36764 14700 36820 14756
rect 36316 14530 36372 14532
rect 36316 14478 36318 14530
rect 36318 14478 36370 14530
rect 36370 14478 36372 14530
rect 36316 14476 36372 14478
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 13074 35252 13076
rect 35196 13022 35198 13074
rect 35198 13022 35250 13074
rect 35250 13022 35252 13074
rect 35196 13020 35252 13022
rect 36540 14418 36596 14420
rect 36540 14366 36542 14418
rect 36542 14366 36594 14418
rect 36594 14366 36596 14418
rect 36540 14364 36596 14366
rect 36540 13746 36596 13748
rect 36540 13694 36542 13746
rect 36542 13694 36594 13746
rect 36594 13694 36596 13746
rect 36540 13692 36596 13694
rect 34860 12236 34916 12292
rect 34412 11452 34468 11508
rect 34076 11170 34132 11172
rect 34076 11118 34078 11170
rect 34078 11118 34130 11170
rect 34130 11118 34132 11170
rect 34076 11116 34132 11118
rect 34636 11170 34692 11172
rect 34636 11118 34638 11170
rect 34638 11118 34690 11170
rect 34690 11118 34692 11170
rect 34636 11116 34692 11118
rect 33964 9324 34020 9380
rect 34972 8988 35028 9044
rect 33628 7644 33684 7700
rect 35644 12348 35700 12404
rect 36092 12348 36148 12404
rect 36316 12290 36372 12292
rect 36316 12238 36318 12290
rect 36318 12238 36370 12290
rect 36370 12238 36372 12290
rect 36316 12236 36372 12238
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35756 11506 35812 11508
rect 35756 11454 35758 11506
rect 35758 11454 35810 11506
rect 35810 11454 35812 11506
rect 35756 11452 35812 11454
rect 35308 11170 35364 11172
rect 35308 11118 35310 11170
rect 35310 11118 35362 11170
rect 35362 11118 35364 11170
rect 35308 11116 35364 11118
rect 36204 11004 36260 11060
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 36092 9772 36148 9828
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35084 5964 35140 6020
rect 33516 5740 33572 5796
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 33852 5122 33908 5124
rect 33852 5070 33854 5122
rect 33854 5070 33906 5122
rect 33906 5070 33908 5122
rect 33852 5068 33908 5070
rect 34636 5122 34692 5124
rect 34636 5070 34638 5122
rect 34638 5070 34690 5122
rect 34690 5070 34692 5122
rect 34636 5068 34692 5070
rect 37212 15314 37268 15316
rect 37212 15262 37214 15314
rect 37214 15262 37266 15314
rect 37266 15262 37268 15314
rect 37212 15260 37268 15262
rect 36988 13916 37044 13972
rect 37100 14924 37156 14980
rect 36764 13132 36820 13188
rect 36876 12684 36932 12740
rect 36876 11788 36932 11844
rect 36652 9660 36708 9716
rect 36876 8930 36932 8932
rect 36876 8878 36878 8930
rect 36878 8878 36930 8930
rect 36930 8878 36932 8930
rect 36876 8876 36932 8878
rect 36316 6130 36372 6132
rect 36316 6078 36318 6130
rect 36318 6078 36370 6130
rect 36370 6078 36372 6130
rect 36316 6076 36372 6078
rect 36428 5234 36484 5236
rect 36428 5182 36430 5234
rect 36430 5182 36482 5234
rect 36482 5182 36484 5234
rect 36428 5180 36484 5182
rect 36876 5068 36932 5124
rect 36204 4284 36260 4340
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 32844 2716 32900 2772
rect 29148 1260 29204 1316
rect 37884 19122 37940 19124
rect 37884 19070 37886 19122
rect 37886 19070 37938 19122
rect 37938 19070 37940 19122
rect 37884 19068 37940 19070
rect 37772 19010 37828 19012
rect 37772 18958 37774 19010
rect 37774 18958 37826 19010
rect 37826 18958 37828 19010
rect 37772 18956 37828 18958
rect 37660 18172 37716 18228
rect 37436 17778 37492 17780
rect 37436 17726 37438 17778
rect 37438 17726 37490 17778
rect 37490 17726 37492 17778
rect 37436 17724 37492 17726
rect 37324 14588 37380 14644
rect 37436 17500 37492 17556
rect 37212 13634 37268 13636
rect 37212 13582 37214 13634
rect 37214 13582 37266 13634
rect 37266 13582 37268 13634
rect 37212 13580 37268 13582
rect 37324 13132 37380 13188
rect 37548 17106 37604 17108
rect 37548 17054 37550 17106
rect 37550 17054 37602 17106
rect 37602 17054 37604 17106
rect 37548 17052 37604 17054
rect 38332 20636 38388 20692
rect 38444 20524 38500 20580
rect 37996 18284 38052 18340
rect 38108 18172 38164 18228
rect 37996 16882 38052 16884
rect 37996 16830 37998 16882
rect 37998 16830 38050 16882
rect 38050 16830 38052 16882
rect 37996 16828 38052 16830
rect 38332 17442 38388 17444
rect 38332 17390 38334 17442
rect 38334 17390 38386 17442
rect 38386 17390 38388 17442
rect 38332 17388 38388 17390
rect 37884 16156 37940 16212
rect 37996 16268 38052 16324
rect 38108 16098 38164 16100
rect 38108 16046 38110 16098
rect 38110 16046 38162 16098
rect 38162 16046 38164 16098
rect 38108 16044 38164 16046
rect 37660 15986 37716 15988
rect 37660 15934 37662 15986
rect 37662 15934 37714 15986
rect 37714 15934 37716 15986
rect 37660 15932 37716 15934
rect 37884 15932 37940 15988
rect 37548 15820 37604 15876
rect 37772 15484 37828 15540
rect 38108 15538 38164 15540
rect 38108 15486 38110 15538
rect 38110 15486 38162 15538
rect 38162 15486 38164 15538
rect 38108 15484 38164 15486
rect 37996 15314 38052 15316
rect 37996 15262 37998 15314
rect 37998 15262 38050 15314
rect 38050 15262 38052 15314
rect 37996 15260 38052 15262
rect 37884 14418 37940 14420
rect 37884 14366 37886 14418
rect 37886 14366 37938 14418
rect 37938 14366 37940 14418
rect 37884 14364 37940 14366
rect 37660 13970 37716 13972
rect 37660 13918 37662 13970
rect 37662 13918 37714 13970
rect 37714 13918 37716 13970
rect 37660 13916 37716 13918
rect 38444 16492 38500 16548
rect 38332 15484 38388 15540
rect 38444 15820 38500 15876
rect 39228 26012 39284 26068
rect 39564 25900 39620 25956
rect 39564 25506 39620 25508
rect 39564 25454 39566 25506
rect 39566 25454 39618 25506
rect 39618 25454 39620 25506
rect 39564 25452 39620 25454
rect 39452 25116 39508 25172
rect 40348 28252 40404 28308
rect 40012 26124 40068 26180
rect 40796 30156 40852 30212
rect 40796 29932 40852 29988
rect 40684 29708 40740 29764
rect 40796 29148 40852 29204
rect 40572 29036 40628 29092
rect 40796 28924 40852 28980
rect 40572 28140 40628 28196
rect 40572 27970 40628 27972
rect 40572 27918 40574 27970
rect 40574 27918 40626 27970
rect 40626 27918 40628 27970
rect 40572 27916 40628 27918
rect 40348 27132 40404 27188
rect 40908 27692 40964 27748
rect 40460 26908 40516 26964
rect 39340 25004 39396 25060
rect 40236 26796 40292 26852
rect 39340 23996 39396 24052
rect 39900 25228 39956 25284
rect 39340 23826 39396 23828
rect 39340 23774 39342 23826
rect 39342 23774 39394 23826
rect 39394 23774 39396 23826
rect 39340 23772 39396 23774
rect 39004 22988 39060 23044
rect 39228 23660 39284 23716
rect 39004 21474 39060 21476
rect 39004 21422 39006 21474
rect 39006 21422 39058 21474
rect 39058 21422 39060 21474
rect 39004 21420 39060 21422
rect 38892 21196 38948 21252
rect 39116 20188 39172 20244
rect 38780 18674 38836 18676
rect 38780 18622 38782 18674
rect 38782 18622 38834 18674
rect 38834 18622 38836 18674
rect 38780 18620 38836 18622
rect 39452 22146 39508 22148
rect 39452 22094 39454 22146
rect 39454 22094 39506 22146
rect 39506 22094 39508 22146
rect 39452 22092 39508 22094
rect 39340 21420 39396 21476
rect 39452 21308 39508 21364
rect 39116 18956 39172 19012
rect 39228 19068 39284 19124
rect 39564 20860 39620 20916
rect 40348 26572 40404 26628
rect 40684 26796 40740 26852
rect 41244 34748 41300 34804
rect 41244 34188 41300 34244
rect 41244 33180 41300 33236
rect 41244 30098 41300 30100
rect 41244 30046 41246 30098
rect 41246 30046 41298 30098
rect 41298 30046 41300 30098
rect 41244 30044 41300 30046
rect 41468 37938 41524 37940
rect 41468 37886 41470 37938
rect 41470 37886 41522 37938
rect 41522 37886 41524 37938
rect 41468 37884 41524 37886
rect 41692 37378 41748 37380
rect 41692 37326 41694 37378
rect 41694 37326 41746 37378
rect 41746 37326 41748 37378
rect 41692 37324 41748 37326
rect 42028 38946 42084 38948
rect 42028 38894 42030 38946
rect 42030 38894 42082 38946
rect 42082 38894 42084 38946
rect 42028 38892 42084 38894
rect 42476 38834 42532 38836
rect 42476 38782 42478 38834
rect 42478 38782 42530 38834
rect 42530 38782 42532 38834
rect 42476 38780 42532 38782
rect 41916 38722 41972 38724
rect 41916 38670 41918 38722
rect 41918 38670 41970 38722
rect 41970 38670 41972 38722
rect 41916 38668 41972 38670
rect 42028 38444 42084 38500
rect 41916 37266 41972 37268
rect 41916 37214 41918 37266
rect 41918 37214 41970 37266
rect 41970 37214 41972 37266
rect 41916 37212 41972 37214
rect 42812 40012 42868 40068
rect 43708 47740 43764 47796
rect 43484 45890 43540 45892
rect 43484 45838 43486 45890
rect 43486 45838 43538 45890
rect 43538 45838 43540 45890
rect 43484 45836 43540 45838
rect 43708 46620 43764 46676
rect 44156 47628 44212 47684
rect 44044 47458 44100 47460
rect 44044 47406 44046 47458
rect 44046 47406 44098 47458
rect 44098 47406 44100 47458
rect 44044 47404 44100 47406
rect 44604 49698 44660 49700
rect 44604 49646 44606 49698
rect 44606 49646 44658 49698
rect 44658 49646 44660 49698
rect 44604 49644 44660 49646
rect 44604 47964 44660 48020
rect 46284 51548 46340 51604
rect 46508 52050 46564 52052
rect 46508 51998 46510 52050
rect 46510 51998 46562 52050
rect 46562 51998 46564 52050
rect 46508 51996 46564 51998
rect 47068 52274 47124 52276
rect 47068 52222 47070 52274
rect 47070 52222 47122 52274
rect 47122 52222 47124 52274
rect 47068 52220 47124 52222
rect 47180 51884 47236 51940
rect 47516 52050 47572 52052
rect 47516 51998 47518 52050
rect 47518 51998 47570 52050
rect 47570 51998 47572 52050
rect 47516 51996 47572 51998
rect 46844 51548 46900 51604
rect 46396 51436 46452 51492
rect 47292 51436 47348 51492
rect 45052 50988 45108 51044
rect 45388 50594 45444 50596
rect 45388 50542 45390 50594
rect 45390 50542 45442 50594
rect 45442 50542 45444 50594
rect 45388 50540 45444 50542
rect 45724 50482 45780 50484
rect 45724 50430 45726 50482
rect 45726 50430 45778 50482
rect 45778 50430 45780 50482
rect 45724 50428 45780 50430
rect 45612 49980 45668 50036
rect 45052 49644 45108 49700
rect 44828 47852 44884 47908
rect 44604 47068 44660 47124
rect 44268 46898 44324 46900
rect 44268 46846 44270 46898
rect 44270 46846 44322 46898
rect 44322 46846 44324 46898
rect 44268 46844 44324 46846
rect 44492 46844 44548 46900
rect 44044 46674 44100 46676
rect 44044 46622 44046 46674
rect 44046 46622 44098 46674
rect 44098 46622 44100 46674
rect 44044 46620 44100 46622
rect 45052 46786 45108 46788
rect 45052 46734 45054 46786
rect 45054 46734 45106 46786
rect 45106 46734 45108 46786
rect 45052 46732 45108 46734
rect 44716 46620 44772 46676
rect 44492 45836 44548 45892
rect 43820 45276 43876 45332
rect 43372 43148 43428 43204
rect 43932 44434 43988 44436
rect 43932 44382 43934 44434
rect 43934 44382 43986 44434
rect 43986 44382 43988 44434
rect 43932 44380 43988 44382
rect 43820 43484 43876 43540
rect 43708 43036 43764 43092
rect 43820 42924 43876 42980
rect 44044 43820 44100 43876
rect 44156 45276 44212 45332
rect 43708 42476 43764 42532
rect 43820 41804 43876 41860
rect 43596 41356 43652 41412
rect 44044 41244 44100 41300
rect 43260 41020 43316 41076
rect 43596 40796 43652 40852
rect 42812 39452 42868 39508
rect 42588 38668 42644 38724
rect 42476 37212 42532 37268
rect 42812 37266 42868 37268
rect 42812 37214 42814 37266
rect 42814 37214 42866 37266
rect 42866 37214 42868 37266
rect 42812 37212 42868 37214
rect 42028 37100 42084 37156
rect 41580 36540 41636 36596
rect 41468 35586 41524 35588
rect 41468 35534 41470 35586
rect 41470 35534 41522 35586
rect 41522 35534 41524 35586
rect 41468 35532 41524 35534
rect 41468 35308 41524 35364
rect 42476 36258 42532 36260
rect 42476 36206 42478 36258
rect 42478 36206 42530 36258
rect 42530 36206 42532 36258
rect 42476 36204 42532 36206
rect 43148 40460 43204 40516
rect 43260 39730 43316 39732
rect 43260 39678 43262 39730
rect 43262 39678 43314 39730
rect 43314 39678 43316 39730
rect 43260 39676 43316 39678
rect 43260 39452 43316 39508
rect 43148 39004 43204 39060
rect 43372 38162 43428 38164
rect 43372 38110 43374 38162
rect 43374 38110 43426 38162
rect 43426 38110 43428 38162
rect 43372 38108 43428 38110
rect 43148 37548 43204 37604
rect 43036 37324 43092 37380
rect 43260 37154 43316 37156
rect 43260 37102 43262 37154
rect 43262 37102 43314 37154
rect 43314 37102 43316 37154
rect 43260 37100 43316 37102
rect 43372 36988 43428 37044
rect 41916 35196 41972 35252
rect 41580 34748 41636 34804
rect 42252 34636 42308 34692
rect 42028 33628 42084 33684
rect 41580 33346 41636 33348
rect 41580 33294 41582 33346
rect 41582 33294 41634 33346
rect 41634 33294 41636 33346
rect 41580 33292 41636 33294
rect 42028 33292 42084 33348
rect 41692 32844 41748 32900
rect 41468 32396 41524 32452
rect 41580 32060 41636 32116
rect 41468 31778 41524 31780
rect 41468 31726 41470 31778
rect 41470 31726 41522 31778
rect 41522 31726 41524 31778
rect 41468 31724 41524 31726
rect 41468 30604 41524 30660
rect 41916 33234 41972 33236
rect 41916 33182 41918 33234
rect 41918 33182 41970 33234
rect 41970 33182 41972 33234
rect 41916 33180 41972 33182
rect 41916 31948 41972 32004
rect 41692 29596 41748 29652
rect 42252 32508 42308 32564
rect 41580 29538 41636 29540
rect 41580 29486 41582 29538
rect 41582 29486 41634 29538
rect 41634 29486 41636 29538
rect 41580 29484 41636 29486
rect 41468 29148 41524 29204
rect 41356 28924 41412 28980
rect 42028 31276 42084 31332
rect 42140 30770 42196 30772
rect 42140 30718 42142 30770
rect 42142 30718 42194 30770
rect 42194 30718 42196 30770
rect 42140 30716 42196 30718
rect 41916 29426 41972 29428
rect 41916 29374 41918 29426
rect 41918 29374 41970 29426
rect 41970 29374 41972 29426
rect 41916 29372 41972 29374
rect 41804 28588 41860 28644
rect 41580 28476 41636 28532
rect 41244 27692 41300 27748
rect 41132 27580 41188 27636
rect 41132 26908 41188 26964
rect 40572 26236 40628 26292
rect 40796 26178 40852 26180
rect 40796 26126 40798 26178
rect 40798 26126 40850 26178
rect 40850 26126 40852 26178
rect 40796 26124 40852 26126
rect 40684 25564 40740 25620
rect 40236 25116 40292 25172
rect 39788 23548 39844 23604
rect 39900 23324 39956 23380
rect 40460 25282 40516 25284
rect 40460 25230 40462 25282
rect 40462 25230 40514 25282
rect 40514 25230 40516 25282
rect 40460 25228 40516 25230
rect 40348 24444 40404 24500
rect 40236 24050 40292 24052
rect 40236 23998 40238 24050
rect 40238 23998 40290 24050
rect 40290 23998 40292 24050
rect 40236 23996 40292 23998
rect 40348 23266 40404 23268
rect 40348 23214 40350 23266
rect 40350 23214 40402 23266
rect 40402 23214 40404 23266
rect 40348 23212 40404 23214
rect 40236 22428 40292 22484
rect 40012 22370 40068 22372
rect 40012 22318 40014 22370
rect 40014 22318 40066 22370
rect 40066 22318 40068 22370
rect 40012 22316 40068 22318
rect 40348 22316 40404 22372
rect 40236 22146 40292 22148
rect 40236 22094 40238 22146
rect 40238 22094 40290 22146
rect 40290 22094 40292 22146
rect 40236 22092 40292 22094
rect 40460 22258 40516 22260
rect 40460 22206 40462 22258
rect 40462 22206 40514 22258
rect 40514 22206 40516 22258
rect 40460 22204 40516 22206
rect 40684 24050 40740 24052
rect 40684 23998 40686 24050
rect 40686 23998 40738 24050
rect 40738 23998 40740 24050
rect 40684 23996 40740 23998
rect 41020 25228 41076 25284
rect 40684 22988 40740 23044
rect 41020 24332 41076 24388
rect 40572 21868 40628 21924
rect 40012 20972 40068 21028
rect 40124 21532 40180 21588
rect 39900 20690 39956 20692
rect 39900 20638 39902 20690
rect 39902 20638 39954 20690
rect 39954 20638 39956 20690
rect 39900 20636 39956 20638
rect 39452 19068 39508 19124
rect 39116 18562 39172 18564
rect 39116 18510 39118 18562
rect 39118 18510 39170 18562
rect 39170 18510 39172 18562
rect 39116 18508 39172 18510
rect 39116 16268 39172 16324
rect 40124 20242 40180 20244
rect 40124 20190 40126 20242
rect 40126 20190 40178 20242
rect 40178 20190 40180 20242
rect 40124 20188 40180 20190
rect 40012 19234 40068 19236
rect 40012 19182 40014 19234
rect 40014 19182 40066 19234
rect 40066 19182 40068 19234
rect 40012 19180 40068 19182
rect 39676 19122 39732 19124
rect 39676 19070 39678 19122
rect 39678 19070 39730 19122
rect 39730 19070 39732 19122
rect 39676 19068 39732 19070
rect 39900 18956 39956 19012
rect 39676 18844 39732 18900
rect 39228 16156 39284 16212
rect 40348 21586 40404 21588
rect 40348 21534 40350 21586
rect 40350 21534 40402 21586
rect 40402 21534 40404 21586
rect 40348 21532 40404 21534
rect 40572 21420 40628 21476
rect 40908 23378 40964 23380
rect 40908 23326 40910 23378
rect 40910 23326 40962 23378
rect 40962 23326 40964 23378
rect 40908 23324 40964 23326
rect 41580 28082 41636 28084
rect 41580 28030 41582 28082
rect 41582 28030 41634 28082
rect 41634 28030 41636 28082
rect 41580 28028 41636 28030
rect 41468 27468 41524 27524
rect 41916 27356 41972 27412
rect 41804 27132 41860 27188
rect 41580 26572 41636 26628
rect 41356 26124 41412 26180
rect 41468 26460 41524 26516
rect 41580 24946 41636 24948
rect 41580 24894 41582 24946
rect 41582 24894 41634 24946
rect 41634 24894 41636 24946
rect 41580 24892 41636 24894
rect 42140 30098 42196 30100
rect 42140 30046 42142 30098
rect 42142 30046 42194 30098
rect 42194 30046 42196 30098
rect 42140 30044 42196 30046
rect 42588 32844 42644 32900
rect 42588 32172 42644 32228
rect 42700 31948 42756 32004
rect 42700 31612 42756 31668
rect 43260 36204 43316 36260
rect 42924 35308 42980 35364
rect 43036 34300 43092 34356
rect 43260 33964 43316 34020
rect 43372 35756 43428 35812
rect 43260 33122 43316 33124
rect 43260 33070 43262 33122
rect 43262 33070 43314 33122
rect 43314 33070 43316 33122
rect 43260 33068 43316 33070
rect 42924 32844 42980 32900
rect 43036 32562 43092 32564
rect 43036 32510 43038 32562
rect 43038 32510 43090 32562
rect 43090 32510 43092 32562
rect 43036 32508 43092 32510
rect 45388 48914 45444 48916
rect 45388 48862 45390 48914
rect 45390 48862 45442 48914
rect 45442 48862 45444 48914
rect 45388 48860 45444 48862
rect 45836 49420 45892 49476
rect 45500 48636 45556 48692
rect 47740 52050 47796 52052
rect 47740 51998 47742 52050
rect 47742 51998 47794 52050
rect 47794 51998 47796 52050
rect 47740 51996 47796 51998
rect 47628 51548 47684 51604
rect 47740 51772 47796 51828
rect 47180 50428 47236 50484
rect 46060 48636 46116 48692
rect 46508 49980 46564 50036
rect 45500 47852 45556 47908
rect 45500 47628 45556 47684
rect 45388 46844 45444 46900
rect 45164 46620 45220 46676
rect 44716 45836 44772 45892
rect 46060 47516 46116 47572
rect 45948 46844 46004 46900
rect 45612 46396 45668 46452
rect 45724 45778 45780 45780
rect 45724 45726 45726 45778
rect 45726 45726 45778 45778
rect 45778 45726 45780 45778
rect 45724 45724 45780 45726
rect 45836 45612 45892 45668
rect 44380 43596 44436 43652
rect 44268 42754 44324 42756
rect 44268 42702 44270 42754
rect 44270 42702 44322 42754
rect 44322 42702 44324 42754
rect 44268 42700 44324 42702
rect 46396 49138 46452 49140
rect 46396 49086 46398 49138
rect 46398 49086 46450 49138
rect 46450 49086 46452 49138
rect 46396 49084 46452 49086
rect 46844 49980 46900 50036
rect 46844 49644 46900 49700
rect 46732 49026 46788 49028
rect 46732 48974 46734 49026
rect 46734 48974 46786 49026
rect 46786 48974 46788 49026
rect 46732 48972 46788 48974
rect 46956 49138 47012 49140
rect 46956 49086 46958 49138
rect 46958 49086 47010 49138
rect 47010 49086 47012 49138
rect 46956 49084 47012 49086
rect 46844 48860 46900 48916
rect 46284 48748 46340 48804
rect 47180 48466 47236 48468
rect 47180 48414 47182 48466
rect 47182 48414 47234 48466
rect 47234 48414 47236 48466
rect 47180 48412 47236 48414
rect 46172 46508 46228 46564
rect 45948 45500 46004 45556
rect 46060 45164 46116 45220
rect 46396 45052 46452 45108
rect 47180 47964 47236 48020
rect 52332 55468 52388 55524
rect 50556 54906 50612 54908
rect 50556 54854 50558 54906
rect 50558 54854 50610 54906
rect 50610 54854 50612 54906
rect 50556 54852 50612 54854
rect 50660 54906 50716 54908
rect 50660 54854 50662 54906
rect 50662 54854 50714 54906
rect 50714 54854 50716 54906
rect 50660 54852 50716 54854
rect 50764 54906 50820 54908
rect 50764 54854 50766 54906
rect 50766 54854 50818 54906
rect 50818 54854 50820 54906
rect 50764 54852 50820 54854
rect 50556 53338 50612 53340
rect 50556 53286 50558 53338
rect 50558 53286 50610 53338
rect 50610 53286 50612 53338
rect 50556 53284 50612 53286
rect 50660 53338 50716 53340
rect 50660 53286 50662 53338
rect 50662 53286 50714 53338
rect 50714 53286 50716 53338
rect 50660 53284 50716 53286
rect 50764 53338 50820 53340
rect 50764 53286 50766 53338
rect 50766 53286 50818 53338
rect 50818 53286 50820 53338
rect 50764 53284 50820 53286
rect 49308 52274 49364 52276
rect 49308 52222 49310 52274
rect 49310 52222 49362 52274
rect 49362 52222 49364 52274
rect 49308 52220 49364 52222
rect 50876 52220 50932 52276
rect 48412 51772 48468 51828
rect 47852 51660 47908 51716
rect 48412 51436 48468 51492
rect 48076 50428 48132 50484
rect 47516 50034 47572 50036
rect 47516 49982 47518 50034
rect 47518 49982 47570 50034
rect 47570 49982 47572 50034
rect 47516 49980 47572 49982
rect 47516 49756 47572 49812
rect 47404 49698 47460 49700
rect 47404 49646 47406 49698
rect 47406 49646 47458 49698
rect 47458 49646 47460 49698
rect 47404 49644 47460 49646
rect 47516 48860 47572 48916
rect 47404 48524 47460 48580
rect 47292 46674 47348 46676
rect 47292 46622 47294 46674
rect 47294 46622 47346 46674
rect 47346 46622 47348 46674
rect 47292 46620 47348 46622
rect 47852 49756 47908 49812
rect 47740 49138 47796 49140
rect 47740 49086 47742 49138
rect 47742 49086 47794 49138
rect 47794 49086 47796 49138
rect 47740 49084 47796 49086
rect 47852 49026 47908 49028
rect 47852 48974 47854 49026
rect 47854 48974 47906 49026
rect 47906 48974 47908 49026
rect 47852 48972 47908 48974
rect 47628 48636 47684 48692
rect 47516 46620 47572 46676
rect 47404 46172 47460 46228
rect 46956 45724 47012 45780
rect 46620 44156 46676 44212
rect 44716 43650 44772 43652
rect 44716 43598 44718 43650
rect 44718 43598 44770 43650
rect 44770 43598 44772 43650
rect 44716 43596 44772 43598
rect 44940 43426 44996 43428
rect 44940 43374 44942 43426
rect 44942 43374 44994 43426
rect 44994 43374 44996 43426
rect 44940 43372 44996 43374
rect 44492 42476 44548 42532
rect 44828 42082 44884 42084
rect 44828 42030 44830 42082
rect 44830 42030 44882 42082
rect 44882 42030 44884 42082
rect 44828 42028 44884 42030
rect 44492 41804 44548 41860
rect 44380 41132 44436 41188
rect 44940 40796 44996 40852
rect 43820 39452 43876 39508
rect 44044 39506 44100 39508
rect 44044 39454 44046 39506
rect 44046 39454 44098 39506
rect 44098 39454 44100 39506
rect 44044 39452 44100 39454
rect 44044 37938 44100 37940
rect 44044 37886 44046 37938
rect 44046 37886 44098 37938
rect 44098 37886 44100 37938
rect 44044 37884 44100 37886
rect 44156 37772 44212 37828
rect 44044 37548 44100 37604
rect 43932 37266 43988 37268
rect 43932 37214 43934 37266
rect 43934 37214 43986 37266
rect 43986 37214 43988 37266
rect 43932 37212 43988 37214
rect 43708 35810 43764 35812
rect 43708 35758 43710 35810
rect 43710 35758 43762 35810
rect 43762 35758 43764 35810
rect 43708 35756 43764 35758
rect 43372 32060 43428 32116
rect 43484 34300 43540 34356
rect 43148 31836 43204 31892
rect 43036 31724 43092 31780
rect 42588 30882 42644 30884
rect 42588 30830 42590 30882
rect 42590 30830 42642 30882
rect 42642 30830 42644 30882
rect 42588 30828 42644 30830
rect 43596 34076 43652 34132
rect 43708 35532 43764 35588
rect 43932 34690 43988 34692
rect 43932 34638 43934 34690
rect 43934 34638 43986 34690
rect 43986 34638 43988 34690
rect 43932 34636 43988 34638
rect 43820 33628 43876 33684
rect 43708 33122 43764 33124
rect 43708 33070 43710 33122
rect 43710 33070 43762 33122
rect 43762 33070 43764 33122
rect 43708 33068 43764 33070
rect 44716 40684 44772 40740
rect 44604 40626 44660 40628
rect 44604 40574 44606 40626
rect 44606 40574 44658 40626
rect 44658 40574 44660 40626
rect 44604 40572 44660 40574
rect 44492 40514 44548 40516
rect 44492 40462 44494 40514
rect 44494 40462 44546 40514
rect 44546 40462 44548 40514
rect 44492 40460 44548 40462
rect 44380 39452 44436 39508
rect 44156 37100 44212 37156
rect 44156 36370 44212 36372
rect 44156 36318 44158 36370
rect 44158 36318 44210 36370
rect 44210 36318 44212 36370
rect 44156 36316 44212 36318
rect 44268 36988 44324 37044
rect 44492 39004 44548 39060
rect 44716 38108 44772 38164
rect 44492 37826 44548 37828
rect 44492 37774 44494 37826
rect 44494 37774 44546 37826
rect 44546 37774 44548 37826
rect 44492 37772 44548 37774
rect 44604 36988 44660 37044
rect 44492 36428 44548 36484
rect 44604 36316 44660 36372
rect 44380 35980 44436 36036
rect 44604 35810 44660 35812
rect 44604 35758 44606 35810
rect 44606 35758 44658 35810
rect 44658 35758 44660 35810
rect 44604 35756 44660 35758
rect 44492 35532 44548 35588
rect 46620 43820 46676 43876
rect 46172 43596 46228 43652
rect 45276 43538 45332 43540
rect 45276 43486 45278 43538
rect 45278 43486 45330 43538
rect 45330 43486 45332 43538
rect 45276 43484 45332 43486
rect 45836 43538 45892 43540
rect 45836 43486 45838 43538
rect 45838 43486 45890 43538
rect 45890 43486 45892 43538
rect 45836 43484 45892 43486
rect 45724 42978 45780 42980
rect 45724 42926 45726 42978
rect 45726 42926 45778 42978
rect 45778 42926 45780 42978
rect 45724 42924 45780 42926
rect 45164 42252 45220 42308
rect 45388 42364 45444 42420
rect 45276 42194 45332 42196
rect 45276 42142 45278 42194
rect 45278 42142 45330 42194
rect 45330 42142 45332 42194
rect 45276 42140 45332 42142
rect 45164 41804 45220 41860
rect 45388 41580 45444 41636
rect 45612 41356 45668 41412
rect 45388 41074 45444 41076
rect 45388 41022 45390 41074
rect 45390 41022 45442 41074
rect 45442 41022 45444 41074
rect 45388 41020 45444 41022
rect 45276 39340 45332 39396
rect 45500 39394 45556 39396
rect 45500 39342 45502 39394
rect 45502 39342 45554 39394
rect 45554 39342 45556 39394
rect 45500 39340 45556 39342
rect 45724 38892 45780 38948
rect 45612 38444 45668 38500
rect 45500 37938 45556 37940
rect 45500 37886 45502 37938
rect 45502 37886 45554 37938
rect 45554 37886 45556 37938
rect 45500 37884 45556 37886
rect 46620 43538 46676 43540
rect 46620 43486 46622 43538
rect 46622 43486 46674 43538
rect 46674 43486 46676 43538
rect 46620 43484 46676 43486
rect 45948 42754 46004 42756
rect 45948 42702 45950 42754
rect 45950 42702 46002 42754
rect 46002 42702 46004 42754
rect 45948 42700 46004 42702
rect 46060 42642 46116 42644
rect 46060 42590 46062 42642
rect 46062 42590 46114 42642
rect 46114 42590 46116 42642
rect 46060 42588 46116 42590
rect 45948 41970 46004 41972
rect 45948 41918 45950 41970
rect 45950 41918 46002 41970
rect 46002 41918 46004 41970
rect 45948 41916 46004 41918
rect 46732 42924 46788 42980
rect 46844 43596 46900 43652
rect 46844 42700 46900 42756
rect 46060 40684 46116 40740
rect 46396 40962 46452 40964
rect 46396 40910 46398 40962
rect 46398 40910 46450 40962
rect 46450 40910 46452 40962
rect 46396 40908 46452 40910
rect 46284 40684 46340 40740
rect 46844 41074 46900 41076
rect 46844 41022 46846 41074
rect 46846 41022 46898 41074
rect 46898 41022 46900 41074
rect 46844 41020 46900 41022
rect 46732 40908 46788 40964
rect 46620 40460 46676 40516
rect 46396 40348 46452 40404
rect 46844 40684 46900 40740
rect 47180 44322 47236 44324
rect 47180 44270 47182 44322
rect 47182 44270 47234 44322
rect 47234 44270 47236 44322
rect 47180 44268 47236 44270
rect 47404 43820 47460 43876
rect 47516 44156 47572 44212
rect 47068 41244 47124 41300
rect 47852 48242 47908 48244
rect 47852 48190 47854 48242
rect 47854 48190 47906 48242
rect 47906 48190 47908 48242
rect 47852 48188 47908 48190
rect 48188 49250 48244 49252
rect 48188 49198 48190 49250
rect 48190 49198 48242 49250
rect 48242 49198 48244 49250
rect 48188 49196 48244 49198
rect 48076 48748 48132 48804
rect 48188 48242 48244 48244
rect 48188 48190 48190 48242
rect 48190 48190 48242 48242
rect 48242 48190 48244 48242
rect 48188 48188 48244 48190
rect 47852 47852 47908 47908
rect 49196 51996 49252 52052
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 49868 51602 49924 51604
rect 49868 51550 49870 51602
rect 49870 51550 49922 51602
rect 49922 51550 49924 51602
rect 49868 51548 49924 51550
rect 48524 49644 48580 49700
rect 48636 49308 48692 49364
rect 48636 48914 48692 48916
rect 48636 48862 48638 48914
rect 48638 48862 48690 48914
rect 48690 48862 48692 48914
rect 48636 48860 48692 48862
rect 47852 45612 47908 45668
rect 48412 46674 48468 46676
rect 48412 46622 48414 46674
rect 48414 46622 48466 46674
rect 48466 46622 48468 46674
rect 48412 46620 48468 46622
rect 48412 45890 48468 45892
rect 48412 45838 48414 45890
rect 48414 45838 48466 45890
rect 48466 45838 48468 45890
rect 48412 45836 48468 45838
rect 48076 45724 48132 45780
rect 48860 48748 48916 48804
rect 49532 50876 49588 50932
rect 49420 49980 49476 50036
rect 50204 50876 50260 50932
rect 49756 49980 49812 50036
rect 48972 48412 49028 48468
rect 49308 46508 49364 46564
rect 48972 46284 49028 46340
rect 48076 45218 48132 45220
rect 48076 45166 48078 45218
rect 48078 45166 48130 45218
rect 48130 45166 48132 45218
rect 48076 45164 48132 45166
rect 47964 45106 48020 45108
rect 47964 45054 47966 45106
rect 47966 45054 48018 45106
rect 48018 45054 48020 45106
rect 47964 45052 48020 45054
rect 48748 45164 48804 45220
rect 48972 45836 49028 45892
rect 49084 45052 49140 45108
rect 48412 44210 48468 44212
rect 48412 44158 48414 44210
rect 48414 44158 48466 44210
rect 48466 44158 48468 44210
rect 48412 44156 48468 44158
rect 47516 42530 47572 42532
rect 47516 42478 47518 42530
rect 47518 42478 47570 42530
rect 47570 42478 47572 42530
rect 47516 42476 47572 42478
rect 47404 40908 47460 40964
rect 48860 44322 48916 44324
rect 48860 44270 48862 44322
rect 48862 44270 48914 44322
rect 48914 44270 48916 44322
rect 48860 44268 48916 44270
rect 48636 43708 48692 43764
rect 48076 43650 48132 43652
rect 48076 43598 48078 43650
rect 48078 43598 48130 43650
rect 48130 43598 48132 43650
rect 48076 43596 48132 43598
rect 48412 43596 48468 43652
rect 48188 43372 48244 43428
rect 47740 41244 47796 41300
rect 47852 42028 47908 42084
rect 47516 40796 47572 40852
rect 47404 40402 47460 40404
rect 47404 40350 47406 40402
rect 47406 40350 47458 40402
rect 47458 40350 47460 40402
rect 47404 40348 47460 40350
rect 46620 39340 46676 39396
rect 46508 38946 46564 38948
rect 46508 38894 46510 38946
rect 46510 38894 46562 38946
rect 46562 38894 46564 38946
rect 46508 38892 46564 38894
rect 47292 38892 47348 38948
rect 47068 38444 47124 38500
rect 45724 37884 45780 37940
rect 45612 37660 45668 37716
rect 45276 37212 45332 37268
rect 46060 37436 46116 37492
rect 45052 36652 45108 36708
rect 45276 36428 45332 36484
rect 45164 36204 45220 36260
rect 45164 35756 45220 35812
rect 44380 34802 44436 34804
rect 44380 34750 44382 34802
rect 44382 34750 44434 34802
rect 44434 34750 44436 34802
rect 44380 34748 44436 34750
rect 44268 33852 44324 33908
rect 44156 33346 44212 33348
rect 44156 33294 44158 33346
rect 44158 33294 44210 33346
rect 44210 33294 44212 33346
rect 44156 33292 44212 33294
rect 43484 31724 43540 31780
rect 43148 31052 43204 31108
rect 43260 31500 43316 31556
rect 43036 30940 43092 30996
rect 42476 30268 42532 30324
rect 42588 29932 42644 29988
rect 42364 29484 42420 29540
rect 43148 30828 43204 30884
rect 42812 29484 42868 29540
rect 42700 29148 42756 29204
rect 42252 28028 42308 28084
rect 42364 29036 42420 29092
rect 42252 27692 42308 27748
rect 42140 27020 42196 27076
rect 42812 29036 42868 29092
rect 42924 30604 42980 30660
rect 43036 29820 43092 29876
rect 41804 26348 41860 26404
rect 42140 26684 42196 26740
rect 42028 26012 42084 26068
rect 41916 24444 41972 24500
rect 41804 24332 41860 24388
rect 41468 23772 41524 23828
rect 40908 22316 40964 22372
rect 41132 22204 41188 22260
rect 42140 25788 42196 25844
rect 42364 26572 42420 26628
rect 42364 26012 42420 26068
rect 42364 25228 42420 25284
rect 42364 24332 42420 24388
rect 41692 24050 41748 24052
rect 41692 23998 41694 24050
rect 41694 23998 41746 24050
rect 41746 23998 41748 24050
rect 41692 23996 41748 23998
rect 42140 24108 42196 24164
rect 41580 23100 41636 23156
rect 40348 20578 40404 20580
rect 40348 20526 40350 20578
rect 40350 20526 40402 20578
rect 40402 20526 40404 20578
rect 40348 20524 40404 20526
rect 40348 20300 40404 20356
rect 40796 20524 40852 20580
rect 40796 20188 40852 20244
rect 40572 19906 40628 19908
rect 40572 19854 40574 19906
rect 40574 19854 40626 19906
rect 40626 19854 40628 19906
rect 40572 19852 40628 19854
rect 40236 18844 40292 18900
rect 40348 19068 40404 19124
rect 40012 16940 40068 16996
rect 40684 18844 40740 18900
rect 40572 18562 40628 18564
rect 40572 18510 40574 18562
rect 40574 18510 40626 18562
rect 40626 18510 40628 18562
rect 40572 18508 40628 18510
rect 40348 17890 40404 17892
rect 40348 17838 40350 17890
rect 40350 17838 40402 17890
rect 40402 17838 40404 17890
rect 40348 17836 40404 17838
rect 40348 17052 40404 17108
rect 40124 16828 40180 16884
rect 39340 16268 39396 16324
rect 38556 15484 38612 15540
rect 38668 15708 38724 15764
rect 37772 13580 37828 13636
rect 38668 14812 38724 14868
rect 38892 14700 38948 14756
rect 38444 14642 38500 14644
rect 38444 14590 38446 14642
rect 38446 14590 38498 14642
rect 38498 14590 38500 14642
rect 38444 14588 38500 14590
rect 38668 14476 38724 14532
rect 39004 14418 39060 14420
rect 39004 14366 39006 14418
rect 39006 14366 39058 14418
rect 39058 14366 39060 14418
rect 39004 14364 39060 14366
rect 38780 13634 38836 13636
rect 38780 13582 38782 13634
rect 38782 13582 38834 13634
rect 38834 13582 38836 13634
rect 38780 13580 38836 13582
rect 38668 13468 38724 13524
rect 38556 13356 38612 13412
rect 37772 11506 37828 11508
rect 37772 11454 37774 11506
rect 37774 11454 37826 11506
rect 37826 11454 37828 11506
rect 37772 11452 37828 11454
rect 37212 7756 37268 7812
rect 37772 9042 37828 9044
rect 37772 8990 37774 9042
rect 37774 8990 37826 9042
rect 37826 8990 37828 9042
rect 37772 8988 37828 8990
rect 37436 8876 37492 8932
rect 37772 6636 37828 6692
rect 37772 6076 37828 6132
rect 37436 5122 37492 5124
rect 37436 5070 37438 5122
rect 37438 5070 37490 5122
rect 37490 5070 37492 5122
rect 37436 5068 37492 5070
rect 37324 3836 37380 3892
rect 37660 3330 37716 3332
rect 37660 3278 37662 3330
rect 37662 3278 37714 3330
rect 37714 3278 37716 3330
rect 37660 3276 37716 3278
rect 37100 2828 37156 2884
rect 37996 11340 38052 11396
rect 37996 10444 38052 10500
rect 38668 12572 38724 12628
rect 38780 11788 38836 11844
rect 38668 11394 38724 11396
rect 38668 11342 38670 11394
rect 38670 11342 38722 11394
rect 38722 11342 38724 11394
rect 38668 11340 38724 11342
rect 38892 11452 38948 11508
rect 39004 14140 39060 14196
rect 39228 15538 39284 15540
rect 39228 15486 39230 15538
rect 39230 15486 39282 15538
rect 39282 15486 39284 15538
rect 39228 15484 39284 15486
rect 39676 16268 39732 16324
rect 39900 15874 39956 15876
rect 39900 15822 39902 15874
rect 39902 15822 39954 15874
rect 39954 15822 39956 15874
rect 39900 15820 39956 15822
rect 39564 15538 39620 15540
rect 39564 15486 39566 15538
rect 39566 15486 39618 15538
rect 39618 15486 39620 15538
rect 39564 15484 39620 15486
rect 40236 16940 40292 16996
rect 40348 16882 40404 16884
rect 40348 16830 40350 16882
rect 40350 16830 40402 16882
rect 40402 16830 40404 16882
rect 40348 16828 40404 16830
rect 39116 13356 39172 13412
rect 39116 12962 39172 12964
rect 39116 12910 39118 12962
rect 39118 12910 39170 12962
rect 39170 12910 39172 12962
rect 39116 12908 39172 12910
rect 39788 14642 39844 14644
rect 39788 14590 39790 14642
rect 39790 14590 39842 14642
rect 39842 14590 39844 14642
rect 39788 14588 39844 14590
rect 39340 14140 39396 14196
rect 39788 13468 39844 13524
rect 39676 13356 39732 13412
rect 39676 13020 39732 13076
rect 39452 12850 39508 12852
rect 39452 12798 39454 12850
rect 39454 12798 39506 12850
rect 39506 12798 39508 12850
rect 39452 12796 39508 12798
rect 39116 11788 39172 11844
rect 39452 11788 39508 11844
rect 38220 10498 38276 10500
rect 38220 10446 38222 10498
rect 38222 10446 38274 10498
rect 38274 10446 38276 10498
rect 38220 10444 38276 10446
rect 37996 7698 38052 7700
rect 37996 7646 37998 7698
rect 37998 7646 38050 7698
rect 38050 7646 38052 7698
rect 37996 7644 38052 7646
rect 38332 8204 38388 8260
rect 38332 7308 38388 7364
rect 38220 6690 38276 6692
rect 38220 6638 38222 6690
rect 38222 6638 38274 6690
rect 38274 6638 38276 6690
rect 38220 6636 38276 6638
rect 39452 10498 39508 10500
rect 39452 10446 39454 10498
rect 39454 10446 39506 10498
rect 39506 10446 39508 10498
rect 39452 10444 39508 10446
rect 40124 14140 40180 14196
rect 40796 17778 40852 17780
rect 40796 17726 40798 17778
rect 40798 17726 40850 17778
rect 40850 17726 40852 17778
rect 40796 17724 40852 17726
rect 41020 17554 41076 17556
rect 41020 17502 41022 17554
rect 41022 17502 41074 17554
rect 41074 17502 41076 17554
rect 41020 17500 41076 17502
rect 40572 16770 40628 16772
rect 40572 16718 40574 16770
rect 40574 16718 40626 16770
rect 40626 16718 40628 16770
rect 40572 16716 40628 16718
rect 41020 16828 41076 16884
rect 40572 16492 40628 16548
rect 40460 16268 40516 16324
rect 40460 15260 40516 15316
rect 40460 14530 40516 14532
rect 40460 14478 40462 14530
rect 40462 14478 40514 14530
rect 40514 14478 40516 14530
rect 40460 14476 40516 14478
rect 40908 16322 40964 16324
rect 40908 16270 40910 16322
rect 40910 16270 40962 16322
rect 40962 16270 40964 16322
rect 40908 16268 40964 16270
rect 41020 15932 41076 15988
rect 40684 15538 40740 15540
rect 40684 15486 40686 15538
rect 40686 15486 40738 15538
rect 40738 15486 40740 15538
rect 40684 15484 40740 15486
rect 40348 13468 40404 13524
rect 40684 15260 40740 15316
rect 40236 12962 40292 12964
rect 40236 12910 40238 12962
rect 40238 12910 40290 12962
rect 40290 12910 40292 12962
rect 40236 12908 40292 12910
rect 40124 12738 40180 12740
rect 40124 12686 40126 12738
rect 40126 12686 40178 12738
rect 40178 12686 40180 12738
rect 40124 12684 40180 12686
rect 40124 11788 40180 11844
rect 39788 10444 39844 10500
rect 38668 9826 38724 9828
rect 38668 9774 38670 9826
rect 38670 9774 38722 9826
rect 38722 9774 38724 9826
rect 38668 9772 38724 9774
rect 39116 8540 39172 8596
rect 38668 7644 38724 7700
rect 39564 8204 39620 8260
rect 39564 7756 39620 7812
rect 38444 6636 38500 6692
rect 38780 7308 38836 7364
rect 40012 7362 40068 7364
rect 40012 7310 40014 7362
rect 40014 7310 40066 7362
rect 40066 7310 40068 7362
rect 40012 7308 40068 7310
rect 40572 13356 40628 13412
rect 40572 12402 40628 12404
rect 40572 12350 40574 12402
rect 40574 12350 40626 12402
rect 40626 12350 40628 12402
rect 40572 12348 40628 12350
rect 41468 21868 41524 21924
rect 41244 20802 41300 20804
rect 41244 20750 41246 20802
rect 41246 20750 41298 20802
rect 41298 20750 41300 20802
rect 41244 20748 41300 20750
rect 42140 22988 42196 23044
rect 41916 22428 41972 22484
rect 41916 21810 41972 21812
rect 41916 21758 41918 21810
rect 41918 21758 41970 21810
rect 41970 21758 41972 21810
rect 41916 21756 41972 21758
rect 41804 21026 41860 21028
rect 41804 20974 41806 21026
rect 41806 20974 41858 21026
rect 41858 20974 41860 21026
rect 41804 20972 41860 20974
rect 41468 19346 41524 19348
rect 41468 19294 41470 19346
rect 41470 19294 41522 19346
rect 41522 19294 41524 19346
rect 41468 19292 41524 19294
rect 41804 20188 41860 20244
rect 41692 19404 41748 19460
rect 41580 18620 41636 18676
rect 42140 21420 42196 21476
rect 41916 19068 41972 19124
rect 42252 20972 42308 21028
rect 42924 27858 42980 27860
rect 42924 27806 42926 27858
rect 42926 27806 42978 27858
rect 42978 27806 42980 27858
rect 42924 27804 42980 27806
rect 43036 27580 43092 27636
rect 42812 26684 42868 26740
rect 43708 31948 43764 32004
rect 43820 32284 43876 32340
rect 43820 31612 43876 31668
rect 44268 32562 44324 32564
rect 44268 32510 44270 32562
rect 44270 32510 44322 32562
rect 44322 32510 44324 32562
rect 44268 32508 44324 32510
rect 44044 31836 44100 31892
rect 44156 31778 44212 31780
rect 44156 31726 44158 31778
rect 44158 31726 44210 31778
rect 44210 31726 44212 31778
rect 44156 31724 44212 31726
rect 43932 31388 43988 31444
rect 43820 30940 43876 30996
rect 43596 30044 43652 30100
rect 44268 31554 44324 31556
rect 44268 31502 44270 31554
rect 44270 31502 44322 31554
rect 44322 31502 44324 31554
rect 44268 31500 44324 31502
rect 44268 31164 44324 31220
rect 45164 34524 45220 34580
rect 45052 34412 45108 34468
rect 45052 34018 45108 34020
rect 45052 33966 45054 34018
rect 45054 33966 45106 34018
rect 45106 33966 45108 34018
rect 45052 33964 45108 33966
rect 44492 32844 44548 32900
rect 44604 32284 44660 32340
rect 44492 31948 44548 32004
rect 44828 32396 44884 32452
rect 43932 30604 43988 30660
rect 43820 30044 43876 30100
rect 43484 29708 43540 29764
rect 43260 29148 43316 29204
rect 43260 27020 43316 27076
rect 43372 26908 43428 26964
rect 43820 29596 43876 29652
rect 43596 29148 43652 29204
rect 43596 28252 43652 28308
rect 43596 27692 43652 27748
rect 43596 27020 43652 27076
rect 43708 27468 43764 27524
rect 43260 25676 43316 25732
rect 42924 25394 42980 25396
rect 42924 25342 42926 25394
rect 42926 25342 42978 25394
rect 42978 25342 42980 25394
rect 42924 25340 42980 25342
rect 42812 25282 42868 25284
rect 42812 25230 42814 25282
rect 42814 25230 42866 25282
rect 42866 25230 42868 25282
rect 42812 25228 42868 25230
rect 43036 25282 43092 25284
rect 43036 25230 43038 25282
rect 43038 25230 43090 25282
rect 43090 25230 43092 25282
rect 43036 25228 43092 25230
rect 43036 25004 43092 25060
rect 42812 24556 42868 24612
rect 42588 23996 42644 24052
rect 42700 24108 42756 24164
rect 42476 23436 42532 23492
rect 42476 23100 42532 23156
rect 42588 22540 42644 22596
rect 42812 23660 42868 23716
rect 42364 20860 42420 20916
rect 42476 21532 42532 21588
rect 42588 21644 42644 21700
rect 42588 21420 42644 21476
rect 42812 20802 42868 20804
rect 42812 20750 42814 20802
rect 42814 20750 42866 20802
rect 42866 20750 42868 20802
rect 42812 20748 42868 20750
rect 42700 20636 42756 20692
rect 42476 20412 42532 20468
rect 42812 20188 42868 20244
rect 42028 19852 42084 19908
rect 42588 19964 42644 20020
rect 41468 17612 41524 17668
rect 41132 16716 41188 16772
rect 41468 16716 41524 16772
rect 42252 18396 42308 18452
rect 41916 18226 41972 18228
rect 41916 18174 41918 18226
rect 41918 18174 41970 18226
rect 41970 18174 41972 18226
rect 41916 18172 41972 18174
rect 42252 18172 42308 18228
rect 41804 18060 41860 18116
rect 41692 16940 41748 16996
rect 41804 17724 41860 17780
rect 41580 16828 41636 16884
rect 41132 15820 41188 15876
rect 41244 15260 41300 15316
rect 40796 15036 40852 15092
rect 41132 14364 41188 14420
rect 40908 13356 40964 13412
rect 41020 12962 41076 12964
rect 41020 12910 41022 12962
rect 41022 12910 41074 12962
rect 41074 12910 41076 12962
rect 41020 12908 41076 12910
rect 40908 12850 40964 12852
rect 40908 12798 40910 12850
rect 40910 12798 40962 12850
rect 40962 12798 40964 12850
rect 40908 12796 40964 12798
rect 41132 12796 41188 12852
rect 41020 12236 41076 12292
rect 40908 11116 40964 11172
rect 40348 9548 40404 9604
rect 41692 14418 41748 14420
rect 41692 14366 41694 14418
rect 41694 14366 41746 14418
rect 41746 14366 41748 14418
rect 41692 14364 41748 14366
rect 41916 17666 41972 17668
rect 41916 17614 41918 17666
rect 41918 17614 41970 17666
rect 41970 17614 41972 17666
rect 41916 17612 41972 17614
rect 42140 17500 42196 17556
rect 41916 17106 41972 17108
rect 41916 17054 41918 17106
rect 41918 17054 41970 17106
rect 41970 17054 41972 17106
rect 41916 17052 41972 17054
rect 42700 19628 42756 19684
rect 43372 26572 43428 26628
rect 43372 25004 43428 25060
rect 43708 26796 43764 26852
rect 44156 29820 44212 29876
rect 44156 28924 44212 28980
rect 43932 26796 43988 26852
rect 43820 26402 43876 26404
rect 43820 26350 43822 26402
rect 43822 26350 43874 26402
rect 43874 26350 43876 26402
rect 43820 26348 43876 26350
rect 43820 25788 43876 25844
rect 44044 26514 44100 26516
rect 44044 26462 44046 26514
rect 44046 26462 44098 26514
rect 44098 26462 44100 26514
rect 44044 26460 44100 26462
rect 44604 30604 44660 30660
rect 45164 33628 45220 33684
rect 46396 37378 46452 37380
rect 46396 37326 46398 37378
rect 46398 37326 46450 37378
rect 46450 37326 46452 37378
rect 46396 37324 46452 37326
rect 46284 37212 46340 37268
rect 46172 36988 46228 37044
rect 45500 36706 45556 36708
rect 45500 36654 45502 36706
rect 45502 36654 45554 36706
rect 45554 36654 45556 36706
rect 45500 36652 45556 36654
rect 45836 36482 45892 36484
rect 45836 36430 45838 36482
rect 45838 36430 45890 36482
rect 45890 36430 45892 36482
rect 45836 36428 45892 36430
rect 45948 36204 46004 36260
rect 46060 35420 46116 35476
rect 45500 33628 45556 33684
rect 45612 34636 45668 34692
rect 45388 33404 45444 33460
rect 45052 32060 45108 32116
rect 45052 31836 45108 31892
rect 44940 31218 44996 31220
rect 44940 31166 44942 31218
rect 44942 31166 44994 31218
rect 44994 31166 44996 31218
rect 44940 31164 44996 31166
rect 44828 31052 44884 31108
rect 45164 30604 45220 30660
rect 45276 31948 45332 32004
rect 44940 29820 44996 29876
rect 44380 28642 44436 28644
rect 44380 28590 44382 28642
rect 44382 28590 44434 28642
rect 44434 28590 44436 28642
rect 44380 28588 44436 28590
rect 44268 27244 44324 27300
rect 44716 27692 44772 27748
rect 44828 27916 44884 27972
rect 44492 27132 44548 27188
rect 44268 26572 44324 26628
rect 44380 26460 44436 26516
rect 44492 25676 44548 25732
rect 43596 24332 43652 24388
rect 43708 25116 43764 25172
rect 43148 23714 43204 23716
rect 43148 23662 43150 23714
rect 43150 23662 43202 23714
rect 43202 23662 43204 23714
rect 43148 23660 43204 23662
rect 43260 22764 43316 22820
rect 43708 23884 43764 23940
rect 43484 23154 43540 23156
rect 43484 23102 43486 23154
rect 43486 23102 43538 23154
rect 43538 23102 43540 23154
rect 43484 23100 43540 23102
rect 44156 25340 44212 25396
rect 43708 22540 43764 22596
rect 43036 20802 43092 20804
rect 43036 20750 43038 20802
rect 43038 20750 43090 20802
rect 43090 20750 43092 20802
rect 43036 20748 43092 20750
rect 43036 20412 43092 20468
rect 42924 19628 42980 19684
rect 42812 19516 42868 19572
rect 42924 19068 42980 19124
rect 42476 18732 42532 18788
rect 42588 18508 42644 18564
rect 43148 18956 43204 19012
rect 43036 18338 43092 18340
rect 43036 18286 43038 18338
rect 43038 18286 43090 18338
rect 43090 18286 43092 18338
rect 43036 18284 43092 18286
rect 43372 22316 43428 22372
rect 43708 20748 43764 20804
rect 43596 20690 43652 20692
rect 43596 20638 43598 20690
rect 43598 20638 43650 20690
rect 43650 20638 43652 20690
rect 43596 20636 43652 20638
rect 43596 20076 43652 20132
rect 43484 19740 43540 19796
rect 43260 18172 43316 18228
rect 42364 16156 42420 16212
rect 42476 16716 42532 16772
rect 42028 15986 42084 15988
rect 42028 15934 42030 15986
rect 42030 15934 42082 15986
rect 42082 15934 42084 15986
rect 42028 15932 42084 15934
rect 42252 15372 42308 15428
rect 42364 15596 42420 15652
rect 42028 15314 42084 15316
rect 42028 15262 42030 15314
rect 42030 15262 42082 15314
rect 42082 15262 42084 15314
rect 42028 15260 42084 15262
rect 42028 14364 42084 14420
rect 41244 9996 41300 10052
rect 41356 13580 41412 13636
rect 41020 9602 41076 9604
rect 41020 9550 41022 9602
rect 41022 9550 41074 9602
rect 41074 9550 41076 9602
rect 41020 9548 41076 9550
rect 40460 9100 40516 9156
rect 40908 8428 40964 8484
rect 41132 9436 41188 9492
rect 40572 6412 40628 6468
rect 37996 5180 38052 5236
rect 40124 4508 40180 4564
rect 40236 5628 40292 5684
rect 39564 4338 39620 4340
rect 39564 4286 39566 4338
rect 39566 4286 39618 4338
rect 39618 4286 39620 4338
rect 39564 4284 39620 4286
rect 40796 5852 40852 5908
rect 40796 5068 40852 5124
rect 40460 4562 40516 4564
rect 40460 4510 40462 4562
rect 40462 4510 40514 4562
rect 40514 4510 40516 4562
rect 40460 4508 40516 4510
rect 40236 4060 40292 4116
rect 38444 3836 38500 3892
rect 39228 3612 39284 3668
rect 41580 12684 41636 12740
rect 41468 12402 41524 12404
rect 41468 12350 41470 12402
rect 41470 12350 41522 12402
rect 41522 12350 41524 12402
rect 41468 12348 41524 12350
rect 41468 12012 41524 12068
rect 43372 17612 43428 17668
rect 43596 19292 43652 19348
rect 43596 18620 43652 18676
rect 43372 17164 43428 17220
rect 42700 16492 42756 16548
rect 42252 13916 42308 13972
rect 42028 13132 42084 13188
rect 41804 12796 41860 12852
rect 42700 14140 42756 14196
rect 43260 15596 43316 15652
rect 42924 15260 42980 15316
rect 43036 15202 43092 15204
rect 43036 15150 43038 15202
rect 43038 15150 43090 15202
rect 43090 15150 43092 15202
rect 43036 15148 43092 15150
rect 42924 14418 42980 14420
rect 42924 14366 42926 14418
rect 42926 14366 42978 14418
rect 42978 14366 42980 14418
rect 42924 14364 42980 14366
rect 42700 13634 42756 13636
rect 42700 13582 42702 13634
rect 42702 13582 42754 13634
rect 42754 13582 42756 13634
rect 42700 13580 42756 13582
rect 43036 13020 43092 13076
rect 42364 12236 42420 12292
rect 41804 11618 41860 11620
rect 41804 11566 41806 11618
rect 41806 11566 41858 11618
rect 41858 11566 41860 11618
rect 41804 11564 41860 11566
rect 41692 11452 41748 11508
rect 42252 11506 42308 11508
rect 42252 11454 42254 11506
rect 42254 11454 42306 11506
rect 42306 11454 42308 11506
rect 42252 11452 42308 11454
rect 41916 9996 41972 10052
rect 42140 9602 42196 9604
rect 42140 9550 42142 9602
rect 42142 9550 42194 9602
rect 42194 9550 42196 9602
rect 42140 9548 42196 9550
rect 41804 9324 41860 9380
rect 41356 8988 41412 9044
rect 41356 8428 41412 8484
rect 42700 12290 42756 12292
rect 42700 12238 42702 12290
rect 42702 12238 42754 12290
rect 42754 12238 42756 12290
rect 42700 12236 42756 12238
rect 42588 11170 42644 11172
rect 42588 11118 42590 11170
rect 42590 11118 42642 11170
rect 42642 11118 42644 11170
rect 42588 11116 42644 11118
rect 42588 10892 42644 10948
rect 42588 9154 42644 9156
rect 42588 9102 42590 9154
rect 42590 9102 42642 9154
rect 42642 9102 42644 9154
rect 42588 9100 42644 9102
rect 41804 8146 41860 8148
rect 41804 8094 41806 8146
rect 41806 8094 41858 8146
rect 41858 8094 41860 8146
rect 41804 8092 41860 8094
rect 43484 16380 43540 16436
rect 43596 16098 43652 16100
rect 43596 16046 43598 16098
rect 43598 16046 43650 16098
rect 43650 16046 43652 16098
rect 43596 16044 43652 16046
rect 43932 25282 43988 25284
rect 43932 25230 43934 25282
rect 43934 25230 43986 25282
rect 43986 25230 43988 25282
rect 43932 25228 43988 25230
rect 44156 24722 44212 24724
rect 44156 24670 44158 24722
rect 44158 24670 44210 24722
rect 44210 24670 44212 24722
rect 44156 24668 44212 24670
rect 44492 24108 44548 24164
rect 44044 23938 44100 23940
rect 44044 23886 44046 23938
rect 44046 23886 44098 23938
rect 44098 23886 44100 23938
rect 44044 23884 44100 23886
rect 44380 22988 44436 23044
rect 44380 22428 44436 22484
rect 43932 21420 43988 21476
rect 44492 22316 44548 22372
rect 44156 21644 44212 21700
rect 44044 20972 44100 21028
rect 43932 20578 43988 20580
rect 43932 20526 43934 20578
rect 43934 20526 43986 20578
rect 43986 20526 43988 20578
rect 43932 20524 43988 20526
rect 43820 19234 43876 19236
rect 43820 19182 43822 19234
rect 43822 19182 43874 19234
rect 43874 19182 43876 19234
rect 43820 19180 43876 19182
rect 43820 17276 43876 17332
rect 44268 20636 44324 20692
rect 44268 20018 44324 20020
rect 44268 19966 44270 20018
rect 44270 19966 44322 20018
rect 44322 19966 44324 20018
rect 44268 19964 44324 19966
rect 44044 19740 44100 19796
rect 45164 27916 45220 27972
rect 44940 27020 44996 27076
rect 45164 26684 45220 26740
rect 44716 26348 44772 26404
rect 44828 22988 44884 23044
rect 44716 22204 44772 22260
rect 44716 21868 44772 21924
rect 44604 20300 44660 20356
rect 44380 19628 44436 19684
rect 44604 19740 44660 19796
rect 44268 19516 44324 19572
rect 44156 19346 44212 19348
rect 44156 19294 44158 19346
rect 44158 19294 44210 19346
rect 44210 19294 44212 19346
rect 44156 19292 44212 19294
rect 44268 18562 44324 18564
rect 44268 18510 44270 18562
rect 44270 18510 44322 18562
rect 44322 18510 44324 18562
rect 44268 18508 44324 18510
rect 44716 19010 44772 19012
rect 44716 18958 44718 19010
rect 44718 18958 44770 19010
rect 44770 18958 44772 19010
rect 44716 18956 44772 18958
rect 44940 25452 44996 25508
rect 45052 25340 45108 25396
rect 45612 32508 45668 32564
rect 45724 31948 45780 32004
rect 45500 31836 45556 31892
rect 46844 37772 46900 37828
rect 46620 37100 46676 37156
rect 46732 35868 46788 35924
rect 47180 36988 47236 37044
rect 47740 41074 47796 41076
rect 47740 41022 47742 41074
rect 47742 41022 47794 41074
rect 47794 41022 47796 41074
rect 47740 41020 47796 41022
rect 47740 40460 47796 40516
rect 48524 43538 48580 43540
rect 48524 43486 48526 43538
rect 48526 43486 48578 43538
rect 48578 43486 48580 43538
rect 48524 43484 48580 43486
rect 49084 43484 49140 43540
rect 49196 43596 49252 43652
rect 48524 42028 48580 42084
rect 48524 41244 48580 41300
rect 48076 40962 48132 40964
rect 48076 40910 48078 40962
rect 48078 40910 48130 40962
rect 48130 40910 48132 40962
rect 48076 40908 48132 40910
rect 47964 40572 48020 40628
rect 48188 40572 48244 40628
rect 48748 40626 48804 40628
rect 48748 40574 48750 40626
rect 48750 40574 48802 40626
rect 48802 40574 48804 40626
rect 48748 40572 48804 40574
rect 48524 40348 48580 40404
rect 48524 39394 48580 39396
rect 48524 39342 48526 39394
rect 48526 39342 48578 39394
rect 48578 39342 48580 39394
rect 48524 39340 48580 39342
rect 49980 49532 50036 49588
rect 49532 49308 49588 49364
rect 49532 49026 49588 49028
rect 49532 48974 49534 49026
rect 49534 48974 49586 49026
rect 49586 48974 49588 49026
rect 49532 48972 49588 48974
rect 49756 48412 49812 48468
rect 49644 46674 49700 46676
rect 49644 46622 49646 46674
rect 49646 46622 49698 46674
rect 49698 46622 49700 46674
rect 49644 46620 49700 46622
rect 49868 48300 49924 48356
rect 49868 47068 49924 47124
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 50988 49868 51044 49924
rect 50764 48860 50820 48916
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 49532 45778 49588 45780
rect 49532 45726 49534 45778
rect 49534 45726 49586 45778
rect 49586 45726 49588 45778
rect 49532 45724 49588 45726
rect 49532 45388 49588 45444
rect 49420 43426 49476 43428
rect 49420 43374 49422 43426
rect 49422 43374 49474 43426
rect 49474 43374 49476 43426
rect 49420 43372 49476 43374
rect 49644 43372 49700 43428
rect 49868 46620 49924 46676
rect 50428 47292 50484 47348
rect 50204 47068 50260 47124
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 50316 46562 50372 46564
rect 50316 46510 50318 46562
rect 50318 46510 50370 46562
rect 50370 46510 50372 46562
rect 50316 46508 50372 46510
rect 50764 46508 50820 46564
rect 50764 46172 50820 46228
rect 49980 45164 50036 45220
rect 50092 45836 50148 45892
rect 50204 44716 50260 44772
rect 50204 44380 50260 44436
rect 50876 46396 50932 46452
rect 51324 49868 51380 49924
rect 51660 49980 51716 50036
rect 51100 48412 51156 48468
rect 51324 48354 51380 48356
rect 51324 48302 51326 48354
rect 51326 48302 51378 48354
rect 51378 48302 51380 48354
rect 51324 48300 51380 48302
rect 50988 46060 51044 46116
rect 51100 47292 51156 47348
rect 50876 45612 50932 45668
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50428 45276 50484 45332
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50204 43596 50260 43652
rect 50316 43708 50372 43764
rect 49756 43260 49812 43316
rect 49420 42028 49476 42084
rect 49756 40572 49812 40628
rect 50092 42866 50148 42868
rect 50092 42814 50094 42866
rect 50094 42814 50146 42866
rect 50146 42814 50148 42866
rect 50092 42812 50148 42814
rect 50876 43596 50932 43652
rect 50988 43708 51044 43764
rect 50316 43148 50372 43204
rect 50428 43484 50484 43540
rect 51996 49698 52052 49700
rect 51996 49646 51998 49698
rect 51998 49646 52050 49698
rect 52050 49646 52052 49698
rect 51996 49644 52052 49646
rect 51996 49308 52052 49364
rect 51436 47292 51492 47348
rect 51548 48242 51604 48244
rect 51548 48190 51550 48242
rect 51550 48190 51602 48242
rect 51602 48190 51604 48242
rect 51548 48188 51604 48190
rect 51548 47458 51604 47460
rect 51548 47406 51550 47458
rect 51550 47406 51602 47458
rect 51602 47406 51604 47458
rect 51548 47404 51604 47406
rect 51660 47740 51716 47796
rect 51212 46562 51268 46564
rect 51212 46510 51214 46562
rect 51214 46510 51266 46562
rect 51266 46510 51268 46562
rect 51212 46508 51268 46510
rect 51212 46060 51268 46116
rect 51100 43484 51156 43540
rect 51212 44604 51268 44660
rect 51100 43036 51156 43092
rect 49868 40908 49924 40964
rect 50428 42642 50484 42644
rect 50428 42590 50430 42642
rect 50430 42590 50482 42642
rect 50482 42590 50484 42642
rect 50428 42588 50484 42590
rect 49532 40514 49588 40516
rect 49532 40462 49534 40514
rect 49534 40462 49586 40514
rect 49586 40462 49588 40514
rect 49532 40460 49588 40462
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 51324 43708 51380 43764
rect 51436 46284 51492 46340
rect 51436 45388 51492 45444
rect 51324 43538 51380 43540
rect 51324 43486 51326 43538
rect 51326 43486 51378 43538
rect 51378 43486 51380 43538
rect 51324 43484 51380 43486
rect 50204 42028 50260 42084
rect 49084 39618 49140 39620
rect 49084 39566 49086 39618
rect 49086 39566 49138 39618
rect 49138 39566 49140 39618
rect 49084 39564 49140 39566
rect 47292 36652 47348 36708
rect 47516 37324 47572 37380
rect 47292 36370 47348 36372
rect 47292 36318 47294 36370
rect 47294 36318 47346 36370
rect 47346 36318 47348 36370
rect 47292 36316 47348 36318
rect 47180 35980 47236 36036
rect 46396 34354 46452 34356
rect 46396 34302 46398 34354
rect 46398 34302 46450 34354
rect 46450 34302 46452 34354
rect 46396 34300 46452 34302
rect 46284 34076 46340 34132
rect 46844 35196 46900 35252
rect 46844 34524 46900 34580
rect 47292 34412 47348 34468
rect 46844 34076 46900 34132
rect 46620 33404 46676 33460
rect 46508 32844 46564 32900
rect 46284 32060 46340 32116
rect 46508 31948 46564 32004
rect 45948 31500 46004 31556
rect 45388 31164 45444 31220
rect 45836 31218 45892 31220
rect 45836 31166 45838 31218
rect 45838 31166 45890 31218
rect 45890 31166 45892 31218
rect 45836 31164 45892 31166
rect 45724 30268 45780 30324
rect 45500 30044 45556 30100
rect 45388 29986 45444 29988
rect 45388 29934 45390 29986
rect 45390 29934 45442 29986
rect 45442 29934 45444 29986
rect 45388 29932 45444 29934
rect 45388 28812 45444 28868
rect 45388 27468 45444 27524
rect 45500 26684 45556 26740
rect 46284 31890 46340 31892
rect 46284 31838 46286 31890
rect 46286 31838 46338 31890
rect 46338 31838 46340 31890
rect 46284 31836 46340 31838
rect 46732 31500 46788 31556
rect 46284 31276 46340 31332
rect 46284 30882 46340 30884
rect 46284 30830 46286 30882
rect 46286 30830 46338 30882
rect 46338 30830 46340 30882
rect 46284 30828 46340 30830
rect 46172 30210 46228 30212
rect 46172 30158 46174 30210
rect 46174 30158 46226 30210
rect 46226 30158 46228 30210
rect 46172 30156 46228 30158
rect 45724 27916 45780 27972
rect 45948 27746 46004 27748
rect 45948 27694 45950 27746
rect 45950 27694 46002 27746
rect 46002 27694 46004 27746
rect 45948 27692 46004 27694
rect 45612 26348 45668 26404
rect 45612 26012 45668 26068
rect 45612 25618 45668 25620
rect 45612 25566 45614 25618
rect 45614 25566 45666 25618
rect 45666 25566 45668 25618
rect 45612 25564 45668 25566
rect 45948 27468 46004 27524
rect 45164 24556 45220 24612
rect 45052 23154 45108 23156
rect 45052 23102 45054 23154
rect 45054 23102 45106 23154
rect 45106 23102 45108 23154
rect 45052 23100 45108 23102
rect 45500 23996 45556 24052
rect 45836 25452 45892 25508
rect 46060 26348 46116 26404
rect 46172 26684 46228 26740
rect 46172 25900 46228 25956
rect 46060 25228 46116 25284
rect 45500 23714 45556 23716
rect 45500 23662 45502 23714
rect 45502 23662 45554 23714
rect 45554 23662 45556 23714
rect 45500 23660 45556 23662
rect 45276 22204 45332 22260
rect 45276 21980 45332 22036
rect 45500 22316 45556 22372
rect 45388 20914 45444 20916
rect 45388 20862 45390 20914
rect 45390 20862 45442 20914
rect 45442 20862 45444 20914
rect 45388 20860 45444 20862
rect 44940 20076 44996 20132
rect 45276 20748 45332 20804
rect 45164 19628 45220 19684
rect 45388 19292 45444 19348
rect 44940 19180 44996 19236
rect 45164 19180 45220 19236
rect 44156 18226 44212 18228
rect 44156 18174 44158 18226
rect 44158 18174 44210 18226
rect 44210 18174 44212 18226
rect 44156 18172 44212 18174
rect 44604 18060 44660 18116
rect 44044 17836 44100 17892
rect 44156 17948 44212 18004
rect 44380 17948 44436 18004
rect 44268 17388 44324 17444
rect 44156 16940 44212 16996
rect 44716 17666 44772 17668
rect 44716 17614 44718 17666
rect 44718 17614 44770 17666
rect 44770 17614 44772 17666
rect 44716 17612 44772 17614
rect 44716 16940 44772 16996
rect 43708 15314 43764 15316
rect 43708 15262 43710 15314
rect 43710 15262 43762 15314
rect 43762 15262 43764 15314
rect 43708 15260 43764 15262
rect 43932 15202 43988 15204
rect 43932 15150 43934 15202
rect 43934 15150 43986 15202
rect 43986 15150 43988 15202
rect 43932 15148 43988 15150
rect 43484 15036 43540 15092
rect 43484 14812 43540 14868
rect 43932 14812 43988 14868
rect 43708 14418 43764 14420
rect 43708 14366 43710 14418
rect 43710 14366 43762 14418
rect 43762 14366 43764 14418
rect 43708 14364 43764 14366
rect 43484 13970 43540 13972
rect 43484 13918 43486 13970
rect 43486 13918 43538 13970
rect 43538 13918 43540 13970
rect 43484 13916 43540 13918
rect 43820 14140 43876 14196
rect 43484 13356 43540 13412
rect 43036 11506 43092 11508
rect 43036 11454 43038 11506
rect 43038 11454 43090 11506
rect 43090 11454 43092 11506
rect 43036 11452 43092 11454
rect 43596 12460 43652 12516
rect 43708 12348 43764 12404
rect 43708 11900 43764 11956
rect 43036 10444 43092 10500
rect 43260 8370 43316 8372
rect 43260 8318 43262 8370
rect 43262 8318 43314 8370
rect 43314 8318 43316 8370
rect 43260 8316 43316 8318
rect 42700 8092 42756 8148
rect 41356 6466 41412 6468
rect 41356 6414 41358 6466
rect 41358 6414 41410 6466
rect 41410 6414 41412 6466
rect 41356 6412 41412 6414
rect 41468 5906 41524 5908
rect 41468 5854 41470 5906
rect 41470 5854 41522 5906
rect 41522 5854 41524 5906
rect 41468 5852 41524 5854
rect 41356 5740 41412 5796
rect 40908 3612 40964 3668
rect 42028 5740 42084 5796
rect 41916 5292 41972 5348
rect 41916 4732 41972 4788
rect 42588 7308 42644 7364
rect 43484 9884 43540 9940
rect 43596 9996 43652 10052
rect 44604 16604 44660 16660
rect 44492 16210 44548 16212
rect 44492 16158 44494 16210
rect 44494 16158 44546 16210
rect 44546 16158 44548 16210
rect 44492 16156 44548 16158
rect 44380 15538 44436 15540
rect 44380 15486 44382 15538
rect 44382 15486 44434 15538
rect 44434 15486 44436 15538
rect 44380 15484 44436 15486
rect 44380 14812 44436 14868
rect 44044 14252 44100 14308
rect 44044 13692 44100 13748
rect 44940 18060 44996 18116
rect 45612 19458 45668 19460
rect 45612 19406 45614 19458
rect 45614 19406 45666 19458
rect 45666 19406 45668 19458
rect 45612 19404 45668 19406
rect 45612 18396 45668 18452
rect 45164 17948 45220 18004
rect 45500 17836 45556 17892
rect 44828 15036 44884 15092
rect 44940 17388 44996 17444
rect 44268 13970 44324 13972
rect 44268 13918 44270 13970
rect 44270 13918 44322 13970
rect 44322 13918 44324 13970
rect 44268 13916 44324 13918
rect 44268 12348 44324 12404
rect 43820 8316 43876 8372
rect 44044 9548 44100 9604
rect 44156 8370 44212 8372
rect 44156 8318 44158 8370
rect 44158 8318 44210 8370
rect 44210 8318 44212 8370
rect 44156 8316 44212 8318
rect 43932 7980 43988 8036
rect 43372 6860 43428 6916
rect 43708 6802 43764 6804
rect 43708 6750 43710 6802
rect 43710 6750 43762 6802
rect 43762 6750 43764 6802
rect 43708 6748 43764 6750
rect 43708 4732 43764 4788
rect 43820 4956 43876 5012
rect 42140 4338 42196 4340
rect 42140 4286 42142 4338
rect 42142 4286 42194 4338
rect 42194 4286 42196 4338
rect 42140 4284 42196 4286
rect 41692 3666 41748 3668
rect 41692 3614 41694 3666
rect 41694 3614 41746 3666
rect 41746 3614 41748 3666
rect 41692 3612 41748 3614
rect 38444 3388 38500 3444
rect 42476 3442 42532 3444
rect 42476 3390 42478 3442
rect 42478 3390 42530 3442
rect 42530 3390 42532 3442
rect 42476 3388 42532 3390
rect 44492 14306 44548 14308
rect 44492 14254 44494 14306
rect 44494 14254 44546 14306
rect 44546 14254 44548 14306
rect 44492 14252 44548 14254
rect 44380 11452 44436 11508
rect 44492 13804 44548 13860
rect 44492 13356 44548 13412
rect 44604 13468 44660 13524
rect 44716 13356 44772 13412
rect 44828 12684 44884 12740
rect 44604 12178 44660 12180
rect 44604 12126 44606 12178
rect 44606 12126 44658 12178
rect 44658 12126 44660 12178
rect 44604 12124 44660 12126
rect 44492 11116 44548 11172
rect 45500 17442 45556 17444
rect 45500 17390 45502 17442
rect 45502 17390 45554 17442
rect 45554 17390 45556 17442
rect 45500 17388 45556 17390
rect 45052 16940 45108 16996
rect 45388 16994 45444 16996
rect 45388 16942 45390 16994
rect 45390 16942 45442 16994
rect 45442 16942 45444 16994
rect 45388 16940 45444 16942
rect 45500 16716 45556 16772
rect 45388 16156 45444 16212
rect 45276 15036 45332 15092
rect 45836 24108 45892 24164
rect 45836 23548 45892 23604
rect 45836 22258 45892 22260
rect 45836 22206 45838 22258
rect 45838 22206 45890 22258
rect 45890 22206 45892 22258
rect 45836 22204 45892 22206
rect 46172 23938 46228 23940
rect 46172 23886 46174 23938
rect 46174 23886 46226 23938
rect 46226 23886 46228 23938
rect 46172 23884 46228 23886
rect 46060 22764 46116 22820
rect 45948 21868 46004 21924
rect 45836 20972 45892 21028
rect 46172 21532 46228 21588
rect 46060 20972 46116 21028
rect 45836 20242 45892 20244
rect 45836 20190 45838 20242
rect 45838 20190 45890 20242
rect 45890 20190 45892 20242
rect 45836 20188 45892 20190
rect 45948 19346 46004 19348
rect 45948 19294 45950 19346
rect 45950 19294 46002 19346
rect 46002 19294 46004 19346
rect 45948 19292 46004 19294
rect 45836 19122 45892 19124
rect 45836 19070 45838 19122
rect 45838 19070 45890 19122
rect 45890 19070 45892 19122
rect 45836 19068 45892 19070
rect 46396 29932 46452 29988
rect 47292 33292 47348 33348
rect 47068 32956 47124 33012
rect 47180 32844 47236 32900
rect 47292 32562 47348 32564
rect 47292 32510 47294 32562
rect 47294 32510 47346 32562
rect 47346 32510 47348 32562
rect 47292 32508 47348 32510
rect 46956 31836 47012 31892
rect 49532 39116 49588 39172
rect 49532 38444 49588 38500
rect 50092 40348 50148 40404
rect 48748 37938 48804 37940
rect 48748 37886 48750 37938
rect 48750 37886 48802 37938
rect 48802 37886 48804 37938
rect 48748 37884 48804 37886
rect 48300 37826 48356 37828
rect 48300 37774 48302 37826
rect 48302 37774 48354 37826
rect 48354 37774 48356 37826
rect 48300 37772 48356 37774
rect 48188 36876 48244 36932
rect 47628 34354 47684 34356
rect 47628 34302 47630 34354
rect 47630 34302 47682 34354
rect 47682 34302 47684 34354
rect 47628 34300 47684 34302
rect 47740 33852 47796 33908
rect 47628 33740 47684 33796
rect 47964 33740 48020 33796
rect 47852 32956 47908 33012
rect 47404 31836 47460 31892
rect 47740 31778 47796 31780
rect 47740 31726 47742 31778
rect 47742 31726 47794 31778
rect 47794 31726 47796 31778
rect 47740 31724 47796 31726
rect 47068 31500 47124 31556
rect 46956 30828 47012 30884
rect 47516 31500 47572 31556
rect 47516 31052 47572 31108
rect 47292 30434 47348 30436
rect 47292 30382 47294 30434
rect 47294 30382 47346 30434
rect 47346 30382 47348 30434
rect 47292 30380 47348 30382
rect 47068 30268 47124 30324
rect 47516 29820 47572 29876
rect 47628 30940 47684 30996
rect 47180 29260 47236 29316
rect 46396 27356 46452 27412
rect 47516 29260 47572 29316
rect 47404 28866 47460 28868
rect 47404 28814 47406 28866
rect 47406 28814 47458 28866
rect 47458 28814 47460 28866
rect 47404 28812 47460 28814
rect 46732 27916 46788 27972
rect 46956 27746 47012 27748
rect 46956 27694 46958 27746
rect 46958 27694 47010 27746
rect 47010 27694 47012 27746
rect 46956 27692 47012 27694
rect 46844 27580 46900 27636
rect 46620 26684 46676 26740
rect 46732 26908 46788 26964
rect 46620 26514 46676 26516
rect 46620 26462 46622 26514
rect 46622 26462 46674 26514
rect 46674 26462 46676 26514
rect 46620 26460 46676 26462
rect 46956 26796 47012 26852
rect 46620 26124 46676 26180
rect 46620 25506 46676 25508
rect 46620 25454 46622 25506
rect 46622 25454 46674 25506
rect 46674 25454 46676 25506
rect 46620 25452 46676 25454
rect 46620 24892 46676 24948
rect 46396 23548 46452 23604
rect 46732 24780 46788 24836
rect 46956 25116 47012 25172
rect 47292 27804 47348 27860
rect 47964 32284 48020 32340
rect 48188 36370 48244 36372
rect 48188 36318 48190 36370
rect 48190 36318 48242 36370
rect 48242 36318 48244 36370
rect 48188 36316 48244 36318
rect 48412 37266 48468 37268
rect 48412 37214 48414 37266
rect 48414 37214 48466 37266
rect 48466 37214 48468 37266
rect 48412 37212 48468 37214
rect 48524 36988 48580 37044
rect 48524 36652 48580 36708
rect 48412 35196 48468 35252
rect 48188 33628 48244 33684
rect 47964 31836 48020 31892
rect 47964 30828 48020 30884
rect 48748 34860 48804 34916
rect 48636 34802 48692 34804
rect 48636 34750 48638 34802
rect 48638 34750 48690 34802
rect 48690 34750 48692 34802
rect 48636 34748 48692 34750
rect 48636 34300 48692 34356
rect 48524 34018 48580 34020
rect 48524 33966 48526 34018
rect 48526 33966 48578 34018
rect 48578 33966 48580 34018
rect 48524 33964 48580 33966
rect 48524 32956 48580 33012
rect 48412 31836 48468 31892
rect 48524 31500 48580 31556
rect 48300 31388 48356 31444
rect 49308 34188 49364 34244
rect 49868 38220 49924 38276
rect 50204 38332 50260 38388
rect 49644 36652 49700 36708
rect 49532 35586 49588 35588
rect 49532 35534 49534 35586
rect 49534 35534 49586 35586
rect 49586 35534 49588 35586
rect 49532 35532 49588 35534
rect 49756 36316 49812 36372
rect 49756 35644 49812 35700
rect 50428 41970 50484 41972
rect 50428 41918 50430 41970
rect 50430 41918 50482 41970
rect 50482 41918 50484 41970
rect 50428 41916 50484 41918
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50764 40402 50820 40404
rect 50764 40350 50766 40402
rect 50766 40350 50818 40402
rect 50818 40350 50820 40402
rect 50764 40348 50820 40350
rect 51100 41970 51156 41972
rect 51100 41918 51102 41970
rect 51102 41918 51154 41970
rect 51154 41918 51156 41970
rect 51100 41916 51156 41918
rect 50876 39564 50932 39620
rect 51100 40348 51156 40404
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50988 39058 51044 39060
rect 50988 39006 50990 39058
rect 50990 39006 51042 39058
rect 51042 39006 51044 39058
rect 50988 39004 51044 39006
rect 50540 38834 50596 38836
rect 50540 38782 50542 38834
rect 50542 38782 50594 38834
rect 50594 38782 50596 38834
rect 50540 38780 50596 38782
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50540 37212 50596 37268
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50540 35810 50596 35812
rect 50540 35758 50542 35810
rect 50542 35758 50594 35810
rect 50594 35758 50596 35810
rect 50540 35756 50596 35758
rect 50204 35644 50260 35700
rect 50428 35698 50484 35700
rect 50428 35646 50430 35698
rect 50430 35646 50482 35698
rect 50482 35646 50484 35698
rect 50428 35644 50484 35646
rect 49980 35532 50036 35588
rect 49644 34242 49700 34244
rect 49644 34190 49646 34242
rect 49646 34190 49698 34242
rect 49698 34190 49700 34242
rect 49644 34188 49700 34190
rect 49420 33964 49476 34020
rect 48188 30716 48244 30772
rect 48188 30268 48244 30324
rect 48300 31052 48356 31108
rect 47964 29650 48020 29652
rect 47964 29598 47966 29650
rect 47966 29598 48018 29650
rect 48018 29598 48020 29650
rect 47964 29596 48020 29598
rect 48076 29538 48132 29540
rect 48076 29486 48078 29538
rect 48078 29486 48130 29538
rect 48130 29486 48132 29538
rect 48076 29484 48132 29486
rect 48300 28588 48356 28644
rect 48076 28028 48132 28084
rect 47740 27858 47796 27860
rect 47740 27806 47742 27858
rect 47742 27806 47794 27858
rect 47794 27806 47796 27858
rect 47740 27804 47796 27806
rect 47852 27298 47908 27300
rect 47852 27246 47854 27298
rect 47854 27246 47906 27298
rect 47906 27246 47908 27298
rect 47852 27244 47908 27246
rect 46844 23548 46900 23604
rect 46508 22930 46564 22932
rect 46508 22878 46510 22930
rect 46510 22878 46562 22930
rect 46562 22878 46564 22930
rect 46508 22876 46564 22878
rect 46396 21868 46452 21924
rect 46284 20188 46340 20244
rect 47404 26684 47460 26740
rect 47740 26402 47796 26404
rect 47740 26350 47742 26402
rect 47742 26350 47794 26402
rect 47794 26350 47796 26402
rect 47740 26348 47796 26350
rect 47852 26236 47908 26292
rect 47628 25228 47684 25284
rect 47404 25004 47460 25060
rect 47180 24332 47236 24388
rect 47292 23826 47348 23828
rect 47292 23774 47294 23826
rect 47294 23774 47346 23826
rect 47346 23774 47348 23826
rect 47292 23772 47348 23774
rect 47180 23436 47236 23492
rect 47068 22204 47124 22260
rect 46620 21196 46676 21252
rect 46620 20748 46676 20804
rect 46172 19628 46228 19684
rect 46620 20300 46676 20356
rect 46732 20188 46788 20244
rect 46172 19458 46228 19460
rect 46172 19406 46174 19458
rect 46174 19406 46226 19458
rect 46226 19406 46228 19458
rect 46172 19404 46228 19406
rect 46172 18956 46228 19012
rect 46060 18620 46116 18676
rect 46172 17948 46228 18004
rect 46508 19852 46564 19908
rect 46396 18844 46452 18900
rect 45836 16940 45892 16996
rect 45836 16604 45892 16660
rect 45836 15820 45892 15876
rect 46172 16882 46228 16884
rect 46172 16830 46174 16882
rect 46174 16830 46226 16882
rect 46226 16830 46228 16882
rect 46172 16828 46228 16830
rect 46060 15596 46116 15652
rect 45276 14140 45332 14196
rect 45276 13916 45332 13972
rect 45052 9996 45108 10052
rect 44716 9602 44772 9604
rect 44716 9550 44718 9602
rect 44718 9550 44770 9602
rect 44770 9550 44772 9602
rect 44716 9548 44772 9550
rect 45612 14418 45668 14420
rect 45612 14366 45614 14418
rect 45614 14366 45666 14418
rect 45666 14366 45668 14418
rect 45612 14364 45668 14366
rect 46396 15596 46452 15652
rect 46620 19292 46676 19348
rect 47516 23660 47572 23716
rect 47292 23378 47348 23380
rect 47292 23326 47294 23378
rect 47294 23326 47346 23378
rect 47346 23326 47348 23378
rect 47292 23324 47348 23326
rect 47292 22316 47348 22372
rect 47180 21980 47236 22036
rect 47404 21756 47460 21812
rect 47740 24332 47796 24388
rect 48300 28140 48356 28196
rect 49868 33404 49924 33460
rect 50204 34130 50260 34132
rect 50204 34078 50206 34130
rect 50206 34078 50258 34130
rect 50258 34078 50260 34130
rect 50204 34076 50260 34078
rect 50876 35084 50932 35140
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50652 34242 50708 34244
rect 50652 34190 50654 34242
rect 50654 34190 50706 34242
rect 50706 34190 50708 34242
rect 50652 34188 50708 34190
rect 49868 33068 49924 33124
rect 49532 32284 49588 32340
rect 49308 31778 49364 31780
rect 49308 31726 49310 31778
rect 49310 31726 49362 31778
rect 49362 31726 49364 31778
rect 49308 31724 49364 31726
rect 49644 32060 49700 32116
rect 49756 31836 49812 31892
rect 49756 31500 49812 31556
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50428 32620 50484 32676
rect 50764 32786 50820 32788
rect 50764 32734 50766 32786
rect 50766 32734 50818 32786
rect 50818 32734 50820 32786
rect 50764 32732 50820 32734
rect 50204 32562 50260 32564
rect 50204 32510 50206 32562
rect 50206 32510 50258 32562
rect 50258 32510 50260 32562
rect 50204 32508 50260 32510
rect 49980 32284 50036 32340
rect 50764 32284 50820 32340
rect 49980 31948 50036 32004
rect 50204 31666 50260 31668
rect 50204 31614 50206 31666
rect 50206 31614 50258 31666
rect 50258 31614 50260 31666
rect 50204 31612 50260 31614
rect 48748 29426 48804 29428
rect 48748 29374 48750 29426
rect 48750 29374 48802 29426
rect 48802 29374 48804 29426
rect 48748 29372 48804 29374
rect 48636 29148 48692 29204
rect 48524 28924 48580 28980
rect 48860 28812 48916 28868
rect 48636 28476 48692 28532
rect 48972 28140 49028 28196
rect 48412 28028 48468 28084
rect 48076 26684 48132 26740
rect 48076 26290 48132 26292
rect 48076 26238 48078 26290
rect 48078 26238 48130 26290
rect 48130 26238 48132 26290
rect 48076 26236 48132 26238
rect 48300 26012 48356 26068
rect 48076 25506 48132 25508
rect 48076 25454 48078 25506
rect 48078 25454 48130 25506
rect 48130 25454 48132 25506
rect 48076 25452 48132 25454
rect 48188 25282 48244 25284
rect 48188 25230 48190 25282
rect 48190 25230 48242 25282
rect 48242 25230 48244 25282
rect 48188 25228 48244 25230
rect 47964 24892 48020 24948
rect 48076 24780 48132 24836
rect 48076 24444 48132 24500
rect 48860 27468 48916 27524
rect 48412 25282 48468 25284
rect 48412 25230 48414 25282
rect 48414 25230 48466 25282
rect 48466 25230 48468 25282
rect 48412 25228 48468 25230
rect 48524 25116 48580 25172
rect 48300 24444 48356 24500
rect 47964 24108 48020 24164
rect 47852 23436 47908 23492
rect 47740 22764 47796 22820
rect 47628 22316 47684 22372
rect 47740 21698 47796 21700
rect 47740 21646 47742 21698
rect 47742 21646 47794 21698
rect 47794 21646 47796 21698
rect 47740 21644 47796 21646
rect 47516 21586 47572 21588
rect 47516 21534 47518 21586
rect 47518 21534 47570 21586
rect 47570 21534 47572 21586
rect 47516 21532 47572 21534
rect 48636 24780 48692 24836
rect 48748 23996 48804 24052
rect 48188 23938 48244 23940
rect 48188 23886 48190 23938
rect 48190 23886 48242 23938
rect 48242 23886 48244 23938
rect 48188 23884 48244 23886
rect 48412 23772 48468 23828
rect 48188 23266 48244 23268
rect 48188 23214 48190 23266
rect 48190 23214 48242 23266
rect 48242 23214 48244 23266
rect 48188 23212 48244 23214
rect 48188 22652 48244 22708
rect 48412 22258 48468 22260
rect 48412 22206 48414 22258
rect 48414 22206 48466 22258
rect 48466 22206 48468 22258
rect 48412 22204 48468 22206
rect 48188 21980 48244 22036
rect 47964 21308 48020 21364
rect 47404 20690 47460 20692
rect 47404 20638 47406 20690
rect 47406 20638 47458 20690
rect 47458 20638 47460 20690
rect 47404 20636 47460 20638
rect 47628 20412 47684 20468
rect 47404 20076 47460 20132
rect 47180 19852 47236 19908
rect 47516 19516 47572 19572
rect 47404 19404 47460 19460
rect 46956 19292 47012 19348
rect 46620 19068 46676 19124
rect 47628 19122 47684 19124
rect 47628 19070 47630 19122
rect 47630 19070 47682 19122
rect 47682 19070 47684 19122
rect 47628 19068 47684 19070
rect 46956 19010 47012 19012
rect 46956 18958 46958 19010
rect 46958 18958 47010 19010
rect 47010 18958 47012 19010
rect 46956 18956 47012 18958
rect 47516 18844 47572 18900
rect 46956 18620 47012 18676
rect 47180 18396 47236 18452
rect 47180 17778 47236 17780
rect 47180 17726 47182 17778
rect 47182 17726 47234 17778
rect 47234 17726 47236 17778
rect 47180 17724 47236 17726
rect 46844 17500 46900 17556
rect 47068 17164 47124 17220
rect 46732 16940 46788 16996
rect 46508 16156 46564 16212
rect 46620 16268 46676 16324
rect 46620 15986 46676 15988
rect 46620 15934 46622 15986
rect 46622 15934 46674 15986
rect 46674 15934 46676 15986
rect 46620 15932 46676 15934
rect 46956 15426 47012 15428
rect 46956 15374 46958 15426
rect 46958 15374 47010 15426
rect 47010 15374 47012 15426
rect 46956 15372 47012 15374
rect 46844 15260 46900 15316
rect 46172 14476 46228 14532
rect 45836 14140 45892 14196
rect 45388 12348 45444 12404
rect 45388 12178 45444 12180
rect 45388 12126 45390 12178
rect 45390 12126 45442 12178
rect 45442 12126 45444 12178
rect 45388 12124 45444 12126
rect 46060 13020 46116 13076
rect 45724 12402 45780 12404
rect 45724 12350 45726 12402
rect 45726 12350 45778 12402
rect 45778 12350 45780 12402
rect 45724 12348 45780 12350
rect 45388 11004 45444 11060
rect 45276 9548 45332 9604
rect 45388 10610 45444 10612
rect 45388 10558 45390 10610
rect 45390 10558 45442 10610
rect 45442 10558 45444 10610
rect 45388 10556 45444 10558
rect 45276 9100 45332 9156
rect 44828 9042 44884 9044
rect 44828 8990 44830 9042
rect 44830 8990 44882 9042
rect 44882 8990 44884 9042
rect 44828 8988 44884 8990
rect 44716 8652 44772 8708
rect 44828 8370 44884 8372
rect 44828 8318 44830 8370
rect 44830 8318 44882 8370
rect 44882 8318 44884 8370
rect 44828 8316 44884 8318
rect 45164 7868 45220 7924
rect 44492 6578 44548 6580
rect 44492 6526 44494 6578
rect 44494 6526 44546 6578
rect 44546 6526 44548 6578
rect 44492 6524 44548 6526
rect 44604 6412 44660 6468
rect 44716 5404 44772 5460
rect 44268 4284 44324 4340
rect 43932 3388 43988 3444
rect 45388 5404 45444 5460
rect 45500 9996 45556 10052
rect 45612 9884 45668 9940
rect 45612 8764 45668 8820
rect 45948 9660 46004 9716
rect 45612 5292 45668 5348
rect 45612 4956 45668 5012
rect 45724 5068 45780 5124
rect 45276 3836 45332 3892
rect 38108 2716 38164 2772
rect 37884 1484 37940 1540
rect 46172 12684 46228 12740
rect 46172 12460 46228 12516
rect 46732 14140 46788 14196
rect 46508 13970 46564 13972
rect 46508 13918 46510 13970
rect 46510 13918 46562 13970
rect 46562 13918 46564 13970
rect 46508 13916 46564 13918
rect 46396 12962 46452 12964
rect 46396 12910 46398 12962
rect 46398 12910 46450 12962
rect 46450 12910 46452 12962
rect 46396 12908 46452 12910
rect 46508 12460 46564 12516
rect 46172 12012 46228 12068
rect 46396 8764 46452 8820
rect 45948 8258 46004 8260
rect 45948 8206 45950 8258
rect 45950 8206 46002 8258
rect 46002 8206 46004 8258
rect 45948 8204 46004 8206
rect 46620 12236 46676 12292
rect 46956 15036 47012 15092
rect 47180 16882 47236 16884
rect 47180 16830 47182 16882
rect 47182 16830 47234 16882
rect 47234 16830 47236 16882
rect 47180 16828 47236 16830
rect 47180 16604 47236 16660
rect 47404 14812 47460 14868
rect 47068 14252 47124 14308
rect 47852 19404 47908 19460
rect 47852 19068 47908 19124
rect 47628 18284 47684 18340
rect 47740 17724 47796 17780
rect 47740 17164 47796 17220
rect 47964 17442 48020 17444
rect 47964 17390 47966 17442
rect 47966 17390 48018 17442
rect 48018 17390 48020 17442
rect 47964 17388 48020 17390
rect 47628 16604 47684 16660
rect 47628 16098 47684 16100
rect 47628 16046 47630 16098
rect 47630 16046 47682 16098
rect 47682 16046 47684 16098
rect 47628 16044 47684 16046
rect 47852 16380 47908 16436
rect 47740 15372 47796 15428
rect 47628 14306 47684 14308
rect 47628 14254 47630 14306
rect 47630 14254 47682 14306
rect 47682 14254 47684 14306
rect 47628 14252 47684 14254
rect 46956 13468 47012 13524
rect 47068 13580 47124 13636
rect 47292 13020 47348 13076
rect 46956 12460 47012 12516
rect 47068 11676 47124 11732
rect 47180 9548 47236 9604
rect 46508 7644 46564 7700
rect 47628 12908 47684 12964
rect 47852 13356 47908 13412
rect 48300 20300 48356 20356
rect 48412 20748 48468 20804
rect 48636 23714 48692 23716
rect 48636 23662 48638 23714
rect 48638 23662 48690 23714
rect 48690 23662 48692 23714
rect 48636 23660 48692 23662
rect 48636 23378 48692 23380
rect 48636 23326 48638 23378
rect 48638 23326 48690 23378
rect 48690 23326 48692 23378
rect 48636 23324 48692 23326
rect 48636 20578 48692 20580
rect 48636 20526 48638 20578
rect 48638 20526 48690 20578
rect 48690 20526 48692 20578
rect 48636 20524 48692 20526
rect 48636 20188 48692 20244
rect 48300 20018 48356 20020
rect 48300 19966 48302 20018
rect 48302 19966 48354 20018
rect 48354 19966 48356 20018
rect 48300 19964 48356 19966
rect 48300 19404 48356 19460
rect 49980 30492 50036 30548
rect 49532 30268 49588 30324
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 51212 39564 51268 39620
rect 51212 37826 51268 37828
rect 51212 37774 51214 37826
rect 51214 37774 51266 37826
rect 51266 37774 51268 37826
rect 51212 37772 51268 37774
rect 52108 48300 52164 48356
rect 52220 49532 52276 49588
rect 51884 47516 51940 47572
rect 51996 46844 52052 46900
rect 52108 46620 52164 46676
rect 54348 55298 54404 55300
rect 54348 55246 54350 55298
rect 54350 55246 54402 55298
rect 54402 55246 54404 55298
rect 54348 55244 54404 55246
rect 55132 55298 55188 55300
rect 55132 55246 55134 55298
rect 55134 55246 55186 55298
rect 55186 55246 55188 55298
rect 55132 55244 55188 55246
rect 56028 54460 56084 54516
rect 56588 53788 56644 53844
rect 56924 55244 56980 55300
rect 55356 50652 55412 50708
rect 53228 49868 53284 49924
rect 52444 49698 52500 49700
rect 52444 49646 52446 49698
rect 52446 49646 52498 49698
rect 52498 49646 52500 49698
rect 52444 49644 52500 49646
rect 52892 49698 52948 49700
rect 52892 49646 52894 49698
rect 52894 49646 52946 49698
rect 52946 49646 52948 49698
rect 52892 49644 52948 49646
rect 52668 49420 52724 49476
rect 52332 47068 52388 47124
rect 52444 48412 52500 48468
rect 52668 47292 52724 47348
rect 52556 47234 52612 47236
rect 52556 47182 52558 47234
rect 52558 47182 52610 47234
rect 52610 47182 52612 47234
rect 52556 47180 52612 47182
rect 52220 46396 52276 46452
rect 52108 45666 52164 45668
rect 52108 45614 52110 45666
rect 52110 45614 52162 45666
rect 52162 45614 52164 45666
rect 52108 45612 52164 45614
rect 51660 43820 51716 43876
rect 51548 43596 51604 43652
rect 51660 42588 51716 42644
rect 51548 42028 51604 42084
rect 51548 41858 51604 41860
rect 51548 41806 51550 41858
rect 51550 41806 51602 41858
rect 51602 41806 51604 41858
rect 51548 41804 51604 41806
rect 51884 43820 51940 43876
rect 51996 43708 52052 43764
rect 52444 46674 52500 46676
rect 52444 46622 52446 46674
rect 52446 46622 52498 46674
rect 52498 46622 52500 46674
rect 52444 46620 52500 46622
rect 53452 48802 53508 48804
rect 53452 48750 53454 48802
rect 53454 48750 53506 48802
rect 53506 48750 53508 48802
rect 53452 48748 53508 48750
rect 53228 47740 53284 47796
rect 53340 48300 53396 48356
rect 52892 46844 52948 46900
rect 52556 45778 52612 45780
rect 52556 45726 52558 45778
rect 52558 45726 52610 45778
rect 52610 45726 52612 45778
rect 52556 45724 52612 45726
rect 52332 44940 52388 44996
rect 52220 43372 52276 43428
rect 52108 43148 52164 43204
rect 51996 42028 52052 42084
rect 52220 41804 52276 41860
rect 51436 40348 51492 40404
rect 51548 40908 51604 40964
rect 51436 39340 51492 39396
rect 51436 38892 51492 38948
rect 51324 37660 51380 37716
rect 52108 41020 52164 41076
rect 51772 40962 51828 40964
rect 51772 40910 51774 40962
rect 51774 40910 51826 40962
rect 51826 40910 51828 40962
rect 51772 40908 51828 40910
rect 51884 40626 51940 40628
rect 51884 40574 51886 40626
rect 51886 40574 51938 40626
rect 51938 40574 51940 40626
rect 51884 40572 51940 40574
rect 52444 41020 52500 41076
rect 52668 44098 52724 44100
rect 52668 44046 52670 44098
rect 52670 44046 52722 44098
rect 52722 44046 52724 44098
rect 52668 44044 52724 44046
rect 53452 48242 53508 48244
rect 53452 48190 53454 48242
rect 53454 48190 53506 48242
rect 53506 48190 53508 48242
rect 53452 48188 53508 48190
rect 53340 47628 53396 47684
rect 52892 46674 52948 46676
rect 52892 46622 52894 46674
rect 52894 46622 52946 46674
rect 52946 46622 52948 46674
rect 52892 46620 52948 46622
rect 54348 48802 54404 48804
rect 54348 48750 54350 48802
rect 54350 48750 54402 48802
rect 54402 48750 54404 48802
rect 54348 48748 54404 48750
rect 53900 48412 53956 48468
rect 54572 48188 54628 48244
rect 55020 48188 55076 48244
rect 55468 48748 55524 48804
rect 54684 48076 54740 48132
rect 54236 47740 54292 47796
rect 53676 47516 53732 47572
rect 53564 47458 53620 47460
rect 53564 47406 53566 47458
rect 53566 47406 53618 47458
rect 53618 47406 53620 47458
rect 54012 47458 54068 47460
rect 53564 47404 53620 47406
rect 53452 47346 53508 47348
rect 53452 47294 53454 47346
rect 53454 47294 53506 47346
rect 53506 47294 53508 47346
rect 53452 47292 53508 47294
rect 54012 47406 54014 47458
rect 54014 47406 54066 47458
rect 54066 47406 54068 47458
rect 54012 47404 54068 47406
rect 53228 45724 53284 45780
rect 53452 45778 53508 45780
rect 53452 45726 53454 45778
rect 53454 45726 53506 45778
rect 53506 45726 53508 45778
rect 53452 45724 53508 45726
rect 53452 45500 53508 45556
rect 53116 44604 53172 44660
rect 53788 46620 53844 46676
rect 53900 46956 53956 47012
rect 53900 45500 53956 45556
rect 54348 46956 54404 47012
rect 54460 47404 54516 47460
rect 54572 47180 54628 47236
rect 54012 45388 54068 45444
rect 53788 45276 53844 45332
rect 54012 45218 54068 45220
rect 54012 45166 54014 45218
rect 54014 45166 54066 45218
rect 54066 45166 54068 45218
rect 54012 45164 54068 45166
rect 53676 44492 53732 44548
rect 53340 43484 53396 43540
rect 53228 43426 53284 43428
rect 53228 43374 53230 43426
rect 53230 43374 53282 43426
rect 53282 43374 53284 43426
rect 53228 43372 53284 43374
rect 53116 42194 53172 42196
rect 53116 42142 53118 42194
rect 53118 42142 53170 42194
rect 53170 42142 53172 42194
rect 53116 42140 53172 42142
rect 52332 40684 52388 40740
rect 52668 40908 52724 40964
rect 52220 40460 52276 40516
rect 52556 40572 52612 40628
rect 52108 40348 52164 40404
rect 52444 40236 52500 40292
rect 52108 39564 52164 39620
rect 52108 39004 52164 39060
rect 51996 38946 52052 38948
rect 51996 38894 51998 38946
rect 51998 38894 52050 38946
rect 52050 38894 52052 38946
rect 51996 38892 52052 38894
rect 51212 37154 51268 37156
rect 51212 37102 51214 37154
rect 51214 37102 51266 37154
rect 51266 37102 51268 37154
rect 51212 37100 51268 37102
rect 51660 35922 51716 35924
rect 51660 35870 51662 35922
rect 51662 35870 51714 35922
rect 51714 35870 51716 35922
rect 51660 35868 51716 35870
rect 51548 35810 51604 35812
rect 51548 35758 51550 35810
rect 51550 35758 51602 35810
rect 51602 35758 51604 35810
rect 51548 35756 51604 35758
rect 51324 34748 51380 34804
rect 50988 34188 51044 34244
rect 51884 37660 51940 37716
rect 51884 35810 51940 35812
rect 51884 35758 51886 35810
rect 51886 35758 51938 35810
rect 51938 35758 51940 35810
rect 51884 35756 51940 35758
rect 52108 37212 52164 37268
rect 52556 40124 52612 40180
rect 52444 40012 52500 40068
rect 52332 39116 52388 39172
rect 52332 38050 52388 38052
rect 52332 37998 52334 38050
rect 52334 37998 52386 38050
rect 52386 37998 52388 38050
rect 52332 37996 52388 37998
rect 52332 37324 52388 37380
rect 52220 36594 52276 36596
rect 52220 36542 52222 36594
rect 52222 36542 52274 36594
rect 52274 36542 52276 36594
rect 52220 36540 52276 36542
rect 52108 36482 52164 36484
rect 52108 36430 52110 36482
rect 52110 36430 52162 36482
rect 52162 36430 52164 36482
rect 52108 36428 52164 36430
rect 52220 35532 52276 35588
rect 51996 35084 52052 35140
rect 52108 35308 52164 35364
rect 51996 34914 52052 34916
rect 51996 34862 51998 34914
rect 51998 34862 52050 34914
rect 52050 34862 52052 34914
rect 51996 34860 52052 34862
rect 51996 34412 52052 34468
rect 51884 34188 51940 34244
rect 51436 33570 51492 33572
rect 51436 33518 51438 33570
rect 51438 33518 51490 33570
rect 51490 33518 51492 33570
rect 51436 33516 51492 33518
rect 51548 33458 51604 33460
rect 51548 33406 51550 33458
rect 51550 33406 51602 33458
rect 51602 33406 51604 33458
rect 51548 33404 51604 33406
rect 50988 33346 51044 33348
rect 50988 33294 50990 33346
rect 50990 33294 51042 33346
rect 51042 33294 51044 33346
rect 50988 33292 51044 33294
rect 50988 33068 51044 33124
rect 51660 32732 51716 32788
rect 51772 32620 51828 32676
rect 50988 31948 51044 32004
rect 51436 31836 51492 31892
rect 50204 30380 50260 30436
rect 50428 31164 50484 31220
rect 50428 30268 50484 30324
rect 50540 31052 50596 31108
rect 50876 30940 50932 30996
rect 51548 31164 51604 31220
rect 50876 30770 50932 30772
rect 50876 30718 50878 30770
rect 50878 30718 50930 30770
rect 50930 30718 50932 30770
rect 50876 30716 50932 30718
rect 51660 30716 51716 30772
rect 50204 29708 50260 29764
rect 49980 29484 50036 29540
rect 49420 26962 49476 26964
rect 49420 26910 49422 26962
rect 49422 26910 49474 26962
rect 49474 26910 49476 26962
rect 49420 26908 49476 26910
rect 49196 26348 49252 26404
rect 49756 29426 49812 29428
rect 49756 29374 49758 29426
rect 49758 29374 49810 29426
rect 49810 29374 49812 29426
rect 49756 29372 49812 29374
rect 50204 29372 50260 29428
rect 50092 28700 50148 28756
rect 49980 28588 50036 28644
rect 49868 28252 49924 28308
rect 49868 28082 49924 28084
rect 49868 28030 49870 28082
rect 49870 28030 49922 28082
rect 49922 28030 49924 28082
rect 49868 28028 49924 28030
rect 49644 27858 49700 27860
rect 49644 27806 49646 27858
rect 49646 27806 49698 27858
rect 49698 27806 49700 27858
rect 49644 27804 49700 27806
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50876 29538 50932 29540
rect 50876 29486 50878 29538
rect 50878 29486 50930 29538
rect 50930 29486 50932 29538
rect 50876 29484 50932 29486
rect 51100 30044 51156 30100
rect 50988 28924 51044 28980
rect 50652 28588 50708 28644
rect 50876 28418 50932 28420
rect 50876 28366 50878 28418
rect 50878 28366 50930 28418
rect 50930 28366 50932 28418
rect 50876 28364 50932 28366
rect 50092 28028 50148 28084
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 51212 29202 51268 29204
rect 51212 29150 51214 29202
rect 51214 29150 51266 29202
rect 51266 29150 51268 29202
rect 51212 29148 51268 29150
rect 51772 29484 51828 29540
rect 51324 29260 51380 29316
rect 51100 28476 51156 28532
rect 51212 28140 51268 28196
rect 50204 27916 50260 27972
rect 50316 27804 50372 27860
rect 49196 25788 49252 25844
rect 48972 25564 49028 25620
rect 49084 25394 49140 25396
rect 49084 25342 49086 25394
rect 49086 25342 49138 25394
rect 49138 25342 49140 25394
rect 49084 25340 49140 25342
rect 48972 25004 49028 25060
rect 49756 25900 49812 25956
rect 49868 26236 49924 26292
rect 50428 26908 50484 26964
rect 50092 26850 50148 26852
rect 50092 26798 50094 26850
rect 50094 26798 50146 26850
rect 50146 26798 50148 26850
rect 50092 26796 50148 26798
rect 50092 26402 50148 26404
rect 50092 26350 50094 26402
rect 50094 26350 50146 26402
rect 50146 26350 50148 26402
rect 50092 26348 50148 26350
rect 50652 27468 50708 27524
rect 50764 27916 50820 27972
rect 50204 26236 50260 26292
rect 50204 25788 50260 25844
rect 49756 25116 49812 25172
rect 49868 25228 49924 25284
rect 49644 24668 49700 24724
rect 49308 24162 49364 24164
rect 49308 24110 49310 24162
rect 49310 24110 49362 24162
rect 49362 24110 49364 24162
rect 49308 24108 49364 24110
rect 49420 23826 49476 23828
rect 49420 23774 49422 23826
rect 49422 23774 49474 23826
rect 49474 23774 49476 23826
rect 49420 23772 49476 23774
rect 49308 23436 49364 23492
rect 49532 23492 49588 23548
rect 50092 23492 50148 23548
rect 50092 23324 50148 23380
rect 49756 23266 49812 23268
rect 49756 23214 49758 23266
rect 49758 23214 49810 23266
rect 49810 23214 49812 23266
rect 49756 23212 49812 23214
rect 49084 22764 49140 22820
rect 48972 22370 49028 22372
rect 48972 22318 48974 22370
rect 48974 22318 49026 22370
rect 49026 22318 49028 22370
rect 48972 22316 49028 22318
rect 49084 20412 49140 20468
rect 49084 20076 49140 20132
rect 48860 20018 48916 20020
rect 48860 19966 48862 20018
rect 48862 19966 48914 20018
rect 48914 19966 48916 20018
rect 48860 19964 48916 19966
rect 48300 18396 48356 18452
rect 48748 19234 48804 19236
rect 48748 19182 48750 19234
rect 48750 19182 48802 19234
rect 48802 19182 48804 19234
rect 48748 19180 48804 19182
rect 48636 18732 48692 18788
rect 48412 18226 48468 18228
rect 48412 18174 48414 18226
rect 48414 18174 48466 18226
rect 48466 18174 48468 18226
rect 48412 18172 48468 18174
rect 48300 17612 48356 17668
rect 48412 17500 48468 17556
rect 48188 16882 48244 16884
rect 48188 16830 48190 16882
rect 48190 16830 48242 16882
rect 48242 16830 48244 16882
rect 48188 16828 48244 16830
rect 48076 16716 48132 16772
rect 48300 16210 48356 16212
rect 48300 16158 48302 16210
rect 48302 16158 48354 16210
rect 48354 16158 48356 16210
rect 48300 16156 48356 16158
rect 48972 19346 49028 19348
rect 48972 19294 48974 19346
rect 48974 19294 49026 19346
rect 49026 19294 49028 19346
rect 48972 19292 49028 19294
rect 48748 17778 48804 17780
rect 48748 17726 48750 17778
rect 48750 17726 48802 17778
rect 48802 17726 48804 17778
rect 48748 17724 48804 17726
rect 49196 17948 49252 18004
rect 50092 22988 50148 23044
rect 49644 22930 49700 22932
rect 49644 22878 49646 22930
rect 49646 22878 49698 22930
rect 49698 22878 49700 22930
rect 49644 22876 49700 22878
rect 49980 22764 50036 22820
rect 49420 21868 49476 21924
rect 49644 21756 49700 21812
rect 49756 22146 49812 22148
rect 49756 22094 49758 22146
rect 49758 22094 49810 22146
rect 49810 22094 49812 22146
rect 49756 22092 49812 22094
rect 49644 21308 49700 21364
rect 49532 19740 49588 19796
rect 49532 19068 49588 19124
rect 49532 18396 49588 18452
rect 49308 17388 49364 17444
rect 49420 18284 49476 18340
rect 49084 17052 49140 17108
rect 48188 15426 48244 15428
rect 48188 15374 48190 15426
rect 48190 15374 48242 15426
rect 48242 15374 48244 15426
rect 48188 15372 48244 15374
rect 48524 15148 48580 15204
rect 48412 14700 48468 14756
rect 48188 14642 48244 14644
rect 48188 14590 48190 14642
rect 48190 14590 48242 14642
rect 48242 14590 48244 14642
rect 48188 14588 48244 14590
rect 48188 14252 48244 14308
rect 49308 16156 49364 16212
rect 48972 15874 49028 15876
rect 48972 15822 48974 15874
rect 48974 15822 49026 15874
rect 49026 15822 49028 15874
rect 48972 15820 49028 15822
rect 48748 15148 48804 15204
rect 48748 14700 48804 14756
rect 48636 14252 48692 14308
rect 48972 14476 49028 14532
rect 48188 13468 48244 13524
rect 47964 12962 48020 12964
rect 47964 12910 47966 12962
rect 47966 12910 48018 12962
rect 48018 12910 48020 12962
rect 47964 12908 48020 12910
rect 47740 12348 47796 12404
rect 47852 12236 47908 12292
rect 47740 12066 47796 12068
rect 47740 12014 47742 12066
rect 47742 12014 47794 12066
rect 47794 12014 47796 12066
rect 47740 12012 47796 12014
rect 47628 11506 47684 11508
rect 47628 11454 47630 11506
rect 47630 11454 47682 11506
rect 47682 11454 47684 11506
rect 47628 11452 47684 11454
rect 47740 11004 47796 11060
rect 47628 10892 47684 10948
rect 47292 7698 47348 7700
rect 47292 7646 47294 7698
rect 47294 7646 47346 7698
rect 47346 7646 47348 7698
rect 47292 7644 47348 7646
rect 46620 7420 46676 7476
rect 45948 6690 46004 6692
rect 45948 6638 45950 6690
rect 45950 6638 46002 6690
rect 46002 6638 46004 6690
rect 45948 6636 46004 6638
rect 46956 7532 47012 7588
rect 47068 6636 47124 6692
rect 45948 4508 46004 4564
rect 46732 4956 46788 5012
rect 46172 3836 46228 3892
rect 46732 3666 46788 3668
rect 46732 3614 46734 3666
rect 46734 3614 46786 3666
rect 46786 3614 46788 3666
rect 46732 3612 46788 3614
rect 48076 11676 48132 11732
rect 47964 9884 48020 9940
rect 48076 9660 48132 9716
rect 48636 12908 48692 12964
rect 48860 13244 48916 13300
rect 49308 15596 49364 15652
rect 49308 15372 49364 15428
rect 49756 21196 49812 21252
rect 49980 20578 50036 20580
rect 49980 20526 49982 20578
rect 49982 20526 50034 20578
rect 50034 20526 50036 20578
rect 49980 20524 50036 20526
rect 49756 20076 49812 20132
rect 49868 19234 49924 19236
rect 49868 19182 49870 19234
rect 49870 19182 49922 19234
rect 49922 19182 49924 19234
rect 49868 19180 49924 19182
rect 49644 17778 49700 17780
rect 49644 17726 49646 17778
rect 49646 17726 49698 17778
rect 49698 17726 49700 17778
rect 49644 17724 49700 17726
rect 49644 16994 49700 16996
rect 49644 16942 49646 16994
rect 49646 16942 49698 16994
rect 49698 16942 49700 16994
rect 49644 16940 49700 16942
rect 49980 18284 50036 18340
rect 49868 17612 49924 17668
rect 49980 17500 50036 17556
rect 49532 16380 49588 16436
rect 49644 16098 49700 16100
rect 49644 16046 49646 16098
rect 49646 16046 49698 16098
rect 49698 16046 49700 16098
rect 49644 16044 49700 16046
rect 49532 14306 49588 14308
rect 49532 14254 49534 14306
rect 49534 14254 49586 14306
rect 49586 14254 49588 14306
rect 49532 14252 49588 14254
rect 49420 14140 49476 14196
rect 49084 13804 49140 13860
rect 49644 13804 49700 13860
rect 48972 13074 49028 13076
rect 48972 13022 48974 13074
rect 48974 13022 49026 13074
rect 49026 13022 49028 13074
rect 48972 13020 49028 13022
rect 48748 12796 48804 12852
rect 48748 12460 48804 12516
rect 48636 11676 48692 11732
rect 48524 10386 48580 10388
rect 48524 10334 48526 10386
rect 48526 10334 48578 10386
rect 48578 10334 48580 10386
rect 48524 10332 48580 10334
rect 48860 11282 48916 11284
rect 48860 11230 48862 11282
rect 48862 11230 48914 11282
rect 48914 11230 48916 11282
rect 48860 11228 48916 11230
rect 50316 24668 50372 24724
rect 50652 26796 50708 26852
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 51212 27020 51268 27076
rect 51660 28588 51716 28644
rect 51324 26908 51380 26964
rect 51100 26572 51156 26628
rect 50764 26514 50820 26516
rect 50764 26462 50766 26514
rect 50766 26462 50818 26514
rect 50818 26462 50820 26514
rect 50764 26460 50820 26462
rect 51100 26236 51156 26292
rect 51324 26684 51380 26740
rect 51212 26012 51268 26068
rect 51212 25506 51268 25508
rect 51212 25454 51214 25506
rect 51214 25454 51266 25506
rect 51266 25454 51268 25506
rect 51212 25452 51268 25454
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 51772 28364 51828 28420
rect 52892 40684 52948 40740
rect 52444 36652 52500 36708
rect 52556 38668 52612 38724
rect 52444 36370 52500 36372
rect 52444 36318 52446 36370
rect 52446 36318 52498 36370
rect 52498 36318 52500 36370
rect 52444 36316 52500 36318
rect 52780 38274 52836 38276
rect 52780 38222 52782 38274
rect 52782 38222 52834 38274
rect 52834 38222 52836 38274
rect 52780 38220 52836 38222
rect 52892 37996 52948 38052
rect 52780 37660 52836 37716
rect 53116 40460 53172 40516
rect 52668 36540 52724 36596
rect 52668 35922 52724 35924
rect 52668 35870 52670 35922
rect 52670 35870 52722 35922
rect 52722 35870 52724 35922
rect 52668 35868 52724 35870
rect 53228 40402 53284 40404
rect 53228 40350 53230 40402
rect 53230 40350 53282 40402
rect 53282 40350 53284 40402
rect 53228 40348 53284 40350
rect 53676 44156 53732 44212
rect 53452 40012 53508 40068
rect 53564 43484 53620 43540
rect 53452 39004 53508 39060
rect 53676 43148 53732 43204
rect 53900 43820 53956 43876
rect 54012 44268 54068 44324
rect 53900 43260 53956 43316
rect 54460 45388 54516 45444
rect 54460 44828 54516 44884
rect 54908 47346 54964 47348
rect 54908 47294 54910 47346
rect 54910 47294 54962 47346
rect 54962 47294 54964 47346
rect 54908 47292 54964 47294
rect 54012 42700 54068 42756
rect 54796 45666 54852 45668
rect 54796 45614 54798 45666
rect 54798 45614 54850 45666
rect 54850 45614 54852 45666
rect 54796 45612 54852 45614
rect 54684 44156 54740 44212
rect 55244 47628 55300 47684
rect 55356 47180 55412 47236
rect 56028 48412 56084 48468
rect 55468 46732 55524 46788
rect 55356 46562 55412 46564
rect 55356 46510 55358 46562
rect 55358 46510 55410 46562
rect 55410 46510 55412 46562
rect 55356 46508 55412 46510
rect 54908 45276 54964 45332
rect 54908 44380 54964 44436
rect 54348 43036 54404 43092
rect 53788 40012 53844 40068
rect 53900 39900 53956 39956
rect 53788 39394 53844 39396
rect 53788 39342 53790 39394
rect 53790 39342 53842 39394
rect 53842 39342 53844 39394
rect 53788 39340 53844 39342
rect 53676 39116 53732 39172
rect 53676 38834 53732 38836
rect 53676 38782 53678 38834
rect 53678 38782 53730 38834
rect 53730 38782 53732 38834
rect 53676 38780 53732 38782
rect 53340 38332 53396 38388
rect 53004 37266 53060 37268
rect 53004 37214 53006 37266
rect 53006 37214 53058 37266
rect 53058 37214 53060 37266
rect 53004 37212 53060 37214
rect 53228 37324 53284 37380
rect 52556 35196 52612 35252
rect 52332 34300 52388 34356
rect 52892 34636 52948 34692
rect 53004 36876 53060 36932
rect 52780 34242 52836 34244
rect 52780 34190 52782 34242
rect 52782 34190 52834 34242
rect 52834 34190 52836 34242
rect 52780 34188 52836 34190
rect 52892 33516 52948 33572
rect 52332 33122 52388 33124
rect 52332 33070 52334 33122
rect 52334 33070 52386 33122
rect 52386 33070 52388 33122
rect 52332 33068 52388 33070
rect 52332 32844 52388 32900
rect 52332 32396 52388 32452
rect 52220 31724 52276 31780
rect 51996 31276 52052 31332
rect 52444 31948 52500 32004
rect 52668 33122 52724 33124
rect 52668 33070 52670 33122
rect 52670 33070 52722 33122
rect 52722 33070 52724 33122
rect 52668 33068 52724 33070
rect 51996 30156 52052 30212
rect 52332 31106 52388 31108
rect 52332 31054 52334 31106
rect 52334 31054 52386 31106
rect 52386 31054 52388 31106
rect 52332 31052 52388 31054
rect 51996 28588 52052 28644
rect 52668 31778 52724 31780
rect 52668 31726 52670 31778
rect 52670 31726 52722 31778
rect 52722 31726 52724 31778
rect 52668 31724 52724 31726
rect 53116 34076 53172 34132
rect 53116 33068 53172 33124
rect 53004 31276 53060 31332
rect 53116 31218 53172 31220
rect 53116 31166 53118 31218
rect 53118 31166 53170 31218
rect 53170 31166 53172 31218
rect 53116 31164 53172 31166
rect 52556 30434 52612 30436
rect 52556 30382 52558 30434
rect 52558 30382 52610 30434
rect 52610 30382 52612 30434
rect 52556 30380 52612 30382
rect 52444 30044 52500 30100
rect 52332 29708 52388 29764
rect 52444 29260 52500 29316
rect 51660 26348 51716 26404
rect 51996 28252 52052 28308
rect 51660 26178 51716 26180
rect 51660 26126 51662 26178
rect 51662 26126 51714 26178
rect 51714 26126 51716 26178
rect 51660 26124 51716 26126
rect 51884 27970 51940 27972
rect 51884 27918 51886 27970
rect 51886 27918 51938 27970
rect 51938 27918 51940 27970
rect 51884 27916 51940 27918
rect 51884 27298 51940 27300
rect 51884 27246 51886 27298
rect 51886 27246 51938 27298
rect 51938 27246 51940 27298
rect 51884 27244 51940 27246
rect 52108 27580 52164 27636
rect 52108 27020 52164 27076
rect 51996 26124 52052 26180
rect 51884 25564 51940 25620
rect 51324 25228 51380 25284
rect 51660 25228 51716 25284
rect 51100 24722 51156 24724
rect 51100 24670 51102 24722
rect 51102 24670 51154 24722
rect 51154 24670 51156 24722
rect 51100 24668 51156 24670
rect 50764 24556 50820 24612
rect 50316 24332 50372 24388
rect 50876 23996 50932 24052
rect 50540 23826 50596 23828
rect 50540 23774 50542 23826
rect 50542 23774 50594 23826
rect 50594 23774 50596 23826
rect 50540 23772 50596 23774
rect 50316 22316 50372 22372
rect 50428 23660 50484 23716
rect 50652 23714 50708 23716
rect 50652 23662 50654 23714
rect 50654 23662 50706 23714
rect 50706 23662 50708 23714
rect 50652 23660 50708 23662
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50540 22988 50596 23044
rect 50652 22428 50708 22484
rect 50540 22204 50596 22260
rect 50764 22258 50820 22260
rect 50764 22206 50766 22258
rect 50766 22206 50818 22258
rect 50818 22206 50820 22258
rect 50764 22204 50820 22206
rect 50428 22092 50484 22148
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 51100 23324 51156 23380
rect 50540 21810 50596 21812
rect 50540 21758 50542 21810
rect 50542 21758 50594 21810
rect 50594 21758 50596 21810
rect 50540 21756 50596 21758
rect 50988 21980 51044 22036
rect 50988 21756 51044 21812
rect 50540 21586 50596 21588
rect 50540 21534 50542 21586
rect 50542 21534 50594 21586
rect 50594 21534 50596 21586
rect 50540 21532 50596 21534
rect 50876 21586 50932 21588
rect 50876 21534 50878 21586
rect 50878 21534 50930 21586
rect 50930 21534 50932 21586
rect 50876 21532 50932 21534
rect 51548 23996 51604 24052
rect 51548 23436 51604 23492
rect 51212 22540 51268 22596
rect 51324 23100 51380 23156
rect 51548 22540 51604 22596
rect 51100 21420 51156 21476
rect 51212 22316 51268 22372
rect 50764 20972 50820 21028
rect 50988 21196 51044 21252
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50316 20018 50372 20020
rect 50316 19966 50318 20018
rect 50318 19966 50370 20018
rect 50370 19966 50372 20018
rect 50316 19964 50372 19966
rect 50764 19964 50820 20020
rect 50652 19794 50708 19796
rect 50652 19742 50654 19794
rect 50654 19742 50706 19794
rect 50706 19742 50708 19794
rect 50652 19740 50708 19742
rect 50540 19180 50596 19236
rect 50204 19068 50260 19124
rect 50652 19068 50708 19124
rect 50988 19180 51044 19236
rect 50204 18844 50260 18900
rect 50556 18842 50612 18844
rect 50316 18732 50372 18788
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50876 18508 50932 18564
rect 50764 18338 50820 18340
rect 50764 18286 50766 18338
rect 50766 18286 50818 18338
rect 50818 18286 50820 18338
rect 50764 18284 50820 18286
rect 51436 21980 51492 22036
rect 51884 23042 51940 23044
rect 51884 22990 51886 23042
rect 51886 22990 51938 23042
rect 51938 22990 51940 23042
rect 51884 22988 51940 22990
rect 52332 27186 52388 27188
rect 52332 27134 52334 27186
rect 52334 27134 52386 27186
rect 52386 27134 52388 27186
rect 52332 27132 52388 27134
rect 52332 25618 52388 25620
rect 52332 25566 52334 25618
rect 52334 25566 52386 25618
rect 52386 25566 52388 25618
rect 52332 25564 52388 25566
rect 52444 25228 52500 25284
rect 52332 25004 52388 25060
rect 52332 24332 52388 24388
rect 51996 22428 52052 22484
rect 52108 22652 52164 22708
rect 51660 21980 51716 22036
rect 51772 21756 51828 21812
rect 52444 23266 52500 23268
rect 52444 23214 52446 23266
rect 52446 23214 52498 23266
rect 52498 23214 52500 23266
rect 52444 23212 52500 23214
rect 52332 22370 52388 22372
rect 52332 22318 52334 22370
rect 52334 22318 52386 22370
rect 52386 22318 52388 22370
rect 52332 22316 52388 22318
rect 51996 21980 52052 22036
rect 52444 22204 52500 22260
rect 51436 20972 51492 21028
rect 51772 21308 51828 21364
rect 51548 20860 51604 20916
rect 51660 20748 51716 20804
rect 51884 20188 51940 20244
rect 51772 20076 51828 20132
rect 51884 20018 51940 20020
rect 51884 19966 51886 20018
rect 51886 19966 51938 20018
rect 51938 19966 51940 20018
rect 51884 19964 51940 19966
rect 51548 19628 51604 19684
rect 51436 19234 51492 19236
rect 51436 19182 51438 19234
rect 51438 19182 51490 19234
rect 51490 19182 51492 19234
rect 51436 19180 51492 19182
rect 51548 19068 51604 19124
rect 51324 18732 51380 18788
rect 51324 18508 51380 18564
rect 50204 17276 50260 17332
rect 50316 17612 50372 17668
rect 50428 17442 50484 17444
rect 50428 17390 50430 17442
rect 50430 17390 50482 17442
rect 50482 17390 50484 17442
rect 50428 17388 50484 17390
rect 50876 17388 50932 17444
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50540 16882 50596 16884
rect 50540 16830 50542 16882
rect 50542 16830 50594 16882
rect 50594 16830 50596 16882
rect 50540 16828 50596 16830
rect 50764 15932 50820 15988
rect 50428 15820 50484 15876
rect 50316 15708 50372 15764
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50428 15372 50484 15428
rect 50316 15036 50372 15092
rect 50316 14642 50372 14644
rect 50316 14590 50318 14642
rect 50318 14590 50370 14642
rect 50370 14590 50372 14642
rect 50316 14588 50372 14590
rect 50652 14306 50708 14308
rect 50652 14254 50654 14306
rect 50654 14254 50706 14306
rect 50706 14254 50708 14306
rect 50652 14252 50708 14254
rect 50876 15202 50932 15204
rect 50876 15150 50878 15202
rect 50878 15150 50930 15202
rect 50930 15150 50932 15202
rect 50876 15148 50932 15150
rect 50988 14476 51044 14532
rect 51548 16994 51604 16996
rect 51548 16942 51550 16994
rect 51550 16942 51602 16994
rect 51602 16942 51604 16994
rect 51548 16940 51604 16942
rect 51212 16098 51268 16100
rect 51212 16046 51214 16098
rect 51214 16046 51266 16098
rect 51266 16046 51268 16098
rect 51212 16044 51268 16046
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 49868 13580 49924 13636
rect 49196 12796 49252 12852
rect 49644 12850 49700 12852
rect 49644 12798 49646 12850
rect 49646 12798 49698 12850
rect 49698 12798 49700 12850
rect 49644 12796 49700 12798
rect 49756 12572 49812 12628
rect 49644 12460 49700 12516
rect 49420 11900 49476 11956
rect 49420 11506 49476 11508
rect 49420 11454 49422 11506
rect 49422 11454 49474 11506
rect 49474 11454 49476 11506
rect 49420 11452 49476 11454
rect 49868 12290 49924 12292
rect 49868 12238 49870 12290
rect 49870 12238 49922 12290
rect 49922 12238 49924 12290
rect 49868 12236 49924 12238
rect 49868 11564 49924 11620
rect 48636 10108 48692 10164
rect 48300 9884 48356 9940
rect 48300 9266 48356 9268
rect 48300 9214 48302 9266
rect 48302 9214 48354 9266
rect 48354 9214 48356 9266
rect 48300 9212 48356 9214
rect 49084 10050 49140 10052
rect 49084 9998 49086 10050
rect 49086 9998 49138 10050
rect 49138 9998 49140 10050
rect 49084 9996 49140 9998
rect 49532 9996 49588 10052
rect 49420 9938 49476 9940
rect 49420 9886 49422 9938
rect 49422 9886 49474 9938
rect 49474 9886 49476 9938
rect 49420 9884 49476 9886
rect 50092 11676 50148 11732
rect 50204 13468 50260 13524
rect 50428 13356 50484 13412
rect 50316 12460 50372 12516
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 50876 12402 50932 12404
rect 50876 12350 50878 12402
rect 50878 12350 50930 12402
rect 50930 12350 50932 12402
rect 50876 12348 50932 12350
rect 50540 11900 50596 11956
rect 50764 11788 50820 11844
rect 50540 11676 50596 11732
rect 49980 10556 50036 10612
rect 50652 11564 50708 11620
rect 47628 6076 47684 6132
rect 48188 6860 48244 6916
rect 48188 5740 48244 5796
rect 49420 8034 49476 8036
rect 49420 7982 49422 8034
rect 49422 7982 49474 8034
rect 49474 7982 49476 8034
rect 49420 7980 49476 7982
rect 49532 7698 49588 7700
rect 49532 7646 49534 7698
rect 49534 7646 49586 7698
rect 49586 7646 49588 7698
rect 49532 7644 49588 7646
rect 49980 8258 50036 8260
rect 49980 8206 49982 8258
rect 49982 8206 50034 8258
rect 50034 8206 50036 8258
rect 49980 8204 50036 8206
rect 50316 11228 50372 11284
rect 50204 11170 50260 11172
rect 50204 11118 50206 11170
rect 50206 11118 50258 11170
rect 50258 11118 50260 11170
rect 50204 11116 50260 11118
rect 50092 7532 50148 7588
rect 50204 10668 50260 10724
rect 49868 7308 49924 7364
rect 49420 7196 49476 7252
rect 49084 6636 49140 6692
rect 50652 11170 50708 11172
rect 50652 11118 50654 11170
rect 50654 11118 50706 11170
rect 50706 11118 50708 11170
rect 50652 11116 50708 11118
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 50988 11452 51044 11508
rect 51100 13468 51156 13524
rect 50988 10892 51044 10948
rect 50876 10108 50932 10164
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 50428 8930 50484 8932
rect 50428 8878 50430 8930
rect 50430 8878 50482 8930
rect 50482 8878 50484 8930
rect 50428 8876 50484 8878
rect 50876 8428 50932 8484
rect 50316 7698 50372 7700
rect 50316 7646 50318 7698
rect 50318 7646 50370 7698
rect 50370 7646 50372 7698
rect 50316 7644 50372 7646
rect 48524 6524 48580 6580
rect 49420 6578 49476 6580
rect 49420 6526 49422 6578
rect 49422 6526 49474 6578
rect 49474 6526 49476 6578
rect 49420 6524 49476 6526
rect 49868 6578 49924 6580
rect 49868 6526 49870 6578
rect 49870 6526 49922 6578
rect 49922 6526 49924 6578
rect 49868 6524 49924 6526
rect 48524 6130 48580 6132
rect 48524 6078 48526 6130
rect 48526 6078 48578 6130
rect 48578 6078 48580 6130
rect 48524 6076 48580 6078
rect 48972 6076 49028 6132
rect 47292 5292 47348 5348
rect 47740 4844 47796 4900
rect 47516 4732 47572 4788
rect 49868 6076 49924 6132
rect 49980 5964 50036 6020
rect 49084 5628 49140 5684
rect 48076 4562 48132 4564
rect 48076 4510 48078 4562
rect 48078 4510 48130 4562
rect 48130 4510 48132 4562
rect 48076 4508 48132 4510
rect 48524 4898 48580 4900
rect 48524 4846 48526 4898
rect 48526 4846 48578 4898
rect 48578 4846 48580 4898
rect 48524 4844 48580 4846
rect 48524 3836 48580 3892
rect 48748 3724 48804 3780
rect 48860 3666 48916 3668
rect 48860 3614 48862 3666
rect 48862 3614 48914 3666
rect 48914 3614 48916 3666
rect 48860 3612 48916 3614
rect 49868 5404 49924 5460
rect 49980 5180 50036 5236
rect 49644 4620 49700 4676
rect 49420 3724 49476 3780
rect 49980 4562 50036 4564
rect 49980 4510 49982 4562
rect 49982 4510 50034 4562
rect 50034 4510 50036 4562
rect 49980 4508 50036 4510
rect 49644 3724 49700 3780
rect 49756 3948 49812 4004
rect 49308 3666 49364 3668
rect 49308 3614 49310 3666
rect 49310 3614 49362 3666
rect 49362 3614 49364 3666
rect 49308 3612 49364 3614
rect 48076 3500 48132 3556
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 50876 7420 50932 7476
rect 50764 7308 50820 7364
rect 50876 6748 50932 6804
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 51212 15820 51268 15876
rect 51324 15708 51380 15764
rect 51436 12850 51492 12852
rect 51436 12798 51438 12850
rect 51438 12798 51490 12850
rect 51490 12798 51492 12850
rect 51436 12796 51492 12798
rect 52220 20524 52276 20580
rect 52332 20300 52388 20356
rect 51996 18956 52052 19012
rect 52108 19852 52164 19908
rect 51884 18562 51940 18564
rect 51884 18510 51886 18562
rect 51886 18510 51938 18562
rect 51938 18510 51940 18562
rect 51884 18508 51940 18510
rect 51772 18284 51828 18340
rect 51884 17948 51940 18004
rect 51772 17052 51828 17108
rect 52220 19068 52276 19124
rect 52444 18562 52500 18564
rect 52444 18510 52446 18562
rect 52446 18510 52498 18562
rect 52498 18510 52500 18562
rect 52444 18508 52500 18510
rect 52332 17778 52388 17780
rect 52332 17726 52334 17778
rect 52334 17726 52386 17778
rect 52386 17726 52388 17778
rect 52332 17724 52388 17726
rect 52220 16210 52276 16212
rect 52220 16158 52222 16210
rect 52222 16158 52274 16210
rect 52274 16158 52276 16210
rect 52220 16156 52276 16158
rect 51884 15708 51940 15764
rect 53564 37378 53620 37380
rect 53564 37326 53566 37378
rect 53566 37326 53618 37378
rect 53618 37326 53620 37378
rect 53564 37324 53620 37326
rect 53452 35420 53508 35476
rect 53788 37660 53844 37716
rect 54124 41356 54180 41412
rect 54572 41580 54628 41636
rect 54348 40908 54404 40964
rect 54236 39730 54292 39732
rect 54236 39678 54238 39730
rect 54238 39678 54290 39730
rect 54290 39678 54292 39730
rect 54236 39676 54292 39678
rect 54124 39004 54180 39060
rect 54460 39452 54516 39508
rect 54460 39004 54516 39060
rect 55020 43484 55076 43540
rect 55356 43596 55412 43652
rect 56028 48130 56084 48132
rect 56028 48078 56030 48130
rect 56030 48078 56082 48130
rect 56082 48078 56084 48130
rect 56028 48076 56084 48078
rect 56476 47628 56532 47684
rect 55692 47234 55748 47236
rect 55692 47182 55694 47234
rect 55694 47182 55746 47234
rect 55746 47182 55748 47234
rect 55692 47180 55748 47182
rect 56028 47068 56084 47124
rect 55692 46898 55748 46900
rect 55692 46846 55694 46898
rect 55694 46846 55746 46898
rect 55746 46846 55748 46898
rect 55692 46844 55748 46846
rect 56252 46956 56308 47012
rect 56588 46732 56644 46788
rect 56812 47068 56868 47124
rect 56588 46562 56644 46564
rect 56588 46510 56590 46562
rect 56590 46510 56642 46562
rect 56642 46510 56644 46562
rect 56588 46508 56644 46510
rect 55580 45836 55636 45892
rect 55804 45666 55860 45668
rect 55804 45614 55806 45666
rect 55806 45614 55858 45666
rect 55858 45614 55860 45666
rect 55804 45612 55860 45614
rect 55580 44828 55636 44884
rect 55916 44380 55972 44436
rect 55580 44322 55636 44324
rect 55580 44270 55582 44322
rect 55582 44270 55634 44322
rect 55634 44270 55636 44322
rect 55580 44268 55636 44270
rect 55468 43260 55524 43316
rect 55356 43036 55412 43092
rect 55132 42700 55188 42756
rect 55132 41132 55188 41188
rect 55244 41970 55300 41972
rect 55244 41918 55246 41970
rect 55246 41918 55298 41970
rect 55298 41918 55300 41970
rect 55244 41916 55300 41918
rect 55244 41020 55300 41076
rect 55132 40514 55188 40516
rect 55132 40462 55134 40514
rect 55134 40462 55186 40514
rect 55186 40462 55188 40514
rect 55132 40460 55188 40462
rect 55020 40402 55076 40404
rect 55020 40350 55022 40402
rect 55022 40350 55074 40402
rect 55074 40350 55076 40402
rect 55020 40348 55076 40350
rect 55580 42028 55636 42084
rect 55468 40908 55524 40964
rect 55580 41580 55636 41636
rect 55356 40348 55412 40404
rect 55468 40684 55524 40740
rect 54908 39506 54964 39508
rect 54908 39454 54910 39506
rect 54910 39454 54962 39506
rect 54962 39454 54964 39506
rect 54908 39452 54964 39454
rect 55020 39004 55076 39060
rect 54012 38220 54068 38276
rect 54908 38722 54964 38724
rect 54908 38670 54910 38722
rect 54910 38670 54962 38722
rect 54962 38670 54964 38722
rect 54908 38668 54964 38670
rect 55244 39618 55300 39620
rect 55244 39566 55246 39618
rect 55246 39566 55298 39618
rect 55298 39566 55300 39618
rect 55244 39564 55300 39566
rect 55244 38946 55300 38948
rect 55244 38894 55246 38946
rect 55246 38894 55298 38946
rect 55298 38894 55300 38946
rect 55244 38892 55300 38894
rect 53676 36370 53732 36372
rect 53676 36318 53678 36370
rect 53678 36318 53730 36370
rect 53730 36318 53732 36370
rect 53676 36316 53732 36318
rect 54124 36764 54180 36820
rect 53900 36482 53956 36484
rect 53900 36430 53902 36482
rect 53902 36430 53954 36482
rect 53954 36430 53956 36482
rect 53900 36428 53956 36430
rect 54012 35868 54068 35924
rect 53788 34914 53844 34916
rect 53788 34862 53790 34914
rect 53790 34862 53842 34914
rect 53842 34862 53844 34914
rect 53788 34860 53844 34862
rect 53564 34802 53620 34804
rect 53564 34750 53566 34802
rect 53566 34750 53618 34802
rect 53618 34750 53620 34802
rect 53564 34748 53620 34750
rect 54684 38220 54740 38276
rect 54460 34914 54516 34916
rect 54460 34862 54462 34914
rect 54462 34862 54514 34914
rect 54514 34862 54516 34914
rect 54460 34860 54516 34862
rect 54908 38050 54964 38052
rect 54908 37998 54910 38050
rect 54910 37998 54962 38050
rect 54962 37998 54964 38050
rect 54908 37996 54964 37998
rect 55020 37938 55076 37940
rect 55020 37886 55022 37938
rect 55022 37886 55074 37938
rect 55074 37886 55076 37938
rect 55020 37884 55076 37886
rect 54796 37826 54852 37828
rect 54796 37774 54798 37826
rect 54798 37774 54850 37826
rect 54850 37774 54852 37826
rect 54796 37772 54852 37774
rect 54796 35308 54852 35364
rect 54684 34690 54740 34692
rect 54684 34638 54686 34690
rect 54686 34638 54738 34690
rect 54738 34638 54740 34690
rect 54684 34636 54740 34638
rect 53676 33740 53732 33796
rect 53564 33516 53620 33572
rect 53340 33122 53396 33124
rect 53340 33070 53342 33122
rect 53342 33070 53394 33122
rect 53394 33070 53396 33122
rect 53340 33068 53396 33070
rect 53452 32732 53508 32788
rect 53340 31948 53396 32004
rect 53452 31500 53508 31556
rect 53900 34412 53956 34468
rect 54348 33458 54404 33460
rect 54348 33406 54350 33458
rect 54350 33406 54402 33458
rect 54402 33406 54404 33458
rect 54348 33404 54404 33406
rect 54012 33292 54068 33348
rect 53676 32396 53732 32452
rect 53676 31948 53732 32004
rect 53676 31666 53732 31668
rect 53676 31614 53678 31666
rect 53678 31614 53730 31666
rect 53730 31614 53732 31666
rect 53676 31612 53732 31614
rect 54012 32060 54068 32116
rect 53900 31724 53956 31780
rect 54124 30828 54180 30884
rect 52780 28252 52836 28308
rect 53340 29986 53396 29988
rect 53340 29934 53342 29986
rect 53342 29934 53394 29986
rect 53394 29934 53396 29986
rect 53340 29932 53396 29934
rect 53228 28812 53284 28868
rect 53116 28252 53172 28308
rect 53116 27804 53172 27860
rect 53004 27244 53060 27300
rect 53564 29260 53620 29316
rect 53788 30268 53844 30324
rect 54236 30492 54292 30548
rect 53564 28418 53620 28420
rect 53564 28366 53566 28418
rect 53566 28366 53618 28418
rect 53618 28366 53620 28418
rect 53564 28364 53620 28366
rect 53564 27298 53620 27300
rect 53564 27246 53566 27298
rect 53566 27246 53618 27298
rect 53618 27246 53620 27298
rect 53564 27244 53620 27246
rect 52780 26066 52836 26068
rect 52780 26014 52782 26066
rect 52782 26014 52834 26066
rect 52834 26014 52836 26066
rect 52780 26012 52836 26014
rect 52892 25900 52948 25956
rect 53004 25676 53060 25732
rect 52780 23884 52836 23940
rect 52780 22204 52836 22260
rect 52668 21474 52724 21476
rect 52668 21422 52670 21474
rect 52670 21422 52722 21474
rect 52722 21422 52724 21474
rect 52668 21420 52724 21422
rect 52892 21308 52948 21364
rect 52668 20860 52724 20916
rect 53004 20524 53060 20580
rect 53228 26348 53284 26404
rect 53340 26124 53396 26180
rect 53340 25564 53396 25620
rect 53452 25452 53508 25508
rect 53228 23042 53284 23044
rect 53228 22990 53230 23042
rect 53230 22990 53282 23042
rect 53282 22990 53284 23042
rect 53228 22988 53284 22990
rect 53676 26796 53732 26852
rect 53900 27804 53956 27860
rect 54236 27916 54292 27972
rect 54684 34130 54740 34132
rect 54684 34078 54686 34130
rect 54686 34078 54738 34130
rect 54738 34078 54740 34130
rect 54684 34076 54740 34078
rect 54572 33180 54628 33236
rect 54908 33852 54964 33908
rect 55132 36258 55188 36260
rect 55132 36206 55134 36258
rect 55134 36206 55186 36258
rect 55186 36206 55188 36258
rect 55132 36204 55188 36206
rect 56364 44994 56420 44996
rect 56364 44942 56366 44994
rect 56366 44942 56418 44994
rect 56418 44942 56420 44994
rect 56364 44940 56420 44942
rect 56140 44044 56196 44100
rect 56364 43260 56420 43316
rect 56252 42754 56308 42756
rect 56252 42702 56254 42754
rect 56254 42702 56306 42754
rect 56306 42702 56308 42754
rect 56252 42700 56308 42702
rect 56140 42082 56196 42084
rect 56140 42030 56142 42082
rect 56142 42030 56194 42082
rect 56194 42030 56196 42082
rect 56140 42028 56196 42030
rect 56028 40684 56084 40740
rect 56140 41132 56196 41188
rect 56588 43708 56644 43764
rect 56588 43426 56644 43428
rect 56588 43374 56590 43426
rect 56590 43374 56642 43426
rect 56642 43374 56644 43426
rect 56588 43372 56644 43374
rect 56476 41580 56532 41636
rect 55692 40460 55748 40516
rect 55804 40402 55860 40404
rect 55804 40350 55806 40402
rect 55806 40350 55858 40402
rect 55858 40350 55860 40402
rect 55804 40348 55860 40350
rect 56252 41074 56308 41076
rect 56252 41022 56254 41074
rect 56254 41022 56306 41074
rect 56306 41022 56308 41074
rect 56252 41020 56308 41022
rect 56364 40962 56420 40964
rect 56364 40910 56366 40962
rect 56366 40910 56418 40962
rect 56418 40910 56420 40962
rect 56364 40908 56420 40910
rect 55916 39676 55972 39732
rect 55804 39506 55860 39508
rect 55804 39454 55806 39506
rect 55806 39454 55858 39506
rect 55858 39454 55860 39506
rect 55804 39452 55860 39454
rect 55692 38892 55748 38948
rect 57148 53788 57204 53844
rect 57036 49644 57092 49700
rect 57932 50764 57988 50820
rect 57484 47740 57540 47796
rect 57372 46562 57428 46564
rect 57372 46510 57374 46562
rect 57374 46510 57426 46562
rect 57426 46510 57428 46562
rect 57372 46508 57428 46510
rect 57596 45948 57652 46004
rect 57484 45218 57540 45220
rect 57484 45166 57486 45218
rect 57486 45166 57538 45218
rect 57538 45166 57540 45218
rect 57484 45164 57540 45166
rect 57148 44604 57204 44660
rect 57596 44492 57652 44548
rect 57820 46786 57876 46788
rect 57820 46734 57822 46786
rect 57822 46734 57874 46786
rect 57874 46734 57876 46786
rect 57820 46732 57876 46734
rect 57820 45948 57876 46004
rect 58828 45612 58884 45668
rect 58044 45164 58100 45220
rect 57148 44098 57204 44100
rect 57148 44046 57150 44098
rect 57150 44046 57202 44098
rect 57202 44046 57204 44098
rect 57148 44044 57204 44046
rect 56924 43372 56980 43428
rect 57820 43372 57876 43428
rect 56812 41356 56868 41412
rect 56476 40124 56532 40180
rect 56812 40012 56868 40068
rect 56140 39676 56196 39732
rect 56700 39788 56756 39844
rect 56140 39116 56196 39172
rect 56364 39340 56420 39396
rect 55804 38556 55860 38612
rect 56252 38610 56308 38612
rect 56252 38558 56254 38610
rect 56254 38558 56306 38610
rect 56306 38558 56308 38610
rect 56252 38556 56308 38558
rect 56140 37772 56196 37828
rect 55804 37212 55860 37268
rect 55692 36988 55748 37044
rect 55580 35532 55636 35588
rect 55468 35420 55524 35476
rect 55132 34972 55188 35028
rect 55132 34300 55188 34356
rect 54572 32060 54628 32116
rect 54908 31388 54964 31444
rect 54796 30380 54852 30436
rect 54684 30210 54740 30212
rect 54684 30158 54686 30210
rect 54686 30158 54738 30210
rect 54738 30158 54740 30210
rect 54684 30156 54740 30158
rect 54684 29932 54740 29988
rect 54684 29036 54740 29092
rect 55692 34972 55748 35028
rect 55356 34914 55412 34916
rect 55356 34862 55358 34914
rect 55358 34862 55410 34914
rect 55410 34862 55412 34914
rect 55356 34860 55412 34862
rect 55804 34860 55860 34916
rect 55580 34748 55636 34804
rect 55692 34690 55748 34692
rect 55692 34638 55694 34690
rect 55694 34638 55746 34690
rect 55746 34638 55748 34690
rect 55692 34636 55748 34638
rect 55244 33852 55300 33908
rect 55244 31836 55300 31892
rect 55580 34188 55636 34244
rect 55468 33740 55524 33796
rect 55356 31164 55412 31220
rect 55132 29986 55188 29988
rect 55132 29934 55134 29986
rect 55134 29934 55186 29986
rect 55186 29934 55188 29986
rect 55132 29932 55188 29934
rect 54460 28252 54516 28308
rect 54348 27580 54404 27636
rect 54460 28028 54516 28084
rect 54124 27020 54180 27076
rect 54348 27132 54404 27188
rect 54236 26908 54292 26964
rect 53676 25676 53732 25732
rect 54684 27916 54740 27972
rect 54460 26908 54516 26964
rect 53676 25228 53732 25284
rect 53564 24722 53620 24724
rect 53564 24670 53566 24722
rect 53566 24670 53618 24722
rect 53618 24670 53620 24722
rect 53564 24668 53620 24670
rect 53452 23938 53508 23940
rect 53452 23886 53454 23938
rect 53454 23886 53506 23938
rect 53506 23886 53508 23938
rect 53452 23884 53508 23886
rect 53676 23436 53732 23492
rect 53452 23324 53508 23380
rect 53452 23100 53508 23156
rect 54012 25116 54068 25172
rect 54124 25004 54180 25060
rect 54348 26796 54404 26852
rect 54012 24946 54068 24948
rect 54012 24894 54014 24946
rect 54014 24894 54066 24946
rect 54066 24894 54068 24946
rect 54012 24892 54068 24894
rect 53900 23884 53956 23940
rect 53788 22146 53844 22148
rect 53788 22094 53790 22146
rect 53790 22094 53842 22146
rect 53842 22094 53844 22146
rect 53788 22092 53844 22094
rect 53452 21532 53508 21588
rect 53340 21474 53396 21476
rect 53340 21422 53342 21474
rect 53342 21422 53394 21474
rect 53394 21422 53396 21474
rect 53340 21420 53396 21422
rect 53788 21586 53844 21588
rect 53788 21534 53790 21586
rect 53790 21534 53842 21586
rect 53842 21534 53844 21586
rect 53788 21532 53844 21534
rect 53340 21084 53396 21140
rect 53564 20242 53620 20244
rect 53564 20190 53566 20242
rect 53566 20190 53618 20242
rect 53618 20190 53620 20242
rect 53564 20188 53620 20190
rect 52780 18732 52836 18788
rect 53116 19852 53172 19908
rect 52668 17948 52724 18004
rect 52892 16156 52948 16212
rect 53004 17724 53060 17780
rect 53004 16940 53060 16996
rect 52220 15708 52276 15764
rect 52780 15708 52836 15764
rect 51884 15538 51940 15540
rect 51884 15486 51886 15538
rect 51886 15486 51938 15538
rect 51938 15486 51940 15538
rect 51884 15484 51940 15486
rect 52220 15372 52276 15428
rect 52444 15202 52500 15204
rect 52444 15150 52446 15202
rect 52446 15150 52498 15202
rect 52498 15150 52500 15202
rect 52444 15148 52500 15150
rect 52332 15036 52388 15092
rect 51772 13916 51828 13972
rect 52108 14140 52164 14196
rect 52108 13692 52164 13748
rect 52332 13746 52388 13748
rect 52332 13694 52334 13746
rect 52334 13694 52386 13746
rect 52386 13694 52388 13746
rect 52332 13692 52388 13694
rect 51660 13634 51716 13636
rect 51660 13582 51662 13634
rect 51662 13582 51714 13634
rect 51714 13582 51716 13634
rect 51660 13580 51716 13582
rect 51772 12962 51828 12964
rect 51772 12910 51774 12962
rect 51774 12910 51826 12962
rect 51826 12910 51828 12962
rect 51772 12908 51828 12910
rect 51212 12066 51268 12068
rect 51212 12014 51214 12066
rect 51214 12014 51266 12066
rect 51266 12014 51268 12066
rect 51212 12012 51268 12014
rect 51324 11394 51380 11396
rect 51324 11342 51326 11394
rect 51326 11342 51378 11394
rect 51378 11342 51380 11394
rect 51324 11340 51380 11342
rect 51212 10610 51268 10612
rect 51212 10558 51214 10610
rect 51214 10558 51266 10610
rect 51266 10558 51268 10610
rect 51212 10556 51268 10558
rect 51324 9996 51380 10052
rect 51436 10108 51492 10164
rect 51100 9266 51156 9268
rect 51100 9214 51102 9266
rect 51102 9214 51154 9266
rect 51154 9214 51156 9266
rect 51100 9212 51156 9214
rect 51100 8988 51156 9044
rect 51660 11676 51716 11732
rect 51660 11004 51716 11060
rect 51772 10834 51828 10836
rect 51772 10782 51774 10834
rect 51774 10782 51826 10834
rect 51826 10782 51828 10834
rect 51772 10780 51828 10782
rect 51996 13580 52052 13636
rect 52332 12850 52388 12852
rect 52332 12798 52334 12850
rect 52334 12798 52386 12850
rect 52386 12798 52388 12850
rect 52332 12796 52388 12798
rect 52108 12684 52164 12740
rect 52332 12572 52388 12628
rect 51996 10780 52052 10836
rect 52108 11564 52164 11620
rect 52108 10668 52164 10724
rect 51884 9884 51940 9940
rect 51212 8428 51268 8484
rect 51548 8876 51604 8932
rect 51212 8258 51268 8260
rect 51212 8206 51214 8258
rect 51214 8206 51266 8258
rect 51266 8206 51268 8258
rect 51212 8204 51268 8206
rect 51660 8092 51716 8148
rect 51884 9436 51940 9492
rect 51212 6690 51268 6692
rect 51212 6638 51214 6690
rect 51214 6638 51266 6690
rect 51266 6638 51268 6690
rect 51212 6636 51268 6638
rect 51772 7644 51828 7700
rect 51884 6636 51940 6692
rect 51436 4844 51492 4900
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50428 3836 50484 3892
rect 49756 3554 49812 3556
rect 49756 3502 49758 3554
rect 49758 3502 49810 3554
rect 49810 3502 49812 3554
rect 49756 3500 49812 3502
rect 50204 3724 50260 3780
rect 51100 3666 51156 3668
rect 51100 3614 51102 3666
rect 51102 3614 51154 3666
rect 51154 3614 51156 3666
rect 51100 3612 51156 3614
rect 52108 9548 52164 9604
rect 52668 12908 52724 12964
rect 53228 19180 53284 19236
rect 53676 20076 53732 20132
rect 53452 19458 53508 19460
rect 53452 19406 53454 19458
rect 53454 19406 53506 19458
rect 53506 19406 53508 19458
rect 53452 19404 53508 19406
rect 53452 19180 53508 19236
rect 53228 18396 53284 18452
rect 53340 18338 53396 18340
rect 53340 18286 53342 18338
rect 53342 18286 53394 18338
rect 53394 18286 53396 18338
rect 53340 18284 53396 18286
rect 53228 17724 53284 17780
rect 54012 21084 54068 21140
rect 54012 20802 54068 20804
rect 54012 20750 54014 20802
rect 54014 20750 54066 20802
rect 54066 20750 54068 20802
rect 54012 20748 54068 20750
rect 54236 23378 54292 23380
rect 54236 23326 54238 23378
rect 54238 23326 54290 23378
rect 54290 23326 54292 23378
rect 54236 23324 54292 23326
rect 54236 21868 54292 21924
rect 54460 26684 54516 26740
rect 54460 26124 54516 26180
rect 54124 20188 54180 20244
rect 54348 20188 54404 20244
rect 54348 20018 54404 20020
rect 54348 19966 54350 20018
rect 54350 19966 54402 20018
rect 54402 19966 54404 20018
rect 54348 19964 54404 19966
rect 54572 23154 54628 23156
rect 54572 23102 54574 23154
rect 54574 23102 54626 23154
rect 54626 23102 54628 23154
rect 54572 23100 54628 23102
rect 54908 29426 54964 29428
rect 54908 29374 54910 29426
rect 54910 29374 54962 29426
rect 54962 29374 54964 29426
rect 54908 29372 54964 29374
rect 55132 29426 55188 29428
rect 55132 29374 55134 29426
rect 55134 29374 55186 29426
rect 55186 29374 55188 29426
rect 55132 29372 55188 29374
rect 55132 28028 55188 28084
rect 55580 30098 55636 30100
rect 55580 30046 55582 30098
rect 55582 30046 55634 30098
rect 55634 30046 55636 30098
rect 55580 30044 55636 30046
rect 55468 29372 55524 29428
rect 55356 28588 55412 28644
rect 55244 27132 55300 27188
rect 55580 29202 55636 29204
rect 55580 29150 55582 29202
rect 55582 29150 55634 29202
rect 55634 29150 55636 29202
rect 55580 29148 55636 29150
rect 56588 37100 56644 37156
rect 56588 35810 56644 35812
rect 56588 35758 56590 35810
rect 56590 35758 56642 35810
rect 56642 35758 56644 35810
rect 56588 35756 56644 35758
rect 56252 35644 56308 35700
rect 56028 35532 56084 35588
rect 55804 33628 55860 33684
rect 55916 33234 55972 33236
rect 55916 33182 55918 33234
rect 55918 33182 55970 33234
rect 55970 33182 55972 33234
rect 55916 33180 55972 33182
rect 56252 35474 56308 35476
rect 56252 35422 56254 35474
rect 56254 35422 56306 35474
rect 56306 35422 56308 35474
rect 56252 35420 56308 35422
rect 56588 34802 56644 34804
rect 56588 34750 56590 34802
rect 56590 34750 56642 34802
rect 56642 34750 56644 34802
rect 56588 34748 56644 34750
rect 56252 34524 56308 34580
rect 57036 39788 57092 39844
rect 57036 39452 57092 39508
rect 56924 37884 56980 37940
rect 57372 42530 57428 42532
rect 57372 42478 57374 42530
rect 57374 42478 57426 42530
rect 57426 42478 57428 42530
rect 57372 42476 57428 42478
rect 57372 41858 57428 41860
rect 57372 41806 57374 41858
rect 57374 41806 57426 41858
rect 57426 41806 57428 41858
rect 57372 41804 57428 41806
rect 57820 41858 57876 41860
rect 57820 41806 57822 41858
rect 57822 41806 57874 41858
rect 57874 41806 57876 41858
rect 57820 41804 57876 41806
rect 58156 43708 58212 43764
rect 57708 39618 57764 39620
rect 57708 39566 57710 39618
rect 57710 39566 57762 39618
rect 57762 39566 57764 39618
rect 57708 39564 57764 39566
rect 57372 39058 57428 39060
rect 57372 39006 57374 39058
rect 57374 39006 57426 39058
rect 57426 39006 57428 39058
rect 57372 39004 57428 39006
rect 57596 39394 57652 39396
rect 57596 39342 57598 39394
rect 57598 39342 57650 39394
rect 57650 39342 57652 39394
rect 57596 39340 57652 39342
rect 57596 39116 57652 39172
rect 57708 38946 57764 38948
rect 57708 38894 57710 38946
rect 57710 38894 57762 38946
rect 57762 38894 57764 38946
rect 57708 38892 57764 38894
rect 57484 38780 57540 38836
rect 57596 38050 57652 38052
rect 57596 37998 57598 38050
rect 57598 37998 57650 38050
rect 57650 37998 57652 38050
rect 57596 37996 57652 37998
rect 57484 37100 57540 37156
rect 56812 36370 56868 36372
rect 56812 36318 56814 36370
rect 56814 36318 56866 36370
rect 56866 36318 56868 36370
rect 56812 36316 56868 36318
rect 57260 36092 57316 36148
rect 57036 35644 57092 35700
rect 56924 35026 56980 35028
rect 56924 34974 56926 35026
rect 56926 34974 56978 35026
rect 56978 34974 56980 35026
rect 56924 34972 56980 34974
rect 56588 34130 56644 34132
rect 56588 34078 56590 34130
rect 56590 34078 56642 34130
rect 56642 34078 56644 34130
rect 56588 34076 56644 34078
rect 56476 33516 56532 33572
rect 56140 31948 56196 32004
rect 56028 31612 56084 31668
rect 55916 30940 55972 30996
rect 56588 32562 56644 32564
rect 56588 32510 56590 32562
rect 56590 32510 56642 32562
rect 56642 32510 56644 32562
rect 56588 32508 56644 32510
rect 57260 33404 57316 33460
rect 56812 32396 56868 32452
rect 56924 33180 56980 33236
rect 56812 31724 56868 31780
rect 56028 29426 56084 29428
rect 56028 29374 56030 29426
rect 56030 29374 56082 29426
rect 56082 29374 56084 29426
rect 56028 29372 56084 29374
rect 55804 29260 55860 29316
rect 56140 29148 56196 29204
rect 54908 26908 54964 26964
rect 55132 26962 55188 26964
rect 55132 26910 55134 26962
rect 55134 26910 55186 26962
rect 55186 26910 55188 26962
rect 55132 26908 55188 26910
rect 56028 28924 56084 28980
rect 55804 28140 55860 28196
rect 55804 27298 55860 27300
rect 55804 27246 55806 27298
rect 55806 27246 55858 27298
rect 55858 27246 55860 27298
rect 55804 27244 55860 27246
rect 55916 28700 55972 28756
rect 56476 29426 56532 29428
rect 56476 29374 56478 29426
rect 56478 29374 56530 29426
rect 56530 29374 56532 29426
rect 56476 29372 56532 29374
rect 56252 28252 56308 28308
rect 56028 28028 56084 28084
rect 55916 27356 55972 27412
rect 55580 27020 55636 27076
rect 54908 26290 54964 26292
rect 54908 26238 54910 26290
rect 54910 26238 54962 26290
rect 54962 26238 54964 26290
rect 54908 26236 54964 26238
rect 55244 25506 55300 25508
rect 55244 25454 55246 25506
rect 55246 25454 55298 25506
rect 55298 25454 55300 25506
rect 55244 25452 55300 25454
rect 54796 25116 54852 25172
rect 55132 24444 55188 24500
rect 56700 30604 56756 30660
rect 56700 30044 56756 30100
rect 56700 29426 56756 29428
rect 56700 29374 56702 29426
rect 56702 29374 56754 29426
rect 56754 29374 56756 29426
rect 56700 29372 56756 29374
rect 56700 28700 56756 28756
rect 57484 35420 57540 35476
rect 57820 38444 57876 38500
rect 57932 38332 57988 38388
rect 57820 36092 57876 36148
rect 57708 35698 57764 35700
rect 57708 35646 57710 35698
rect 57710 35646 57762 35698
rect 57762 35646 57764 35698
rect 57708 35644 57764 35646
rect 57148 32508 57204 32564
rect 57148 32060 57204 32116
rect 56812 28028 56868 28084
rect 57372 31836 57428 31892
rect 58156 38108 58212 38164
rect 58268 37212 58324 37268
rect 58044 34972 58100 35028
rect 58156 36316 58212 36372
rect 58044 34690 58100 34692
rect 58044 34638 58046 34690
rect 58046 34638 58098 34690
rect 58098 34638 58100 34690
rect 58044 34636 58100 34638
rect 58044 34018 58100 34020
rect 58044 33966 58046 34018
rect 58046 33966 58098 34018
rect 58098 33966 58100 34018
rect 58044 33964 58100 33966
rect 57932 33292 57988 33348
rect 57932 32620 57988 32676
rect 57820 32562 57876 32564
rect 57820 32510 57822 32562
rect 57822 32510 57874 32562
rect 57874 32510 57876 32562
rect 57820 32508 57876 32510
rect 57484 31778 57540 31780
rect 57484 31726 57486 31778
rect 57486 31726 57538 31778
rect 57538 31726 57540 31778
rect 57484 31724 57540 31726
rect 57484 30268 57540 30324
rect 57596 30940 57652 30996
rect 57820 31500 57876 31556
rect 57260 29372 57316 29428
rect 57148 28364 57204 28420
rect 57148 28028 57204 28084
rect 56588 27916 56644 27972
rect 57596 28418 57652 28420
rect 57596 28366 57598 28418
rect 57598 28366 57650 28418
rect 57650 28366 57652 28418
rect 57596 28364 57652 28366
rect 58044 28700 58100 28756
rect 57484 27970 57540 27972
rect 57484 27918 57486 27970
rect 57486 27918 57538 27970
rect 57538 27918 57540 27970
rect 57484 27916 57540 27918
rect 56476 27356 56532 27412
rect 56028 26908 56084 26964
rect 56028 25564 56084 25620
rect 55692 24892 55748 24948
rect 56812 27244 56868 27300
rect 56588 26178 56644 26180
rect 56588 26126 56590 26178
rect 56590 26126 56642 26178
rect 56642 26126 56644 26178
rect 56588 26124 56644 26126
rect 56588 25506 56644 25508
rect 56588 25454 56590 25506
rect 56590 25454 56642 25506
rect 56642 25454 56644 25506
rect 56588 25452 56644 25454
rect 56588 25228 56644 25284
rect 55804 24834 55860 24836
rect 55804 24782 55806 24834
rect 55806 24782 55858 24834
rect 55858 24782 55860 24834
rect 55804 24780 55860 24782
rect 55916 24108 55972 24164
rect 54684 22316 54740 22372
rect 54908 23996 54964 24052
rect 54684 21474 54740 21476
rect 54684 21422 54686 21474
rect 54686 21422 54738 21474
rect 54738 21422 54740 21474
rect 54684 21420 54740 21422
rect 54572 20524 54628 20580
rect 54460 19852 54516 19908
rect 54012 19346 54068 19348
rect 54012 19294 54014 19346
rect 54014 19294 54066 19346
rect 54066 19294 54068 19346
rect 54012 19292 54068 19294
rect 53788 19234 53844 19236
rect 53788 19182 53790 19234
rect 53790 19182 53842 19234
rect 53842 19182 53844 19234
rect 53788 19180 53844 19182
rect 53676 18508 53732 18564
rect 53788 18338 53844 18340
rect 53788 18286 53790 18338
rect 53790 18286 53842 18338
rect 53842 18286 53844 18338
rect 53788 18284 53844 18286
rect 53564 17836 53620 17892
rect 53452 17724 53508 17780
rect 54684 19010 54740 19012
rect 54684 18958 54686 19010
rect 54686 18958 54738 19010
rect 54738 18958 54740 19010
rect 54684 18956 54740 18958
rect 55244 23378 55300 23380
rect 55244 23326 55246 23378
rect 55246 23326 55298 23378
rect 55298 23326 55300 23378
rect 55244 23324 55300 23326
rect 55132 22988 55188 23044
rect 55580 23100 55636 23156
rect 55916 22988 55972 23044
rect 55020 22370 55076 22372
rect 55020 22318 55022 22370
rect 55022 22318 55074 22370
rect 55074 22318 55076 22370
rect 55020 22316 55076 22318
rect 55020 20802 55076 20804
rect 55020 20750 55022 20802
rect 55022 20750 55074 20802
rect 55074 20750 55076 20802
rect 55020 20748 55076 20750
rect 54908 18732 54964 18788
rect 54796 18674 54852 18676
rect 54796 18622 54798 18674
rect 54798 18622 54850 18674
rect 54850 18622 54852 18674
rect 54796 18620 54852 18622
rect 54012 18508 54068 18564
rect 53228 16268 53284 16324
rect 53340 16716 53396 16772
rect 53004 15426 53060 15428
rect 53004 15374 53006 15426
rect 53006 15374 53058 15426
rect 53058 15374 53060 15426
rect 53004 15372 53060 15374
rect 53900 17276 53956 17332
rect 53564 17106 53620 17108
rect 53564 17054 53566 17106
rect 53566 17054 53618 17106
rect 53618 17054 53620 17106
rect 53564 17052 53620 17054
rect 53564 16828 53620 16884
rect 53676 16716 53732 16772
rect 53564 16156 53620 16212
rect 53788 16380 53844 16436
rect 53676 15708 53732 15764
rect 53340 14252 53396 14308
rect 53228 13858 53284 13860
rect 53228 13806 53230 13858
rect 53230 13806 53282 13858
rect 53282 13806 53284 13858
rect 53228 13804 53284 13806
rect 53116 13692 53172 13748
rect 53564 14140 53620 14196
rect 53340 12012 53396 12068
rect 53340 11676 53396 11732
rect 53340 11282 53396 11284
rect 53340 11230 53342 11282
rect 53342 11230 53394 11282
rect 53394 11230 53396 11282
rect 53340 11228 53396 11230
rect 52668 10834 52724 10836
rect 52668 10782 52670 10834
rect 52670 10782 52722 10834
rect 52722 10782 52724 10834
rect 52668 10780 52724 10782
rect 52444 9938 52500 9940
rect 52444 9886 52446 9938
rect 52446 9886 52498 9938
rect 52498 9886 52500 9938
rect 52444 9884 52500 9886
rect 52332 9660 52388 9716
rect 53004 10220 53060 10276
rect 53564 10834 53620 10836
rect 53564 10782 53566 10834
rect 53566 10782 53618 10834
rect 53618 10782 53620 10834
rect 53564 10780 53620 10782
rect 52556 9436 52612 9492
rect 52892 9660 52948 9716
rect 52556 9212 52612 9268
rect 52220 8428 52276 8484
rect 52332 8652 52388 8708
rect 52108 8146 52164 8148
rect 52108 8094 52110 8146
rect 52110 8094 52162 8146
rect 52162 8094 52164 8146
rect 52108 8092 52164 8094
rect 52108 7644 52164 7700
rect 52108 6412 52164 6468
rect 51996 4060 52052 4116
rect 51996 3836 52052 3892
rect 50540 3500 50596 3556
rect 51772 3388 51828 3444
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 52780 7980 52836 8036
rect 52556 6802 52612 6804
rect 52556 6750 52558 6802
rect 52558 6750 52610 6802
rect 52610 6750 52612 6802
rect 52556 6748 52612 6750
rect 53788 14476 53844 14532
rect 54908 18562 54964 18564
rect 54908 18510 54910 18562
rect 54910 18510 54962 18562
rect 54962 18510 54964 18562
rect 54908 18508 54964 18510
rect 54236 18450 54292 18452
rect 54236 18398 54238 18450
rect 54238 18398 54290 18450
rect 54290 18398 54292 18450
rect 54236 18396 54292 18398
rect 54684 18450 54740 18452
rect 54684 18398 54686 18450
rect 54686 18398 54738 18450
rect 54738 18398 54740 18450
rect 54684 18396 54740 18398
rect 54796 17836 54852 17892
rect 54684 17500 54740 17556
rect 54572 17442 54628 17444
rect 54572 17390 54574 17442
rect 54574 17390 54626 17442
rect 54626 17390 54628 17442
rect 54572 17388 54628 17390
rect 54572 17164 54628 17220
rect 54460 17052 54516 17108
rect 54012 16828 54068 16884
rect 54124 16492 54180 16548
rect 54012 15484 54068 15540
rect 54124 16098 54180 16100
rect 54124 16046 54126 16098
rect 54126 16046 54178 16098
rect 54178 16046 54180 16098
rect 54124 16044 54180 16046
rect 54684 16210 54740 16212
rect 54684 16158 54686 16210
rect 54686 16158 54738 16210
rect 54738 16158 54740 16210
rect 54684 16156 54740 16158
rect 54684 15426 54740 15428
rect 54684 15374 54686 15426
rect 54686 15374 54738 15426
rect 54738 15374 54740 15426
rect 54684 15372 54740 15374
rect 54236 15036 54292 15092
rect 54684 14924 54740 14980
rect 53900 13522 53956 13524
rect 53900 13470 53902 13522
rect 53902 13470 53954 13522
rect 53954 13470 53956 13522
rect 53900 13468 53956 13470
rect 54236 13634 54292 13636
rect 54236 13582 54238 13634
rect 54238 13582 54290 13634
rect 54290 13582 54292 13634
rect 54236 13580 54292 13582
rect 54124 12684 54180 12740
rect 54460 13746 54516 13748
rect 54460 13694 54462 13746
rect 54462 13694 54514 13746
rect 54514 13694 54516 13746
rect 54460 13692 54516 13694
rect 54348 12572 54404 12628
rect 54348 12066 54404 12068
rect 54348 12014 54350 12066
rect 54350 12014 54402 12066
rect 54402 12014 54404 12066
rect 54348 12012 54404 12014
rect 54236 11900 54292 11956
rect 53676 9266 53732 9268
rect 53676 9214 53678 9266
rect 53678 9214 53730 9266
rect 53730 9214 53732 9266
rect 53676 9212 53732 9214
rect 53788 9996 53844 10052
rect 54012 9212 54068 9268
rect 53116 7980 53172 8036
rect 53228 8652 53284 8708
rect 53004 6524 53060 6580
rect 53116 7756 53172 7812
rect 53340 8370 53396 8372
rect 53340 8318 53342 8370
rect 53342 8318 53394 8370
rect 53394 8318 53396 8370
rect 53340 8316 53396 8318
rect 53452 8204 53508 8260
rect 53788 8764 53844 8820
rect 53564 7644 53620 7700
rect 53564 6636 53620 6692
rect 52444 5292 52500 5348
rect 53340 5292 53396 5348
rect 53788 5292 53844 5348
rect 52444 5122 52500 5124
rect 52444 5070 52446 5122
rect 52446 5070 52498 5122
rect 52498 5070 52500 5122
rect 52444 5068 52500 5070
rect 52332 4508 52388 4564
rect 52556 4338 52612 4340
rect 52556 4286 52558 4338
rect 52558 4286 52610 4338
rect 52610 4286 52612 4338
rect 52556 4284 52612 4286
rect 52556 3948 52612 4004
rect 52892 4172 52948 4228
rect 52892 3612 52948 3668
rect 52780 3554 52836 3556
rect 52780 3502 52782 3554
rect 52782 3502 52834 3554
rect 52834 3502 52836 3554
rect 52780 3500 52836 3502
rect 53452 3388 53508 3444
rect 52220 2716 52276 2772
rect 54348 9266 54404 9268
rect 54348 9214 54350 9266
rect 54350 9214 54402 9266
rect 54402 9214 54404 9266
rect 54348 9212 54404 9214
rect 54236 8204 54292 8260
rect 54236 8034 54292 8036
rect 54236 7982 54238 8034
rect 54238 7982 54290 8034
rect 54290 7982 54292 8034
rect 54236 7980 54292 7982
rect 54684 12796 54740 12852
rect 55244 19852 55300 19908
rect 55468 22540 55524 22596
rect 55692 22540 55748 22596
rect 55804 22482 55860 22484
rect 55804 22430 55806 22482
rect 55806 22430 55858 22482
rect 55858 22430 55860 22482
rect 55804 22428 55860 22430
rect 55692 22092 55748 22148
rect 55580 20636 55636 20692
rect 55916 21980 55972 22036
rect 56588 23938 56644 23940
rect 56588 23886 56590 23938
rect 56590 23886 56642 23938
rect 56642 23886 56644 23938
rect 56588 23884 56644 23886
rect 56476 23212 56532 23268
rect 56476 22988 56532 23044
rect 56588 22594 56644 22596
rect 56588 22542 56590 22594
rect 56590 22542 56642 22594
rect 56642 22542 56644 22594
rect 56588 22540 56644 22542
rect 56700 22146 56756 22148
rect 56700 22094 56702 22146
rect 56702 22094 56754 22146
rect 56754 22094 56756 22146
rect 56700 22092 56756 22094
rect 56364 21698 56420 21700
rect 56364 21646 56366 21698
rect 56366 21646 56418 21698
rect 56418 21646 56420 21698
rect 56364 21644 56420 21646
rect 55692 21532 55748 21588
rect 55468 19852 55524 19908
rect 54908 17442 54964 17444
rect 54908 17390 54910 17442
rect 54910 17390 54962 17442
rect 54962 17390 54964 17442
rect 54908 17388 54964 17390
rect 55020 16604 55076 16660
rect 54908 15820 54964 15876
rect 54908 14476 54964 14532
rect 54908 13580 54964 13636
rect 55020 13692 55076 13748
rect 56028 20188 56084 20244
rect 56364 20524 56420 20580
rect 55468 19010 55524 19012
rect 55468 18958 55470 19010
rect 55470 18958 55522 19010
rect 55522 18958 55524 19010
rect 55468 18956 55524 18958
rect 55804 19964 55860 20020
rect 55804 19122 55860 19124
rect 55804 19070 55806 19122
rect 55806 19070 55858 19122
rect 55858 19070 55860 19122
rect 55804 19068 55860 19070
rect 56252 19010 56308 19012
rect 56252 18958 56254 19010
rect 56254 18958 56306 19010
rect 56306 18958 56308 19010
rect 56252 18956 56308 18958
rect 55356 17164 55412 17220
rect 55804 18508 55860 18564
rect 55580 18060 55636 18116
rect 55916 18396 55972 18452
rect 56252 17948 56308 18004
rect 56700 21586 56756 21588
rect 56700 21534 56702 21586
rect 56702 21534 56754 21586
rect 56754 21534 56756 21586
rect 56700 21532 56756 21534
rect 56588 21308 56644 21364
rect 56476 20076 56532 20132
rect 56700 20130 56756 20132
rect 56700 20078 56702 20130
rect 56702 20078 56754 20130
rect 56754 20078 56756 20130
rect 56700 20076 56756 20078
rect 57148 26850 57204 26852
rect 57148 26798 57150 26850
rect 57150 26798 57202 26850
rect 57202 26798 57204 26850
rect 57148 26796 57204 26798
rect 57484 26850 57540 26852
rect 57484 26798 57486 26850
rect 57486 26798 57538 26850
rect 57538 26798 57540 26850
rect 57484 26796 57540 26798
rect 57484 25004 57540 25060
rect 57260 24668 57316 24724
rect 56924 22258 56980 22260
rect 56924 22206 56926 22258
rect 56926 22206 56978 22258
rect 56978 22206 56980 22258
rect 56924 22204 56980 22206
rect 56812 19292 56868 19348
rect 56588 19180 56644 19236
rect 56924 19122 56980 19124
rect 56924 19070 56926 19122
rect 56926 19070 56978 19122
rect 56978 19070 56980 19122
rect 56924 19068 56980 19070
rect 57148 23714 57204 23716
rect 57148 23662 57150 23714
rect 57150 23662 57202 23714
rect 57202 23662 57204 23714
rect 57148 23660 57204 23662
rect 57820 27970 57876 27972
rect 57820 27918 57822 27970
rect 57822 27918 57874 27970
rect 57874 27918 57876 27970
rect 57820 27916 57876 27918
rect 57932 27186 57988 27188
rect 57932 27134 57934 27186
rect 57934 27134 57986 27186
rect 57986 27134 57988 27186
rect 57932 27132 57988 27134
rect 57708 26572 57764 26628
rect 57820 26796 57876 26852
rect 57820 25900 57876 25956
rect 57932 26012 57988 26068
rect 57708 25282 57764 25284
rect 57708 25230 57710 25282
rect 57710 25230 57762 25282
rect 57762 25230 57764 25282
rect 57708 25228 57764 25230
rect 57484 24108 57540 24164
rect 57484 23884 57540 23940
rect 56476 18674 56532 18676
rect 56476 18622 56478 18674
rect 56478 18622 56530 18674
rect 56530 18622 56532 18674
rect 56476 18620 56532 18622
rect 57036 18620 57092 18676
rect 55692 17554 55748 17556
rect 55692 17502 55694 17554
rect 55694 17502 55746 17554
rect 55746 17502 55748 17554
rect 55692 17500 55748 17502
rect 55580 17442 55636 17444
rect 55580 17390 55582 17442
rect 55582 17390 55634 17442
rect 55634 17390 55636 17442
rect 55580 17388 55636 17390
rect 55356 16044 55412 16100
rect 56252 17388 56308 17444
rect 55916 16828 55972 16884
rect 55468 15426 55524 15428
rect 55468 15374 55470 15426
rect 55470 15374 55522 15426
rect 55522 15374 55524 15426
rect 55468 15372 55524 15374
rect 55580 15484 55636 15540
rect 55356 14140 55412 14196
rect 55692 15090 55748 15092
rect 55692 15038 55694 15090
rect 55694 15038 55746 15090
rect 55746 15038 55748 15090
rect 55692 15036 55748 15038
rect 55692 14364 55748 14420
rect 55692 13746 55748 13748
rect 55692 13694 55694 13746
rect 55694 13694 55746 13746
rect 55746 13694 55748 13746
rect 55692 13692 55748 13694
rect 56252 15820 56308 15876
rect 55916 15314 55972 15316
rect 55916 15262 55918 15314
rect 55918 15262 55970 15314
rect 55970 15262 55972 15314
rect 55916 15260 55972 15262
rect 56700 18508 56756 18564
rect 56476 17500 56532 17556
rect 57372 23324 57428 23380
rect 57708 23324 57764 23380
rect 57372 22764 57428 22820
rect 57484 23100 57540 23156
rect 57260 21532 57316 21588
rect 57596 21532 57652 21588
rect 57708 20972 57764 21028
rect 57372 20802 57428 20804
rect 57372 20750 57374 20802
rect 57374 20750 57426 20802
rect 57426 20750 57428 20802
rect 57372 20748 57428 20750
rect 57484 20130 57540 20132
rect 57484 20078 57486 20130
rect 57486 20078 57538 20130
rect 57538 20078 57540 20130
rect 57484 20076 57540 20078
rect 57820 20914 57876 20916
rect 57820 20862 57822 20914
rect 57822 20862 57874 20914
rect 57874 20862 57876 20914
rect 57820 20860 57876 20862
rect 57932 20524 57988 20580
rect 58044 23996 58100 24052
rect 57260 19122 57316 19124
rect 57260 19070 57262 19122
rect 57262 19070 57314 19122
rect 57314 19070 57316 19122
rect 57260 19068 57316 19070
rect 58044 20076 58100 20132
rect 57820 18674 57876 18676
rect 57820 18622 57822 18674
rect 57822 18622 57874 18674
rect 57874 18622 57876 18674
rect 57820 18620 57876 18622
rect 57708 18508 57764 18564
rect 57484 18172 57540 18228
rect 57372 17612 57428 17668
rect 56588 15538 56644 15540
rect 56588 15486 56590 15538
rect 56590 15486 56642 15538
rect 56642 15486 56644 15538
rect 56588 15484 56644 15486
rect 56364 15260 56420 15316
rect 57708 17442 57764 17444
rect 57708 17390 57710 17442
rect 57710 17390 57762 17442
rect 57762 17390 57764 17442
rect 57708 17388 57764 17390
rect 57484 16994 57540 16996
rect 57484 16942 57486 16994
rect 57486 16942 57538 16994
rect 57538 16942 57540 16994
rect 57484 16940 57540 16942
rect 57372 16268 57428 16324
rect 56924 15874 56980 15876
rect 56924 15822 56926 15874
rect 56926 15822 56978 15874
rect 56978 15822 56980 15874
rect 56924 15820 56980 15822
rect 56140 14476 56196 14532
rect 57260 15260 57316 15316
rect 56028 14252 56084 14308
rect 56364 13916 56420 13972
rect 56140 13804 56196 13860
rect 55580 13522 55636 13524
rect 55580 13470 55582 13522
rect 55582 13470 55634 13522
rect 55634 13470 55636 13522
rect 55580 13468 55636 13470
rect 55580 13244 55636 13300
rect 55916 13132 55972 13188
rect 54796 11340 54852 11396
rect 55804 13020 55860 13076
rect 54908 11170 54964 11172
rect 54908 11118 54910 11170
rect 54910 11118 54962 11170
rect 54962 11118 54964 11170
rect 54908 11116 54964 11118
rect 54908 10444 54964 10500
rect 55692 12012 55748 12068
rect 55356 11564 55412 11620
rect 55356 10834 55412 10836
rect 55356 10782 55358 10834
rect 55358 10782 55410 10834
rect 55410 10782 55412 10834
rect 55356 10780 55412 10782
rect 55580 9938 55636 9940
rect 55580 9886 55582 9938
rect 55582 9886 55634 9938
rect 55634 9886 55636 9938
rect 55580 9884 55636 9886
rect 54684 9436 54740 9492
rect 54684 8316 54740 8372
rect 55468 9324 55524 9380
rect 54796 7980 54852 8036
rect 54460 6748 54516 6804
rect 54124 6636 54180 6692
rect 54908 6690 54964 6692
rect 54908 6638 54910 6690
rect 54910 6638 54962 6690
rect 54962 6638 54964 6690
rect 54908 6636 54964 6638
rect 54236 6524 54292 6580
rect 54460 6578 54516 6580
rect 54460 6526 54462 6578
rect 54462 6526 54514 6578
rect 54514 6526 54516 6578
rect 54460 6524 54516 6526
rect 55020 6412 55076 6468
rect 55132 8316 55188 8372
rect 54684 6130 54740 6132
rect 54684 6078 54686 6130
rect 54686 6078 54738 6130
rect 54738 6078 54740 6130
rect 54684 6076 54740 6078
rect 55356 8092 55412 8148
rect 55244 7586 55300 7588
rect 55244 7534 55246 7586
rect 55246 7534 55298 7586
rect 55298 7534 55300 7586
rect 55244 7532 55300 7534
rect 55356 6578 55412 6580
rect 55356 6526 55358 6578
rect 55358 6526 55410 6578
rect 55410 6526 55412 6578
rect 55356 6524 55412 6526
rect 54572 5292 54628 5348
rect 54124 4226 54180 4228
rect 54124 4174 54126 4226
rect 54126 4174 54178 4226
rect 54178 4174 54180 4226
rect 54124 4172 54180 4174
rect 54908 4172 54964 4228
rect 55244 3666 55300 3668
rect 55244 3614 55246 3666
rect 55246 3614 55298 3666
rect 55298 3614 55300 3666
rect 55244 3612 55300 3614
rect 55356 2716 55412 2772
rect 56252 11506 56308 11508
rect 56252 11454 56254 11506
rect 56254 11454 56306 11506
rect 56306 11454 56308 11506
rect 56252 11452 56308 11454
rect 57036 14812 57092 14868
rect 56700 14418 56756 14420
rect 56700 14366 56702 14418
rect 56702 14366 56754 14418
rect 56754 14366 56756 14418
rect 56700 14364 56756 14366
rect 56588 12402 56644 12404
rect 56588 12350 56590 12402
rect 56590 12350 56642 12402
rect 56642 12350 56644 12402
rect 56588 12348 56644 12350
rect 57148 14588 57204 14644
rect 57036 12850 57092 12852
rect 57036 12798 57038 12850
rect 57038 12798 57090 12850
rect 57090 12798 57092 12850
rect 57036 12796 57092 12798
rect 56924 11676 56980 11732
rect 57484 15820 57540 15876
rect 57820 15708 57876 15764
rect 57932 15820 57988 15876
rect 57708 15314 57764 15316
rect 57708 15262 57710 15314
rect 57710 15262 57762 15314
rect 57762 15262 57764 15314
rect 57708 15260 57764 15262
rect 57708 14924 57764 14980
rect 57596 14476 57652 14532
rect 56700 11394 56756 11396
rect 56700 11342 56702 11394
rect 56702 11342 56754 11394
rect 56754 11342 56756 11394
rect 56700 11340 56756 11342
rect 56476 11004 56532 11060
rect 56588 10556 56644 10612
rect 56476 10498 56532 10500
rect 56476 10446 56478 10498
rect 56478 10446 56530 10498
rect 56530 10446 56532 10498
rect 56476 10444 56532 10446
rect 56252 9938 56308 9940
rect 56252 9886 56254 9938
rect 56254 9886 56306 9938
rect 56306 9886 56308 9938
rect 56252 9884 56308 9886
rect 55916 9212 55972 9268
rect 56140 9266 56196 9268
rect 56140 9214 56142 9266
rect 56142 9214 56194 9266
rect 56194 9214 56196 9266
rect 56140 9212 56196 9214
rect 57148 11788 57204 11844
rect 56700 9324 56756 9380
rect 56140 8652 56196 8708
rect 56252 8316 56308 8372
rect 55692 7196 55748 7252
rect 55580 6748 55636 6804
rect 56588 8370 56644 8372
rect 56588 8318 56590 8370
rect 56590 8318 56642 8370
rect 56642 8318 56644 8370
rect 56588 8316 56644 8318
rect 56588 7698 56644 7700
rect 56588 7646 56590 7698
rect 56590 7646 56642 7698
rect 56642 7646 56644 7698
rect 56588 7644 56644 7646
rect 57372 12402 57428 12404
rect 57372 12350 57374 12402
rect 57374 12350 57426 12402
rect 57426 12350 57428 12402
rect 57372 12348 57428 12350
rect 57820 13074 57876 13076
rect 57820 13022 57822 13074
rect 57822 13022 57874 13074
rect 57874 13022 57876 13074
rect 57820 13020 57876 13022
rect 57932 12796 57988 12852
rect 57372 11452 57428 11508
rect 57596 11506 57652 11508
rect 57596 11454 57598 11506
rect 57598 11454 57650 11506
rect 57650 11454 57652 11506
rect 57596 11452 57652 11454
rect 57372 11228 57428 11284
rect 57372 10444 57428 10500
rect 57484 11340 57540 11396
rect 57260 9996 57316 10052
rect 57260 8764 57316 8820
rect 56700 7308 56756 7364
rect 55804 6690 55860 6692
rect 55804 6638 55806 6690
rect 55806 6638 55858 6690
rect 55858 6638 55860 6690
rect 55804 6636 55860 6638
rect 56700 6690 56756 6692
rect 56700 6638 56702 6690
rect 56702 6638 56754 6690
rect 56754 6638 56756 6690
rect 56700 6636 56756 6638
rect 58044 9938 58100 9940
rect 58044 9886 58046 9938
rect 58046 9886 58098 9938
rect 58098 9886 58100 9938
rect 58044 9884 58100 9886
rect 57484 8652 57540 8708
rect 57708 8540 57764 8596
rect 57596 8034 57652 8036
rect 57596 7982 57598 8034
rect 57598 7982 57650 8034
rect 57650 7982 57652 8034
rect 57596 7980 57652 7982
rect 57484 7644 57540 7700
rect 57372 6636 57428 6692
rect 56476 6130 56532 6132
rect 56476 6078 56478 6130
rect 56478 6078 56530 6130
rect 56530 6078 56532 6130
rect 56476 6076 56532 6078
rect 57596 6466 57652 6468
rect 57596 6414 57598 6466
rect 57598 6414 57650 6466
rect 57650 6414 57652 6466
rect 57596 6412 57652 6414
rect 55916 5794 55972 5796
rect 55916 5742 55918 5794
rect 55918 5742 55970 5794
rect 55970 5742 55972 5794
rect 55916 5740 55972 5742
rect 57148 5628 57204 5684
rect 56700 5234 56756 5236
rect 56700 5182 56702 5234
rect 56702 5182 56754 5234
rect 56754 5182 56756 5234
rect 56700 5180 56756 5182
rect 57820 7362 57876 7364
rect 57820 7310 57822 7362
rect 57822 7310 57874 7362
rect 57874 7310 57876 7362
rect 57820 7308 57876 7310
rect 58044 6860 58100 6916
rect 57820 6412 57876 6468
rect 56252 5010 56308 5012
rect 56252 4958 56254 5010
rect 56254 4958 56306 5010
rect 56306 4958 56308 5010
rect 56252 4956 56308 4958
rect 56140 4396 56196 4452
rect 57484 4450 57540 4452
rect 57484 4398 57486 4450
rect 57486 4398 57538 4450
rect 57538 4398 57540 4450
rect 57484 4396 57540 4398
rect 56588 4060 56644 4116
rect 56700 4172 56756 4228
rect 57484 3948 57540 4004
rect 57148 3612 57204 3668
rect 56252 2828 56308 2884
rect 55468 1596 55524 1652
rect 53900 1484 53956 1540
rect 57708 3276 57764 3332
rect 58044 4898 58100 4900
rect 58044 4846 58046 4898
rect 58046 4846 58098 4898
rect 58098 4846 58100 4898
rect 58044 4844 58100 4846
rect 57932 3724 57988 3780
rect 58268 34748 58324 34804
rect 58268 20972 58324 21028
rect 58268 16716 58324 16772
rect 58268 16156 58324 16212
rect 58604 38444 58660 38500
rect 58716 41804 58772 41860
rect 58716 37548 58772 37604
rect 58716 33180 58772 33236
rect 58492 31388 58548 31444
rect 58716 32508 58772 32564
rect 58492 27916 58548 27972
rect 58604 25282 58660 25284
rect 58604 25230 58606 25282
rect 58606 25230 58658 25282
rect 58658 25230 58660 25282
rect 58604 25228 58660 25230
rect 58492 16716 58548 16772
rect 58604 20972 58660 21028
rect 58380 14252 58436 14308
rect 58492 16492 58548 16548
rect 58380 12796 58436 12852
rect 58492 12348 58548 12404
rect 58380 5628 58436 5684
rect 58940 42476 58996 42532
rect 58940 34636 58996 34692
rect 58828 29484 58884 29540
rect 59500 29484 59556 29540
rect 59164 29372 59220 29428
rect 59052 28700 59108 28756
rect 58940 25900 58996 25956
rect 58716 20076 58772 20132
rect 58828 22988 58884 23044
rect 58828 18844 58884 18900
rect 58716 18172 58772 18228
rect 58828 16492 58884 16548
rect 58716 10780 58772 10836
rect 58828 14812 58884 14868
rect 59052 21980 59108 22036
rect 59276 23660 59332 23716
rect 59052 20412 59108 20468
rect 59052 13020 59108 13076
rect 59164 18956 59220 19012
rect 58940 11452 58996 11508
rect 59276 14812 59332 14868
rect 59500 13468 59556 13524
rect 59164 9884 59220 9940
rect 58828 7980 58884 8036
rect 59612 7868 59668 7924
rect 58604 4956 58660 5012
rect 58268 3276 58324 3332
rect 57820 2604 57876 2660
<< metal3 >>
rect 200 57204 800 57232
rect 200 57148 1932 57204
rect 1988 57148 1998 57204
rect 200 57120 800 57148
rect 43026 57036 43036 57092
rect 43092 57036 43596 57092
rect 43652 57036 43662 57092
rect 19826 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20110 56476
rect 50546 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50830 56476
rect 4162 56252 4172 56308
rect 4228 56252 4732 56308
rect 4788 56252 33628 56308
rect 33684 56252 33694 56308
rect 29922 56140 29932 56196
rect 29988 56140 54236 56196
rect 54292 56140 54684 56196
rect 54740 56140 54750 56196
rect 57810 56140 57820 56196
rect 57876 56140 59836 56196
rect 59892 56140 59902 56196
rect 14130 56028 14140 56084
rect 14196 56028 15148 56084
rect 15204 56028 15214 56084
rect 40002 56028 40012 56084
rect 40068 56028 41244 56084
rect 41300 56028 41310 56084
rect 46946 56028 46956 56084
rect 47012 56028 48860 56084
rect 48916 56028 48926 56084
rect 10098 55916 10108 55972
rect 10164 55916 13916 55972
rect 13972 55916 14364 55972
rect 14420 55916 14430 55972
rect 27010 55916 27020 55972
rect 27076 55916 27580 55972
rect 27636 55916 27692 55972
rect 27748 55916 27758 55972
rect 36866 55916 36876 55972
rect 36932 55916 42476 55972
rect 42532 55916 42924 55972
rect 42980 55916 42990 55972
rect 48402 55916 48412 55972
rect 48468 55916 49532 55972
rect 49588 55916 49598 55972
rect 54450 55916 54460 55972
rect 54516 55916 55468 55972
rect 55524 55916 55534 55972
rect 23650 55804 23660 55860
rect 23716 55804 36428 55860
rect 36484 55804 37212 55860
rect 37268 55804 37278 55860
rect 4466 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4750 55692
rect 35186 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35470 55692
rect 41234 55580 41244 55636
rect 41300 55580 49308 55636
rect 49364 55580 49374 55636
rect 31042 55468 31052 55524
rect 31108 55468 52332 55524
rect 52388 55468 52398 55524
rect 27122 55244 27132 55300
rect 27188 55244 36876 55300
rect 36932 55244 36942 55300
rect 41122 55244 41132 55300
rect 41188 55244 43708 55300
rect 43764 55244 43774 55300
rect 54338 55244 54348 55300
rect 54404 55244 55132 55300
rect 55188 55244 56924 55300
rect 56980 55244 56990 55300
rect 33618 55132 33628 55188
rect 33684 55132 37548 55188
rect 37604 55132 37614 55188
rect 44146 55132 44156 55188
rect 44212 55132 46620 55188
rect 46676 55132 46686 55188
rect 3042 55020 3052 55076
rect 3108 55020 3500 55076
rect 3556 55020 4060 55076
rect 4116 55020 4126 55076
rect 13570 55020 13580 55076
rect 13636 55020 22876 55076
rect 22932 55020 23324 55076
rect 23380 55020 23390 55076
rect 19826 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20110 54908
rect 50546 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50830 54908
rect 42130 54572 42140 54628
rect 42196 54572 43708 54628
rect 43764 54572 43774 54628
rect 59200 54516 59800 54544
rect 38210 54460 38220 54516
rect 38276 54460 39116 54516
rect 39172 54460 39182 54516
rect 40786 54460 40796 54516
rect 40852 54460 41580 54516
rect 41636 54460 43260 54516
rect 43316 54460 43326 54516
rect 56018 54460 56028 54516
rect 56084 54460 59800 54516
rect 59200 54432 59800 54460
rect 38434 54348 38444 54404
rect 38500 54348 39004 54404
rect 39060 54348 39340 54404
rect 39396 54348 39406 54404
rect 40450 54348 40460 54404
rect 40516 54348 42252 54404
rect 42308 54348 42318 54404
rect 42466 54348 42476 54404
rect 42532 54348 43148 54404
rect 43204 54348 43820 54404
rect 43876 54348 43886 54404
rect 42700 54292 42756 54348
rect 42690 54236 42700 54292
rect 42756 54236 42766 54292
rect 4466 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4750 54124
rect 35186 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35470 54124
rect 31892 53788 39228 53844
rect 39284 53788 39294 53844
rect 41570 53788 41580 53844
rect 41636 53788 42812 53844
rect 42868 53788 42878 53844
rect 56578 53788 56588 53844
rect 56644 53788 57148 53844
rect 57204 53788 57214 53844
rect 31892 53620 31948 53788
rect 39330 53676 39340 53732
rect 39396 53676 40348 53732
rect 40404 53676 40414 53732
rect 42914 53676 42924 53732
rect 42980 53676 43932 53732
rect 43988 53676 43998 53732
rect 2706 53564 2716 53620
rect 2772 53564 3164 53620
rect 3220 53564 31948 53620
rect 35970 53564 35980 53620
rect 36036 53564 40460 53620
rect 40516 53564 40526 53620
rect 43586 53452 43596 53508
rect 43652 53452 44380 53508
rect 44436 53452 45388 53508
rect 45444 53452 45454 53508
rect 42466 53340 42476 53396
rect 42532 53340 43820 53396
rect 43876 53340 43886 53396
rect 19826 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20110 53340
rect 50546 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50830 53340
rect 28018 53228 28028 53284
rect 28084 53228 29596 53284
rect 29652 53228 29662 53284
rect 43362 53228 43372 53284
rect 43428 53228 43932 53284
rect 43988 53228 43998 53284
rect 35074 53116 35084 53172
rect 35140 53116 35980 53172
rect 36036 53116 36046 53172
rect 40898 53116 40908 53172
rect 40964 53116 42588 53172
rect 42644 53116 42654 53172
rect 44370 53116 44380 53172
rect 44436 53116 47068 53172
rect 47124 53116 47134 53172
rect 32274 52780 32284 52836
rect 32340 52780 33740 52836
rect 33796 52780 33806 52836
rect 34738 52780 34748 52836
rect 34804 52780 34972 52836
rect 35028 52780 35644 52836
rect 35700 52780 42700 52836
rect 42756 52780 42766 52836
rect 34290 52668 34300 52724
rect 34356 52668 37716 52724
rect 37874 52668 37884 52724
rect 37940 52668 39788 52724
rect 39844 52668 39854 52724
rect 37660 52612 37716 52668
rect 37660 52556 40908 52612
rect 40964 52556 42028 52612
rect 42084 52556 42094 52612
rect 4466 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4750 52556
rect 35186 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35470 52556
rect 32722 52332 32732 52388
rect 32788 52332 34860 52388
rect 34916 52332 34926 52388
rect 42018 52332 42028 52388
rect 42084 52332 42420 52388
rect 42802 52332 42812 52388
rect 42868 52332 43036 52388
rect 43092 52332 45948 52388
rect 46004 52332 46014 52388
rect 42364 52276 42420 52332
rect 33842 52220 33852 52276
rect 33908 52220 34972 52276
rect 35028 52220 35038 52276
rect 36306 52220 36316 52276
rect 36372 52220 36652 52276
rect 36708 52220 37996 52276
rect 38052 52220 38332 52276
rect 38388 52220 40460 52276
rect 40516 52220 42140 52276
rect 42196 52220 42206 52276
rect 42364 52220 43708 52276
rect 43764 52220 43774 52276
rect 44146 52220 44156 52276
rect 44212 52220 47068 52276
rect 47124 52220 47134 52276
rect 49298 52220 49308 52276
rect 49364 52220 50876 52276
rect 50932 52220 50942 52276
rect 33170 52108 33180 52164
rect 33236 52108 33964 52164
rect 34020 52108 34188 52164
rect 34244 52108 34254 52164
rect 38098 52108 38108 52164
rect 38164 52108 39116 52164
rect 39172 52108 39182 52164
rect 42242 52108 42252 52164
rect 42308 52108 43932 52164
rect 43988 52108 43998 52164
rect 33618 51996 33628 52052
rect 33684 51996 34524 52052
rect 34580 51996 34590 52052
rect 35858 51996 35868 52052
rect 35924 51996 36540 52052
rect 36596 51996 36606 52052
rect 40338 51996 40348 52052
rect 40404 51996 41468 52052
rect 41524 51996 41534 52052
rect 46498 51996 46508 52052
rect 46564 51996 47516 52052
rect 47572 51996 47582 52052
rect 47730 51996 47740 52052
rect 47796 51996 49196 52052
rect 49252 51996 49262 52052
rect 47740 51940 47796 51996
rect 31938 51884 31948 51940
rect 32004 51884 36092 51940
rect 36148 51884 37436 51940
rect 37492 51884 38892 51940
rect 38948 51884 41356 51940
rect 41412 51884 42588 51940
rect 42644 51884 42654 51940
rect 46050 51884 46060 51940
rect 46116 51884 47180 51940
rect 47236 51884 47796 51940
rect 200 51828 800 51856
rect 200 51772 1932 51828
rect 1988 51772 1998 51828
rect 47730 51772 47740 51828
rect 47796 51772 48412 51828
rect 48468 51772 48478 51828
rect 200 51744 800 51772
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 45042 51660 45052 51716
rect 45108 51660 47852 51716
rect 47908 51660 47918 51716
rect 37538 51548 37548 51604
rect 37604 51548 38332 51604
rect 38388 51548 38398 51604
rect 38994 51548 39004 51604
rect 39060 51548 43260 51604
rect 43316 51548 43326 51604
rect 46274 51548 46284 51604
rect 46340 51548 46844 51604
rect 46900 51548 47628 51604
rect 47684 51548 49868 51604
rect 49924 51548 49934 51604
rect 38210 51436 38220 51492
rect 38276 51436 41468 51492
rect 41524 51436 43820 51492
rect 43876 51436 43886 51492
rect 46386 51436 46396 51492
rect 46452 51436 47292 51492
rect 47348 51436 48412 51492
rect 48468 51436 48478 51492
rect 24098 51324 24108 51380
rect 24164 51324 24668 51380
rect 24724 51324 24734 51380
rect 31602 51324 31612 51380
rect 31668 51324 32396 51380
rect 32452 51324 32462 51380
rect 34178 51324 34188 51380
rect 34244 51324 35308 51380
rect 35364 51324 35374 51380
rect 36418 51324 36428 51380
rect 36484 51324 37436 51380
rect 37492 51324 40124 51380
rect 40180 51324 40190 51380
rect 41010 51324 41020 51380
rect 41076 51324 44380 51380
rect 44436 51324 44446 51380
rect 29026 51212 29036 51268
rect 29092 51212 34636 51268
rect 34692 51212 34702 51268
rect 38770 51212 38780 51268
rect 38836 51212 39340 51268
rect 39396 51212 40012 51268
rect 40068 51212 42028 51268
rect 42084 51212 42252 51268
rect 42308 51212 42318 51268
rect 24210 51100 24220 51156
rect 24276 51100 26124 51156
rect 26180 51100 28252 51156
rect 28308 51100 28318 51156
rect 42690 50988 42700 51044
rect 42756 50988 45052 51044
rect 45108 50988 45118 51044
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 26114 50876 26124 50932
rect 26180 50876 26460 50932
rect 26516 50876 26796 50932
rect 26852 50876 27468 50932
rect 27524 50876 27534 50932
rect 39778 50876 39788 50932
rect 39844 50876 42476 50932
rect 42532 50876 42542 50932
rect 49522 50876 49532 50932
rect 49588 50876 50204 50932
rect 50260 50876 50270 50932
rect 32722 50764 32732 50820
rect 32788 50764 57932 50820
rect 57988 50764 57998 50820
rect 29474 50652 29484 50708
rect 29540 50652 55356 50708
rect 55412 50652 55422 50708
rect 22754 50540 22764 50596
rect 22820 50540 26348 50596
rect 26404 50540 26414 50596
rect 36082 50540 36092 50596
rect 36148 50540 36158 50596
rect 36754 50540 36764 50596
rect 36820 50540 38220 50596
rect 38276 50540 38286 50596
rect 41122 50540 41132 50596
rect 41188 50540 42700 50596
rect 42756 50540 42766 50596
rect 44034 50540 44044 50596
rect 44100 50540 45388 50596
rect 45444 50540 45454 50596
rect 36092 50484 36148 50540
rect 25218 50428 25228 50484
rect 25284 50428 26124 50484
rect 26180 50428 26190 50484
rect 34738 50428 34748 50484
rect 34804 50428 35196 50484
rect 35252 50428 36372 50484
rect 38658 50428 38668 50484
rect 38724 50428 39228 50484
rect 39284 50428 41020 50484
rect 41076 50428 41086 50484
rect 43250 50428 43260 50484
rect 43316 50428 44716 50484
rect 44772 50428 45724 50484
rect 45780 50428 45790 50484
rect 47170 50428 47180 50484
rect 47236 50428 48076 50484
rect 48132 50428 48142 50484
rect 36316 50372 36372 50428
rect 23650 50316 23660 50372
rect 23716 50316 23996 50372
rect 24052 50316 24062 50372
rect 31154 50316 31164 50372
rect 31220 50316 31836 50372
rect 31892 50316 31902 50372
rect 32498 50316 32508 50372
rect 32564 50316 33516 50372
rect 33572 50316 33582 50372
rect 36306 50316 36316 50372
rect 36372 50316 36382 50372
rect 38994 50316 39004 50372
rect 39060 50316 39788 50372
rect 39844 50316 39854 50372
rect 39666 50204 39676 50260
rect 39732 50204 39900 50260
rect 39956 50204 39966 50260
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 43586 49980 43596 50036
rect 43652 49980 45612 50036
rect 45668 49980 45678 50036
rect 46498 49980 46508 50036
rect 46564 49980 46844 50036
rect 46900 49980 47516 50036
rect 47572 49980 49420 50036
rect 49476 49980 49486 50036
rect 49746 49980 49756 50036
rect 49812 49980 51660 50036
rect 51716 49980 51726 50036
rect 3266 49868 3276 49924
rect 3332 49868 23716 49924
rect 24994 49868 25004 49924
rect 25060 49868 26796 49924
rect 26852 49868 26862 49924
rect 27010 49868 27020 49924
rect 27076 49868 28140 49924
rect 28196 49868 28206 49924
rect 30034 49868 30044 49924
rect 30100 49868 33740 49924
rect 33796 49868 33806 49924
rect 34738 49868 34748 49924
rect 34804 49868 40684 49924
rect 40740 49868 50988 49924
rect 51044 49868 51054 49924
rect 51314 49868 51324 49924
rect 51380 49868 53228 49924
rect 53284 49868 53294 49924
rect 23660 49812 23716 49868
rect 27020 49812 27076 49868
rect 21522 49756 21532 49812
rect 21588 49756 22204 49812
rect 22260 49756 22270 49812
rect 22418 49756 22428 49812
rect 22484 49756 23436 49812
rect 23492 49756 23502 49812
rect 23660 49756 26124 49812
rect 26180 49756 26190 49812
rect 26562 49756 26572 49812
rect 26628 49756 27076 49812
rect 47506 49756 47516 49812
rect 47572 49756 47852 49812
rect 47908 49756 47918 49812
rect 17602 49644 17612 49700
rect 17668 49644 19964 49700
rect 20020 49644 20636 49700
rect 20692 49644 20702 49700
rect 26674 49644 26684 49700
rect 26740 49644 27692 49700
rect 27748 49644 27758 49700
rect 32162 49644 32172 49700
rect 32228 49644 33068 49700
rect 33124 49644 33134 49700
rect 37650 49644 37660 49700
rect 37716 49644 38892 49700
rect 38948 49644 39340 49700
rect 39396 49644 39900 49700
rect 39956 49644 40460 49700
rect 40516 49644 40526 49700
rect 43362 49644 43372 49700
rect 43428 49644 44604 49700
rect 44660 49644 45052 49700
rect 45108 49644 45118 49700
rect 46834 49644 46844 49700
rect 46900 49644 47404 49700
rect 47460 49644 48524 49700
rect 48580 49644 48590 49700
rect 51986 49644 51996 49700
rect 52052 49644 52444 49700
rect 52500 49644 52892 49700
rect 52948 49644 57036 49700
rect 57092 49644 57102 49700
rect 9538 49532 9548 49588
rect 9604 49532 10108 49588
rect 10164 49532 10174 49588
rect 13234 49532 13244 49588
rect 13300 49532 13692 49588
rect 13748 49532 13758 49588
rect 23426 49532 23436 49588
rect 23492 49532 24668 49588
rect 24724 49532 24734 49588
rect 34066 49532 34076 49588
rect 34132 49532 35644 49588
rect 35700 49532 35710 49588
rect 49970 49532 49980 49588
rect 50036 49532 52220 49588
rect 52276 49532 52286 49588
rect 43922 49420 43932 49476
rect 43988 49420 45836 49476
rect 45892 49420 52668 49476
rect 52724 49420 52734 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 13458 49308 13468 49364
rect 13524 49308 13916 49364
rect 13972 49308 14476 49364
rect 14532 49308 14542 49364
rect 40002 49308 40012 49364
rect 40068 49308 40460 49364
rect 40516 49308 40526 49364
rect 48626 49308 48636 49364
rect 48692 49308 49532 49364
rect 49588 49308 51996 49364
rect 52052 49308 52062 49364
rect 9762 49196 9772 49252
rect 9828 49196 15820 49252
rect 15876 49196 17052 49252
rect 17108 49196 17118 49252
rect 32722 49196 32732 49252
rect 32788 49196 34188 49252
rect 34244 49196 34254 49252
rect 34412 49196 48188 49252
rect 48244 49196 48254 49252
rect 34412 49140 34468 49196
rect 12572 49084 13692 49140
rect 13748 49084 13758 49140
rect 21746 49084 21756 49140
rect 21812 49084 23660 49140
rect 23716 49084 23996 49140
rect 24052 49084 24062 49140
rect 26786 49084 26796 49140
rect 26852 49084 27916 49140
rect 27972 49084 27982 49140
rect 30258 49084 30268 49140
rect 30324 49084 31276 49140
rect 31332 49084 31342 49140
rect 31490 49084 31500 49140
rect 31556 49084 34468 49140
rect 36092 49084 46396 49140
rect 46452 49084 46462 49140
rect 46946 49084 46956 49140
rect 47012 49084 47740 49140
rect 47796 49084 47806 49140
rect 12572 49028 12628 49084
rect 31500 49028 31556 49084
rect 12562 48972 12572 49028
rect 12628 48972 12638 49028
rect 12786 48972 12796 49028
rect 12852 48972 16044 49028
rect 16100 48972 16940 49028
rect 16996 48972 17006 49028
rect 20850 48972 20860 49028
rect 20916 48972 21644 49028
rect 21700 48972 21710 49028
rect 30594 48972 30604 49028
rect 30660 48972 31556 49028
rect 31612 48972 32396 49028
rect 32452 48972 33628 49028
rect 33684 48972 33694 49028
rect 34514 48972 34524 49028
rect 34580 48972 35084 49028
rect 35140 48972 35150 49028
rect 31612 48916 31668 48972
rect 10322 48860 10332 48916
rect 10388 48860 11452 48916
rect 11508 48860 12684 48916
rect 12740 48860 12750 48916
rect 29586 48860 29596 48916
rect 29652 48860 30044 48916
rect 30100 48860 30492 48916
rect 30548 48860 31276 48916
rect 31332 48860 31342 48916
rect 31602 48860 31612 48916
rect 31668 48860 31678 48916
rect 33730 48860 33740 48916
rect 33796 48860 35868 48916
rect 35924 48860 35934 48916
rect 36092 48804 36148 49084
rect 37874 48972 37884 49028
rect 37940 48972 39228 49028
rect 39284 48972 39788 49028
rect 39844 48972 39854 49028
rect 40226 48972 40236 49028
rect 40292 48972 40684 49028
rect 40740 48972 40750 49028
rect 46722 48972 46732 49028
rect 46788 48972 47852 49028
rect 47908 48972 49532 49028
rect 49588 48972 49598 49028
rect 40002 48860 40012 48916
rect 40068 48860 41692 48916
rect 41748 48860 41758 48916
rect 42476 48860 45388 48916
rect 45444 48860 46844 48916
rect 46900 48860 46910 48916
rect 47506 48860 47516 48916
rect 47572 48860 48636 48916
rect 48692 48860 50764 48916
rect 50820 48860 50830 48916
rect 42476 48804 42532 48860
rect 12898 48748 12908 48804
rect 12964 48748 13804 48804
rect 13860 48748 13870 48804
rect 24882 48748 24892 48804
rect 24948 48748 26908 48804
rect 26964 48748 26974 48804
rect 31378 48748 31388 48804
rect 31444 48748 32172 48804
rect 32228 48748 32238 48804
rect 33954 48748 33964 48804
rect 34020 48748 35196 48804
rect 35252 48748 35262 48804
rect 35420 48748 36148 48804
rect 39442 48748 39452 48804
rect 39508 48748 42476 48804
rect 42532 48748 42542 48804
rect 43810 48748 43820 48804
rect 43876 48748 44380 48804
rect 44436 48748 46284 48804
rect 46340 48748 48076 48804
rect 48132 48748 48860 48804
rect 48916 48748 48926 48804
rect 53442 48748 53452 48804
rect 53508 48748 54348 48804
rect 54404 48748 55468 48804
rect 55524 48748 55534 48804
rect 34710 48636 34748 48692
rect 34804 48636 34814 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 35420 48580 35476 48748
rect 43586 48636 43596 48692
rect 43652 48636 45500 48692
rect 45556 48636 46060 48692
rect 46116 48636 46126 48692
rect 47404 48636 47628 48692
rect 47684 48636 47694 48692
rect 47404 48580 47460 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 35074 48524 35084 48580
rect 35140 48524 35476 48580
rect 47394 48524 47404 48580
rect 47460 48524 47470 48580
rect 59200 48468 59800 48496
rect 16258 48412 16268 48468
rect 16324 48412 17724 48468
rect 17780 48412 17790 48468
rect 17938 48412 17948 48468
rect 18004 48412 18732 48468
rect 18788 48412 18798 48468
rect 21186 48412 21196 48468
rect 21252 48412 21868 48468
rect 21924 48412 22428 48468
rect 22484 48412 22494 48468
rect 36754 48412 36764 48468
rect 36820 48412 37324 48468
rect 37380 48412 37772 48468
rect 37828 48412 37838 48468
rect 47170 48412 47180 48468
rect 47236 48412 48972 48468
rect 49028 48412 49038 48468
rect 49746 48412 49756 48468
rect 49812 48412 51100 48468
rect 51156 48412 51166 48468
rect 52434 48412 52444 48468
rect 52500 48412 53900 48468
rect 53956 48412 53966 48468
rect 56018 48412 56028 48468
rect 56084 48412 59800 48468
rect 48972 48356 49028 48412
rect 59200 48384 59800 48412
rect 10434 48300 10444 48356
rect 10500 48300 12460 48356
rect 12516 48300 12526 48356
rect 17266 48300 17276 48356
rect 17332 48300 18956 48356
rect 19012 48300 19022 48356
rect 21970 48300 21980 48356
rect 22036 48300 22316 48356
rect 22372 48300 24332 48356
rect 24388 48300 24398 48356
rect 27122 48300 27132 48356
rect 27188 48300 29484 48356
rect 29540 48300 29550 48356
rect 48972 48300 49868 48356
rect 49924 48300 49934 48356
rect 51314 48300 51324 48356
rect 51380 48300 52108 48356
rect 52164 48300 53340 48356
rect 53396 48300 53406 48356
rect 8754 48188 8764 48244
rect 8820 48188 9772 48244
rect 9828 48188 9838 48244
rect 12002 48188 12012 48244
rect 12068 48188 13804 48244
rect 13860 48188 13870 48244
rect 16594 48188 16604 48244
rect 16660 48188 17948 48244
rect 18004 48188 18014 48244
rect 23426 48188 23436 48244
rect 23492 48188 24108 48244
rect 24164 48188 24174 48244
rect 29698 48188 29708 48244
rect 29764 48188 31164 48244
rect 31220 48188 34076 48244
rect 34132 48188 34142 48244
rect 35746 48188 35756 48244
rect 35812 48188 36988 48244
rect 37044 48188 37548 48244
rect 37604 48188 38332 48244
rect 38388 48188 38398 48244
rect 40338 48188 40348 48244
rect 40404 48188 40908 48244
rect 40964 48188 41244 48244
rect 41300 48188 41310 48244
rect 41682 48188 41692 48244
rect 41748 48188 47852 48244
rect 47908 48188 47918 48244
rect 48178 48188 48188 48244
rect 48244 48188 51548 48244
rect 51604 48188 51614 48244
rect 53442 48188 53452 48244
rect 53508 48188 53900 48244
rect 53956 48188 54572 48244
rect 54628 48188 54638 48244
rect 55010 48188 55020 48244
rect 55076 48188 55086 48244
rect 55020 48132 55076 48188
rect 1138 48076 1148 48132
rect 1204 48076 15932 48132
rect 15988 48076 15998 48132
rect 22418 48076 22428 48132
rect 22484 48076 23212 48132
rect 23268 48076 24892 48132
rect 24948 48076 25340 48132
rect 25396 48076 25406 48132
rect 29922 48076 29932 48132
rect 29988 48076 30940 48132
rect 30996 48076 31006 48132
rect 32162 48076 32172 48132
rect 32228 48076 33628 48132
rect 33684 48076 33694 48132
rect 40114 48076 40124 48132
rect 40180 48076 40684 48132
rect 40740 48076 42364 48132
rect 42420 48076 42924 48132
rect 42980 48076 44660 48132
rect 54674 48076 54684 48132
rect 54740 48076 56028 48132
rect 56084 48076 56094 48132
rect 44604 48020 44660 48076
rect 13122 47964 13132 48020
rect 13188 47964 14028 48020
rect 14084 47964 14094 48020
rect 19394 47964 19404 48020
rect 19460 47964 26124 48020
rect 26180 47964 27468 48020
rect 27524 47964 27534 48020
rect 30818 47964 30828 48020
rect 30884 47964 32508 48020
rect 32564 47964 33292 48020
rect 33348 47964 33964 48020
rect 34020 47964 34030 48020
rect 35522 47964 35532 48020
rect 35588 47964 35980 48020
rect 36036 47964 37100 48020
rect 37156 47964 42700 48020
rect 42756 47964 42766 48020
rect 44594 47964 44604 48020
rect 44660 47964 47180 48020
rect 47236 47964 47246 48020
rect 33842 47852 33852 47908
rect 33908 47852 34748 47908
rect 34804 47852 34814 47908
rect 39442 47852 39452 47908
rect 39508 47852 41580 47908
rect 41636 47852 41646 47908
rect 43026 47852 43036 47908
rect 43092 47852 44828 47908
rect 44884 47852 45500 47908
rect 45556 47852 47852 47908
rect 47908 47852 47918 47908
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 19506 47740 19516 47796
rect 19572 47740 24892 47796
rect 24948 47740 25564 47796
rect 25620 47740 25630 47796
rect 33730 47740 33740 47796
rect 33796 47740 34524 47796
rect 34580 47740 34590 47796
rect 36082 47740 36092 47796
rect 36148 47740 36652 47796
rect 36708 47740 43708 47796
rect 43764 47740 43774 47796
rect 51650 47740 51660 47796
rect 51716 47740 53228 47796
rect 53284 47740 54236 47796
rect 54292 47740 57484 47796
rect 57540 47740 57550 47796
rect 7746 47628 7756 47684
rect 7812 47628 8988 47684
rect 9044 47628 10220 47684
rect 10276 47628 10286 47684
rect 32050 47628 32060 47684
rect 32116 47628 38108 47684
rect 38164 47628 38174 47684
rect 40898 47628 40908 47684
rect 40964 47628 42028 47684
rect 42084 47628 44156 47684
rect 44212 47628 45500 47684
rect 45556 47628 45566 47684
rect 53330 47628 53340 47684
rect 53396 47628 55244 47684
rect 55300 47628 56476 47684
rect 56532 47628 56542 47684
rect 11778 47516 11788 47572
rect 11844 47516 12460 47572
rect 12516 47516 12684 47572
rect 12740 47516 13860 47572
rect 18274 47516 18284 47572
rect 18340 47516 19740 47572
rect 19796 47516 19806 47572
rect 34412 47516 34860 47572
rect 34916 47516 46060 47572
rect 46116 47516 46126 47572
rect 51874 47516 51884 47572
rect 51940 47516 53676 47572
rect 53732 47516 53742 47572
rect 13804 47460 13860 47516
rect 7186 47404 7196 47460
rect 7252 47404 8764 47460
rect 8820 47404 8830 47460
rect 10322 47404 10332 47460
rect 10388 47404 10398 47460
rect 11666 47404 11676 47460
rect 11732 47404 12236 47460
rect 12292 47404 12302 47460
rect 13794 47404 13804 47460
rect 13860 47404 13870 47460
rect 14018 47404 14028 47460
rect 14084 47404 15148 47460
rect 15204 47404 15214 47460
rect 21858 47404 21868 47460
rect 21924 47404 23436 47460
rect 23492 47404 23502 47460
rect 23762 47404 23772 47460
rect 23828 47404 26684 47460
rect 26740 47404 26750 47460
rect 10332 47348 10388 47404
rect 12236 47348 12292 47404
rect 34412 47348 34468 47516
rect 38658 47404 38668 47460
rect 38724 47404 39676 47460
rect 39732 47404 41692 47460
rect 41748 47404 41758 47460
rect 42914 47404 42924 47460
rect 42980 47404 44044 47460
rect 44100 47404 44110 47460
rect 51538 47404 51548 47460
rect 51604 47404 53564 47460
rect 53620 47404 53630 47460
rect 54002 47404 54012 47460
rect 54068 47404 54460 47460
rect 54516 47404 54526 47460
rect 10332 47292 11788 47348
rect 11844 47292 11854 47348
rect 12236 47292 13020 47348
rect 13076 47292 13916 47348
rect 13972 47292 13982 47348
rect 22978 47292 22988 47348
rect 23044 47292 23548 47348
rect 23604 47292 24444 47348
rect 24500 47292 24510 47348
rect 30930 47292 30940 47348
rect 30996 47292 32620 47348
rect 32676 47292 32686 47348
rect 33618 47292 33628 47348
rect 33684 47292 34300 47348
rect 34356 47292 34468 47348
rect 35074 47292 35084 47348
rect 35140 47292 37660 47348
rect 37716 47292 37726 47348
rect 38668 47236 38724 47404
rect 50418 47292 50428 47348
rect 50484 47292 51100 47348
rect 51156 47292 51436 47348
rect 51492 47292 51502 47348
rect 52658 47292 52668 47348
rect 52724 47292 53452 47348
rect 53508 47292 54908 47348
rect 54964 47292 54974 47348
rect 9314 47180 9324 47236
rect 9380 47180 9660 47236
rect 9716 47180 10332 47236
rect 10388 47180 10398 47236
rect 17042 47180 17052 47236
rect 17108 47180 18172 47236
rect 18228 47180 18238 47236
rect 28466 47180 28476 47236
rect 28532 47180 30156 47236
rect 30212 47180 30222 47236
rect 37762 47180 37772 47236
rect 37828 47180 38724 47236
rect 51436 47236 51492 47292
rect 51436 47180 52556 47236
rect 52612 47180 52622 47236
rect 54562 47180 54572 47236
rect 54628 47180 55356 47236
rect 55412 47180 55692 47236
rect 55748 47180 55758 47236
rect 14914 47068 14924 47124
rect 14980 47068 15148 47124
rect 15204 47068 18956 47124
rect 19012 47068 19022 47124
rect 35634 47068 35644 47124
rect 35700 47068 35710 47124
rect 40226 47068 40236 47124
rect 40292 47068 40684 47124
rect 40740 47068 40750 47124
rect 41794 47068 41804 47124
rect 41860 47068 42812 47124
rect 42868 47068 44604 47124
rect 44660 47068 44670 47124
rect 49858 47068 49868 47124
rect 49924 47068 50204 47124
rect 50260 47068 50270 47124
rect 52322 47068 52332 47124
rect 52388 47068 56028 47124
rect 56084 47068 56812 47124
rect 56868 47068 56878 47124
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 35644 47012 35700 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 34290 46956 34300 47012
rect 34356 46956 35700 47012
rect 40684 46956 41020 47012
rect 41076 46956 41916 47012
rect 41972 46956 50428 47012
rect 53890 46956 53900 47012
rect 53956 46956 54348 47012
rect 54404 46956 56252 47012
rect 56308 46956 56318 47012
rect 40684 46900 40740 46956
rect 50372 46900 50428 46956
rect 14354 46844 14364 46900
rect 14420 46844 16268 46900
rect 16324 46844 16828 46900
rect 16884 46844 16894 46900
rect 22642 46844 22652 46900
rect 22708 46844 23212 46900
rect 23268 46844 24108 46900
rect 24164 46844 24174 46900
rect 33954 46844 33964 46900
rect 34020 46844 36988 46900
rect 37044 46844 37548 46900
rect 37604 46844 37614 46900
rect 40674 46844 40684 46900
rect 40740 46844 40750 46900
rect 44258 46844 44268 46900
rect 44324 46844 44492 46900
rect 44548 46844 45388 46900
rect 45444 46844 45948 46900
rect 46004 46844 46014 46900
rect 50372 46844 51996 46900
rect 52052 46844 52062 46900
rect 52882 46844 52892 46900
rect 52948 46844 55692 46900
rect 55748 46844 55758 46900
rect 33730 46732 33740 46788
rect 33796 46732 34860 46788
rect 34916 46732 34926 46788
rect 40786 46732 40796 46788
rect 40852 46732 45052 46788
rect 45108 46732 45118 46788
rect 55458 46732 55468 46788
rect 55524 46732 56588 46788
rect 56644 46732 57820 46788
rect 57876 46732 57886 46788
rect 43036 46676 43092 46732
rect 14018 46620 14028 46676
rect 14084 46620 14476 46676
rect 14532 46620 14542 46676
rect 18610 46620 18620 46676
rect 18676 46620 19516 46676
rect 19572 46620 19582 46676
rect 23314 46620 23324 46676
rect 23380 46620 24668 46676
rect 24724 46620 24734 46676
rect 25442 46620 25452 46676
rect 25508 46620 27244 46676
rect 27300 46620 27310 46676
rect 29698 46620 29708 46676
rect 29764 46620 30268 46676
rect 30324 46620 30334 46676
rect 32386 46620 32396 46676
rect 32452 46620 34412 46676
rect 34468 46620 36316 46676
rect 36372 46620 37996 46676
rect 38052 46620 38062 46676
rect 39554 46620 39564 46676
rect 39620 46620 40012 46676
rect 40068 46620 40572 46676
rect 40628 46620 41132 46676
rect 41188 46620 41198 46676
rect 43026 46620 43036 46676
rect 43092 46620 43102 46676
rect 43698 46620 43708 46676
rect 43764 46620 44044 46676
rect 44100 46620 44716 46676
rect 44772 46620 45164 46676
rect 45220 46620 45230 46676
rect 47282 46620 47292 46676
rect 47348 46620 47516 46676
rect 47572 46620 48412 46676
rect 48468 46620 49644 46676
rect 49700 46620 49868 46676
rect 49924 46620 49934 46676
rect 52098 46620 52108 46676
rect 52164 46620 52444 46676
rect 52500 46620 52510 46676
rect 52882 46620 52892 46676
rect 52948 46620 53788 46676
rect 53844 46620 53854 46676
rect 24668 46564 24724 46620
rect 17826 46508 17836 46564
rect 17892 46508 19740 46564
rect 19796 46508 19806 46564
rect 24668 46508 26124 46564
rect 26180 46508 26190 46564
rect 32498 46508 32508 46564
rect 32564 46508 33628 46564
rect 33684 46508 33694 46564
rect 40338 46508 40348 46564
rect 40404 46508 40908 46564
rect 40964 46508 40974 46564
rect 41458 46508 41468 46564
rect 41524 46508 41692 46564
rect 41748 46508 46172 46564
rect 46228 46508 46238 46564
rect 49298 46508 49308 46564
rect 49364 46508 50316 46564
rect 50372 46508 50382 46564
rect 50754 46508 50764 46564
rect 50820 46508 51212 46564
rect 51268 46508 51278 46564
rect 55346 46508 55356 46564
rect 55412 46508 55804 46564
rect 55860 46508 56588 46564
rect 56644 46508 56654 46564
rect 57362 46508 57372 46564
rect 57428 46508 57708 46564
rect 57764 46508 57774 46564
rect 9100 46396 19068 46452
rect 19124 46396 19134 46452
rect 20178 46396 20188 46452
rect 20244 46396 20282 46452
rect 41682 46396 41692 46452
rect 41748 46396 42252 46452
rect 42308 46396 45612 46452
rect 45668 46396 45678 46452
rect 50866 46396 50876 46452
rect 50932 46396 52220 46452
rect 52276 46396 52286 46452
rect 9100 46340 9156 46396
rect 5842 46284 5852 46340
rect 5908 46284 6412 46340
rect 6468 46284 9100 46340
rect 9156 46284 9166 46340
rect 18386 46284 18396 46340
rect 18452 46284 19180 46340
rect 19236 46284 19246 46340
rect 48962 46284 48972 46340
rect 49028 46284 51436 46340
rect 51492 46284 51502 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 10770 46172 10780 46228
rect 10836 46172 25004 46228
rect 25060 46172 25070 46228
rect 28242 46172 28252 46228
rect 28308 46172 29372 46228
rect 29428 46172 29820 46228
rect 29876 46172 29886 46228
rect 47394 46172 47404 46228
rect 47460 46172 50764 46228
rect 50820 46172 50830 46228
rect 3378 46060 3388 46116
rect 3444 46060 31836 46116
rect 31892 46060 31902 46116
rect 37650 46060 37660 46116
rect 37716 46060 38332 46116
rect 38388 46060 40348 46116
rect 40404 46060 40796 46116
rect 40852 46060 40862 46116
rect 50306 46060 50316 46116
rect 50372 46060 50988 46116
rect 51044 46060 51212 46116
rect 51268 46060 57708 46116
rect 57764 46060 57774 46116
rect 24770 45948 24780 46004
rect 24836 45948 26124 46004
rect 26180 45948 26190 46004
rect 27010 45948 27020 46004
rect 27076 45948 57596 46004
rect 57652 45948 57820 46004
rect 57876 45948 57886 46004
rect 3490 45836 3500 45892
rect 3556 45836 8428 45892
rect 23202 45836 23212 45892
rect 23268 45836 24220 45892
rect 24276 45836 24892 45892
rect 24948 45836 24958 45892
rect 28466 45836 28476 45892
rect 28532 45836 29932 45892
rect 29988 45836 29998 45892
rect 37202 45836 37212 45892
rect 37268 45836 37772 45892
rect 37828 45836 38780 45892
rect 38836 45836 39116 45892
rect 39172 45836 39182 45892
rect 39330 45836 39340 45892
rect 39396 45836 40460 45892
rect 40516 45836 41692 45892
rect 41748 45836 41758 45892
rect 43474 45836 43484 45892
rect 43540 45836 44492 45892
rect 44548 45836 44558 45892
rect 44706 45836 44716 45892
rect 44772 45836 48412 45892
rect 48468 45836 48972 45892
rect 49028 45836 49038 45892
rect 50082 45836 50092 45892
rect 50148 45836 55580 45892
rect 55636 45836 55646 45892
rect 200 45780 800 45808
rect 200 45724 1932 45780
rect 1988 45724 1998 45780
rect 200 45696 800 45724
rect 8372 45668 8428 45836
rect 9090 45724 9100 45780
rect 9156 45724 11116 45780
rect 11172 45724 11182 45780
rect 19058 45724 19068 45780
rect 19124 45724 19964 45780
rect 20020 45724 20030 45780
rect 36642 45724 36652 45780
rect 36708 45724 39452 45780
rect 39508 45724 39518 45780
rect 45714 45724 45724 45780
rect 45780 45724 46956 45780
rect 47012 45724 48076 45780
rect 48132 45724 49532 45780
rect 49588 45724 49598 45780
rect 52546 45724 52556 45780
rect 52612 45724 53228 45780
rect 53284 45724 53452 45780
rect 53508 45724 53518 45780
rect 38780 45668 38836 45724
rect 3154 45612 3164 45668
rect 3220 45612 5628 45668
rect 5684 45612 5694 45668
rect 8372 45612 28700 45668
rect 28756 45612 28766 45668
rect 36530 45612 36540 45668
rect 36596 45612 37436 45668
rect 37492 45612 37502 45668
rect 38770 45612 38780 45668
rect 38836 45612 38846 45668
rect 45826 45612 45836 45668
rect 45892 45612 47852 45668
rect 47908 45612 50876 45668
rect 50932 45612 50942 45668
rect 52098 45612 52108 45668
rect 52164 45612 54796 45668
rect 54852 45612 54862 45668
rect 55794 45612 55804 45668
rect 55860 45612 58828 45668
rect 58884 45612 58894 45668
rect 16594 45500 16604 45556
rect 16660 45500 18508 45556
rect 18564 45500 19292 45556
rect 19348 45500 19358 45556
rect 36642 45500 36652 45556
rect 36708 45500 37660 45556
rect 37716 45500 37726 45556
rect 45938 45500 45948 45556
rect 46004 45500 50484 45556
rect 53442 45500 53452 45556
rect 53508 45500 53900 45556
rect 53956 45500 53966 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 24210 45388 24220 45444
rect 24276 45388 27356 45444
rect 27412 45388 27422 45444
rect 33730 45388 33740 45444
rect 33796 45388 34524 45444
rect 34580 45388 35196 45444
rect 35252 45388 38220 45444
rect 38276 45388 49532 45444
rect 49588 45388 49598 45444
rect 50428 45332 50484 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 51426 45388 51436 45444
rect 51492 45388 54012 45444
rect 54068 45388 54460 45444
rect 54516 45388 54526 45444
rect 5730 45276 5740 45332
rect 5796 45276 8428 45332
rect 8484 45276 9772 45332
rect 9828 45276 9838 45332
rect 12674 45276 12684 45332
rect 12740 45276 13132 45332
rect 13188 45276 13580 45332
rect 13636 45276 14028 45332
rect 14084 45276 14700 45332
rect 14756 45276 14766 45332
rect 21410 45276 21420 45332
rect 21476 45276 28140 45332
rect 28196 45276 28206 45332
rect 28914 45276 28924 45332
rect 28980 45276 30268 45332
rect 30324 45276 30716 45332
rect 30772 45276 30782 45332
rect 43810 45276 43820 45332
rect 43876 45276 44156 45332
rect 44212 45276 44222 45332
rect 50418 45276 50428 45332
rect 50484 45276 50494 45332
rect 53778 45276 53788 45332
rect 53844 45276 54908 45332
rect 54964 45276 54974 45332
rect 2706 45164 2716 45220
rect 2772 45164 3276 45220
rect 3332 45164 3342 45220
rect 9650 45164 9660 45220
rect 9716 45164 12012 45220
rect 12068 45164 12572 45220
rect 12628 45164 18564 45220
rect 20962 45164 20972 45220
rect 21028 45164 22988 45220
rect 23044 45164 23054 45220
rect 35522 45164 35532 45220
rect 35588 45164 36428 45220
rect 36484 45164 36494 45220
rect 46050 45164 46060 45220
rect 46116 45164 48076 45220
rect 48132 45164 48748 45220
rect 48804 45164 48814 45220
rect 49970 45164 49980 45220
rect 50036 45164 54012 45220
rect 54068 45164 54078 45220
rect 57474 45164 57484 45220
rect 57540 45164 58044 45220
rect 58100 45164 58110 45220
rect 18508 45108 18564 45164
rect 10098 45052 10108 45108
rect 10164 45052 10556 45108
rect 10612 45052 14588 45108
rect 14644 45052 14654 45108
rect 18498 45052 18508 45108
rect 18564 45052 18732 45108
rect 18788 45052 19964 45108
rect 20020 45052 20030 45108
rect 29922 45052 29932 45108
rect 29988 45052 31724 45108
rect 31780 45052 31790 45108
rect 38546 45052 38556 45108
rect 38612 45052 39564 45108
rect 39620 45052 41132 45108
rect 41188 45052 41804 45108
rect 41860 45052 41870 45108
rect 46386 45052 46396 45108
rect 46452 45052 47964 45108
rect 48020 45052 49084 45108
rect 49140 45052 49150 45108
rect 10658 44940 10668 44996
rect 10724 44940 11564 44996
rect 11620 44940 12796 44996
rect 12852 44940 14028 44996
rect 14084 44940 14252 44996
rect 14308 44940 14318 44996
rect 20290 44940 20300 44996
rect 20356 44940 20524 44996
rect 20580 44940 20860 44996
rect 20916 44940 20926 44996
rect 40898 44940 40908 44996
rect 40964 44940 52332 44996
rect 52388 44940 52398 44996
rect 55570 44940 55580 44996
rect 55636 44940 56364 44996
rect 56420 44940 56430 44996
rect 36194 44828 36204 44884
rect 36260 44828 40684 44884
rect 40740 44828 54460 44884
rect 54516 44828 54526 44884
rect 55458 44828 55468 44884
rect 55524 44828 55580 44884
rect 55636 44828 55646 44884
rect 14690 44716 14700 44772
rect 14756 44716 17948 44772
rect 18004 44716 18014 44772
rect 41234 44716 41244 44772
rect 41300 44716 50204 44772
rect 50260 44716 50270 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 36418 44604 36428 44660
rect 36484 44604 38668 44660
rect 38724 44604 51212 44660
rect 51268 44604 51278 44660
rect 53106 44604 53116 44660
rect 53172 44604 57148 44660
rect 57204 44604 57214 44660
rect 34178 44492 34188 44548
rect 34244 44492 36316 44548
rect 36372 44492 36382 44548
rect 39666 44492 39676 44548
rect 39732 44492 40236 44548
rect 40292 44492 53676 44548
rect 53732 44492 53742 44548
rect 54226 44492 54236 44548
rect 54292 44492 57596 44548
rect 57652 44492 57662 44548
rect 24658 44380 24668 44436
rect 24724 44380 25564 44436
rect 25620 44380 26124 44436
rect 26180 44380 26190 44436
rect 34178 44380 34188 44436
rect 34244 44380 35084 44436
rect 35140 44380 35150 44436
rect 41570 44380 41580 44436
rect 41636 44380 43260 44436
rect 43316 44380 43932 44436
rect 43988 44380 43998 44436
rect 50194 44380 50204 44436
rect 50260 44380 54908 44436
rect 54964 44380 55916 44436
rect 55972 44380 55982 44436
rect 7858 44268 7868 44324
rect 7924 44268 8540 44324
rect 8596 44268 8606 44324
rect 8754 44268 8764 44324
rect 8820 44268 14252 44324
rect 14308 44268 14812 44324
rect 14868 44268 14878 44324
rect 18162 44268 18172 44324
rect 18228 44268 19068 44324
rect 19124 44268 19134 44324
rect 23090 44268 23100 44324
rect 23156 44268 23660 44324
rect 23716 44268 23726 44324
rect 24322 44268 24332 44324
rect 24388 44268 25900 44324
rect 25956 44268 25966 44324
rect 33618 44268 33628 44324
rect 33684 44268 35420 44324
rect 35476 44268 35486 44324
rect 47170 44268 47180 44324
rect 47236 44268 48860 44324
rect 48916 44268 48926 44324
rect 54002 44268 54012 44324
rect 54068 44268 55580 44324
rect 55636 44268 55646 44324
rect 8372 44156 8988 44212
rect 9044 44156 9324 44212
rect 9380 44156 11116 44212
rect 11172 44156 13132 44212
rect 13188 44156 13198 44212
rect 17714 44156 17724 44212
rect 17780 44156 18396 44212
rect 18452 44156 18844 44212
rect 18900 44156 18910 44212
rect 30370 44156 30380 44212
rect 30436 44156 31164 44212
rect 31220 44156 31230 44212
rect 32162 44156 32172 44212
rect 32228 44156 32732 44212
rect 32788 44156 32798 44212
rect 35074 44156 35084 44212
rect 35140 44156 36204 44212
rect 36260 44156 36270 44212
rect 46610 44156 46620 44212
rect 46676 44156 47516 44212
rect 47572 44156 48412 44212
rect 48468 44156 48478 44212
rect 53666 44156 53676 44212
rect 53732 44156 54684 44212
rect 54740 44156 54750 44212
rect 8372 44100 8428 44156
rect 17724 44100 17780 44156
rect 5058 44044 5068 44100
rect 5124 44044 5964 44100
rect 6020 44044 6030 44100
rect 6738 44044 6748 44100
rect 6804 44044 8428 44100
rect 11442 44044 11452 44100
rect 11508 44044 11900 44100
rect 11956 44044 17780 44100
rect 25106 44044 25116 44100
rect 25172 44044 25788 44100
rect 25844 44044 25854 44100
rect 30594 44044 30604 44100
rect 30660 44044 31500 44100
rect 31556 44044 32844 44100
rect 32900 44044 32910 44100
rect 33170 44044 33180 44100
rect 33236 44044 39116 44100
rect 39172 44044 39182 44100
rect 40674 44044 40684 44100
rect 40740 44044 42252 44100
rect 42308 44044 42318 44100
rect 52658 44044 52668 44100
rect 52724 44044 55468 44100
rect 55524 44044 55534 44100
rect 56130 44044 56140 44100
rect 56196 44044 57148 44100
rect 57204 44044 57214 44100
rect 15026 43932 15036 43988
rect 15092 43932 17276 43988
rect 17332 43932 17342 43988
rect 32610 43932 32620 43988
rect 32676 43932 32956 43988
rect 33012 43932 38780 43988
rect 38836 43932 38846 43988
rect 16604 43876 16660 43932
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 13570 43820 13580 43876
rect 13636 43820 13646 43876
rect 16594 43820 16604 43876
rect 16660 43820 16670 43876
rect 18610 43820 18620 43876
rect 18676 43820 18956 43876
rect 19012 43820 19022 43876
rect 36642 43820 36652 43876
rect 36708 43820 42364 43876
rect 42420 43820 44044 43876
rect 44100 43820 44110 43876
rect 46610 43820 46620 43876
rect 46676 43820 47404 43876
rect 47460 43820 47470 43876
rect 51650 43820 51660 43876
rect 51716 43820 51884 43876
rect 51940 43820 53900 43876
rect 53956 43820 53966 43876
rect 13580 43764 13636 43820
rect 13580 43708 14364 43764
rect 14420 43708 15036 43764
rect 15092 43708 15102 43764
rect 22418 43708 22428 43764
rect 22484 43708 23100 43764
rect 23156 43708 23166 43764
rect 37986 43708 37996 43764
rect 38052 43708 38444 43764
rect 38500 43708 39676 43764
rect 39732 43708 39742 43764
rect 40002 43708 40012 43764
rect 40068 43708 41244 43764
rect 41300 43708 41310 43764
rect 41906 43708 41916 43764
rect 41972 43708 42812 43764
rect 42868 43708 42878 43764
rect 48626 43708 48636 43764
rect 48692 43708 50316 43764
rect 50372 43708 50382 43764
rect 50978 43708 50988 43764
rect 51044 43708 51324 43764
rect 51380 43708 51996 43764
rect 52052 43708 52062 43764
rect 56578 43708 56588 43764
rect 56644 43708 58156 43764
rect 58212 43708 58222 43764
rect 5404 43596 8092 43652
rect 8148 43596 8158 43652
rect 10546 43596 10556 43652
rect 10612 43596 11788 43652
rect 11844 43596 11854 43652
rect 17826 43596 17836 43652
rect 17892 43596 18508 43652
rect 18564 43596 18574 43652
rect 34514 43596 34524 43652
rect 34580 43596 35868 43652
rect 35924 43596 35934 43652
rect 41122 43596 41132 43652
rect 41188 43596 41468 43652
rect 41524 43596 41534 43652
rect 44370 43596 44380 43652
rect 44436 43596 44716 43652
rect 44772 43596 46172 43652
rect 46228 43596 46238 43652
rect 46834 43596 46844 43652
rect 46900 43596 48076 43652
rect 48132 43596 48412 43652
rect 48468 43596 49196 43652
rect 49252 43596 50204 43652
rect 50260 43596 50270 43652
rect 50866 43596 50876 43652
rect 50932 43596 51548 43652
rect 51604 43596 51614 43652
rect 52546 43596 52556 43652
rect 52612 43596 55356 43652
rect 55412 43596 55422 43652
rect 5404 43540 5460 43596
rect 2818 43484 2828 43540
rect 2884 43484 5404 43540
rect 5460 43484 5470 43540
rect 6962 43484 6972 43540
rect 7028 43484 10220 43540
rect 10276 43484 10286 43540
rect 11106 43484 11116 43540
rect 11172 43484 12012 43540
rect 12068 43484 12572 43540
rect 12628 43484 12638 43540
rect 15138 43484 15148 43540
rect 15204 43484 15820 43540
rect 15876 43484 16268 43540
rect 16324 43484 16334 43540
rect 20290 43484 20300 43540
rect 20356 43484 21420 43540
rect 21476 43484 21486 43540
rect 23090 43484 23100 43540
rect 23156 43484 24556 43540
rect 24612 43484 25676 43540
rect 25732 43484 25742 43540
rect 29810 43484 29820 43540
rect 29876 43484 31276 43540
rect 31332 43484 31342 43540
rect 31948 43484 32284 43540
rect 32340 43484 32350 43540
rect 40786 43484 40796 43540
rect 40852 43484 43820 43540
rect 43876 43484 43886 43540
rect 45266 43484 45276 43540
rect 45332 43484 45836 43540
rect 45892 43484 45902 43540
rect 46610 43484 46620 43540
rect 46676 43484 48524 43540
rect 48580 43484 48590 43540
rect 49074 43484 49084 43540
rect 49140 43484 49700 43540
rect 50418 43484 50428 43540
rect 50484 43484 51100 43540
rect 51156 43484 51324 43540
rect 51380 43484 51390 43540
rect 53330 43484 53340 43540
rect 53396 43484 53564 43540
rect 53620 43484 55020 43540
rect 55076 43484 55086 43540
rect 31948 43428 32004 43484
rect 45836 43428 45892 43484
rect 49644 43428 49700 43484
rect 6738 43372 6748 43428
rect 6804 43372 7644 43428
rect 7700 43372 7980 43428
rect 8036 43372 8428 43428
rect 8484 43372 8494 43428
rect 10668 43372 14252 43428
rect 14308 43372 14318 43428
rect 31938 43372 31948 43428
rect 32004 43372 32014 43428
rect 35074 43372 35084 43428
rect 35140 43372 37436 43428
rect 37492 43372 37502 43428
rect 39330 43372 39340 43428
rect 39396 43372 40236 43428
rect 40292 43372 40302 43428
rect 41010 43372 41020 43428
rect 41076 43372 42140 43428
rect 42196 43372 42476 43428
rect 42532 43372 42542 43428
rect 43026 43372 43036 43428
rect 43092 43372 44940 43428
rect 44996 43372 45006 43428
rect 45836 43372 48188 43428
rect 48244 43372 49420 43428
rect 49476 43372 49486 43428
rect 49634 43372 49644 43428
rect 49700 43372 52220 43428
rect 52276 43372 52286 43428
rect 53218 43372 53228 43428
rect 53284 43372 53340 43428
rect 53396 43372 53406 43428
rect 56578 43372 56588 43428
rect 56644 43372 56700 43428
rect 56756 43372 56924 43428
rect 56980 43372 57820 43428
rect 57876 43372 57886 43428
rect 10668 43204 10724 43372
rect 8306 43148 8316 43204
rect 8372 43148 10724 43204
rect 10780 43260 20692 43316
rect 20850 43260 20860 43316
rect 20916 43260 23884 43316
rect 23940 43260 23950 43316
rect 31042 43260 31052 43316
rect 31108 43260 31118 43316
rect 32722 43260 32732 43316
rect 32788 43260 33404 43316
rect 33460 43260 33470 43316
rect 38882 43260 38892 43316
rect 38948 43260 39452 43316
rect 39508 43260 40684 43316
rect 40740 43260 41580 43316
rect 41636 43260 41646 43316
rect 49746 43260 49756 43316
rect 49812 43260 52556 43316
rect 52612 43260 52622 43316
rect 53890 43260 53900 43316
rect 53956 43260 55468 43316
rect 55524 43260 56364 43316
rect 56420 43260 56430 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 10780 43092 10836 43260
rect 20636 43204 20692 43260
rect 31052 43204 31108 43260
rect 53900 43204 53956 43260
rect 20636 43148 21196 43204
rect 21252 43148 21262 43204
rect 31052 43148 31276 43204
rect 31332 43148 31342 43204
rect 41654 43148 41692 43204
rect 41748 43148 41758 43204
rect 43334 43148 43372 43204
rect 43428 43148 43438 43204
rect 50306 43148 50316 43204
rect 50372 43148 52108 43204
rect 52164 43148 52174 43204
rect 53666 43148 53676 43204
rect 53732 43148 53956 43204
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 59200 43092 59800 43120
rect 8082 43036 8092 43092
rect 8148 43036 10836 43092
rect 11106 43036 11116 43092
rect 11172 43036 12124 43092
rect 12180 43036 12190 43092
rect 12348 43036 13972 43092
rect 14242 43036 14252 43092
rect 14308 43036 26124 43092
rect 26180 43036 26190 43092
rect 43698 43036 43708 43092
rect 43764 43036 51100 43092
rect 51156 43036 51166 43092
rect 54012 43036 54348 43092
rect 54404 43036 54414 43092
rect 55346 43036 55356 43092
rect 55412 43036 59800 43092
rect 12348 42980 12404 43036
rect 13916 42980 13972 43036
rect 4946 42924 4956 42980
rect 5012 42924 6412 42980
rect 6468 42924 7084 42980
rect 7140 42924 7150 42980
rect 9762 42924 9772 42980
rect 9828 42924 12404 42980
rect 12674 42924 12684 42980
rect 12740 42924 13692 42980
rect 13748 42924 13758 42980
rect 13916 42924 28476 42980
rect 28532 42924 28542 42980
rect 39890 42924 39900 42980
rect 39956 42924 40236 42980
rect 40292 42924 40302 42980
rect 43810 42924 43820 42980
rect 43876 42924 45724 42980
rect 45780 42924 46732 42980
rect 46788 42924 46798 42980
rect 12898 42812 12908 42868
rect 12964 42812 13804 42868
rect 13860 42812 13870 42868
rect 23314 42812 23324 42868
rect 23380 42812 24108 42868
rect 24164 42812 24174 42868
rect 24994 42812 25004 42868
rect 25060 42812 26348 42868
rect 26404 42812 26908 42868
rect 26964 42812 26974 42868
rect 36082 42812 36092 42868
rect 36148 42812 36652 42868
rect 36708 42812 36718 42868
rect 38556 42812 39788 42868
rect 39844 42812 40460 42868
rect 40516 42812 41804 42868
rect 41860 42812 50092 42868
rect 50148 42812 50158 42868
rect 38556 42756 38612 42812
rect 54012 42756 54068 43036
rect 59200 43008 59800 43036
rect 3826 42700 3836 42756
rect 3892 42700 6300 42756
rect 6356 42700 6860 42756
rect 6916 42700 6926 42756
rect 10322 42700 10332 42756
rect 10388 42700 11004 42756
rect 11060 42700 11452 42756
rect 11508 42700 12348 42756
rect 12404 42700 12414 42756
rect 28130 42700 28140 42756
rect 28196 42700 29596 42756
rect 29652 42700 29662 42756
rect 30370 42700 30380 42756
rect 30436 42700 31052 42756
rect 31108 42700 31118 42756
rect 31714 42700 31724 42756
rect 31780 42700 32508 42756
rect 32564 42700 32574 42756
rect 32722 42700 32732 42756
rect 32788 42700 33852 42756
rect 33908 42700 33918 42756
rect 36754 42700 36764 42756
rect 36820 42700 37660 42756
rect 37716 42700 38332 42756
rect 38388 42700 38398 42756
rect 38546 42700 38556 42756
rect 38612 42700 38622 42756
rect 39442 42700 39452 42756
rect 39508 42700 39676 42756
rect 39732 42700 40684 42756
rect 40740 42700 40750 42756
rect 42802 42700 42812 42756
rect 42868 42700 44268 42756
rect 44324 42700 44334 42756
rect 45938 42700 45948 42756
rect 46004 42700 46844 42756
rect 46900 42700 46910 42756
rect 54002 42700 54012 42756
rect 54068 42700 54078 42756
rect 55122 42700 55132 42756
rect 55188 42700 56252 42756
rect 56308 42700 56318 42756
rect 3714 42588 3724 42644
rect 3780 42588 4844 42644
rect 4900 42588 4910 42644
rect 13682 42588 13692 42644
rect 13748 42588 14140 42644
rect 14196 42588 19516 42644
rect 19572 42588 19582 42644
rect 28802 42588 28812 42644
rect 28868 42588 29372 42644
rect 29428 42588 29438 42644
rect 30258 42588 30268 42644
rect 30324 42588 30940 42644
rect 30996 42588 32620 42644
rect 32676 42588 32686 42644
rect 37202 42588 37212 42644
rect 37268 42588 38220 42644
rect 38276 42588 39004 42644
rect 39060 42588 39172 42644
rect 39330 42588 39340 42644
rect 39396 42588 46060 42644
rect 46116 42588 46126 42644
rect 50418 42588 50428 42644
rect 50484 42588 51660 42644
rect 51716 42588 51726 42644
rect 39116 42532 39172 42588
rect 7746 42476 7756 42532
rect 7812 42476 8092 42532
rect 8148 42476 8158 42532
rect 15250 42476 15260 42532
rect 15316 42476 16268 42532
rect 16324 42476 16334 42532
rect 17154 42476 17164 42532
rect 17220 42476 18060 42532
rect 18116 42476 18126 42532
rect 19170 42476 19180 42532
rect 19236 42476 19740 42532
rect 19796 42476 20748 42532
rect 20804 42476 21308 42532
rect 21364 42476 21374 42532
rect 31378 42476 31388 42532
rect 31444 42476 32956 42532
rect 33012 42476 33516 42532
rect 33572 42476 33582 42532
rect 35410 42476 35420 42532
rect 35476 42476 35644 42532
rect 35700 42476 35710 42532
rect 35858 42476 35868 42532
rect 35924 42476 36652 42532
rect 36708 42476 36718 42532
rect 37874 42476 37884 42532
rect 37940 42476 38892 42532
rect 38948 42476 38958 42532
rect 39116 42476 41132 42532
rect 41188 42476 41198 42532
rect 41346 42476 41356 42532
rect 41412 42476 41580 42532
rect 41636 42476 43708 42532
rect 43764 42476 43774 42532
rect 44482 42476 44492 42532
rect 44548 42476 47516 42532
rect 47572 42476 47582 42532
rect 57362 42476 57372 42532
rect 57428 42476 58940 42532
rect 58996 42476 59006 42532
rect 7410 42364 7420 42420
rect 7476 42364 8204 42420
rect 8260 42364 14700 42420
rect 14756 42364 15596 42420
rect 15652 42364 18844 42420
rect 18900 42364 18910 42420
rect 27234 42364 27244 42420
rect 27300 42364 45388 42420
rect 45444 42364 45454 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 3154 42252 3164 42308
rect 3220 42252 17612 42308
rect 17668 42252 17678 42308
rect 34738 42252 34748 42308
rect 34804 42252 36092 42308
rect 36148 42252 36158 42308
rect 36642 42252 36652 42308
rect 36708 42252 38108 42308
rect 38164 42252 38174 42308
rect 39974 42252 40012 42308
rect 40068 42252 40078 42308
rect 42802 42252 42812 42308
rect 42868 42252 45164 42308
rect 45220 42252 45230 42308
rect 12786 42140 12796 42196
rect 12852 42140 13356 42196
rect 13412 42140 13422 42196
rect 20178 42140 20188 42196
rect 20244 42140 22876 42196
rect 22932 42140 24332 42196
rect 24388 42140 24398 42196
rect 25218 42140 25228 42196
rect 25284 42140 26012 42196
rect 26068 42140 26078 42196
rect 31602 42140 31612 42196
rect 31668 42140 36988 42196
rect 37044 42140 37054 42196
rect 38882 42140 38892 42196
rect 38948 42140 41244 42196
rect 41300 42140 41310 42196
rect 41468 42140 45276 42196
rect 45332 42140 49476 42196
rect 53106 42140 53116 42196
rect 53172 42140 54012 42196
rect 54068 42140 54078 42196
rect 41468 42084 41524 42140
rect 49420 42084 49476 42140
rect 13122 42028 13132 42084
rect 13188 42028 13916 42084
rect 13972 42028 14924 42084
rect 14980 42028 14990 42084
rect 16482 42028 16492 42084
rect 16548 42028 17052 42084
rect 17108 42028 23324 42084
rect 23380 42028 23390 42084
rect 28578 42028 28588 42084
rect 28644 42028 29596 42084
rect 29652 42028 30380 42084
rect 30436 42028 30446 42084
rect 31826 42028 31836 42084
rect 31892 42028 34076 42084
rect 34132 42028 34142 42084
rect 35746 42028 35756 42084
rect 35812 42028 35980 42084
rect 36036 42028 40684 42084
rect 40740 42028 41524 42084
rect 42466 42028 42476 42084
rect 42532 42028 44828 42084
rect 44884 42028 44894 42084
rect 47842 42028 47852 42084
rect 47908 42028 48524 42084
rect 48580 42028 48590 42084
rect 49410 42028 49420 42084
rect 49476 42028 50204 42084
rect 50260 42028 50270 42084
rect 51538 42028 51548 42084
rect 51604 42028 51996 42084
rect 52052 42028 52444 42084
rect 52500 42028 52510 42084
rect 55570 42028 55580 42084
rect 55636 42028 56140 42084
rect 56196 42028 56206 42084
rect 5954 41916 5964 41972
rect 6020 41916 6972 41972
rect 7028 41916 7038 41972
rect 8978 41916 8988 41972
rect 9044 41916 9772 41972
rect 9828 41916 9838 41972
rect 15698 41916 15708 41972
rect 15764 41916 16716 41972
rect 16772 41916 18060 41972
rect 18116 41916 18126 41972
rect 33618 41916 33628 41972
rect 33684 41916 35644 41972
rect 35700 41916 35756 41972
rect 35812 41916 35822 41972
rect 37090 41916 37100 41972
rect 37156 41916 37772 41972
rect 37828 41916 37838 41972
rect 38882 41916 38892 41972
rect 38948 41916 39900 41972
rect 39956 41916 39966 41972
rect 40338 41916 40348 41972
rect 40404 41916 45948 41972
rect 46004 41916 46014 41972
rect 50306 41916 50316 41972
rect 50372 41916 50428 41972
rect 50484 41916 50494 41972
rect 51090 41916 51100 41972
rect 51156 41916 55244 41972
rect 55300 41916 55310 41972
rect 5730 41804 5740 41860
rect 5796 41804 6748 41860
rect 6804 41804 6814 41860
rect 9996 41804 10780 41860
rect 10836 41804 19404 41860
rect 19460 41804 19470 41860
rect 34962 41804 34972 41860
rect 35028 41804 41692 41860
rect 41748 41804 41758 41860
rect 42242 41804 42252 41860
rect 42308 41804 43820 41860
rect 43876 41804 44492 41860
rect 44548 41804 45164 41860
rect 45220 41804 45230 41860
rect 51538 41804 51548 41860
rect 51604 41804 52220 41860
rect 52276 41804 52286 41860
rect 56130 41804 56140 41860
rect 56196 41804 57372 41860
rect 57428 41804 57438 41860
rect 57810 41804 57820 41860
rect 57876 41804 58716 41860
rect 58772 41804 58782 41860
rect 9996 41748 10052 41804
rect 3938 41692 3948 41748
rect 4004 41692 5516 41748
rect 5572 41692 7084 41748
rect 7140 41692 7150 41748
rect 9986 41692 9996 41748
rect 10052 41692 10062 41748
rect 16034 41692 16044 41748
rect 16100 41692 18284 41748
rect 18340 41692 18350 41748
rect 20738 41692 20748 41748
rect 20804 41692 25900 41748
rect 25956 41692 25966 41748
rect 34290 41692 34300 41748
rect 34356 41692 35756 41748
rect 35812 41692 35822 41748
rect 45378 41580 45388 41636
rect 45444 41580 54572 41636
rect 54628 41580 54638 41636
rect 55570 41580 55580 41636
rect 55636 41580 56476 41636
rect 56532 41580 56542 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 40226 41468 40236 41524
rect 40292 41468 52332 41524
rect 52388 41468 52398 41524
rect 26002 41356 26012 41412
rect 26068 41356 27244 41412
rect 27300 41356 27310 41412
rect 43026 41356 43036 41412
rect 43092 41356 43596 41412
rect 43652 41356 45612 41412
rect 45668 41356 45678 41412
rect 54114 41356 54124 41412
rect 54180 41356 56812 41412
rect 56868 41356 56878 41412
rect 2930 41244 2940 41300
rect 2996 41244 3724 41300
rect 3780 41244 3790 41300
rect 8372 41244 8988 41300
rect 9044 41244 9054 41300
rect 16594 41244 16604 41300
rect 16660 41244 17836 41300
rect 17892 41244 17902 41300
rect 36866 41244 36876 41300
rect 36932 41244 37884 41300
rect 37940 41244 41020 41300
rect 41076 41244 41086 41300
rect 44034 41244 44044 41300
rect 44100 41244 47068 41300
rect 47124 41244 47134 41300
rect 47730 41244 47740 41300
rect 47796 41244 48524 41300
rect 48580 41244 48590 41300
rect 8372 41188 8428 41244
rect 2594 41132 2604 41188
rect 2660 41132 3276 41188
rect 3332 41132 8428 41188
rect 8530 41132 8540 41188
rect 8596 41132 9436 41188
rect 9492 41132 9884 41188
rect 9940 41132 10220 41188
rect 10276 41132 10286 41188
rect 24994 41132 25004 41188
rect 25060 41132 26684 41188
rect 26740 41132 27804 41188
rect 27860 41132 27870 41188
rect 35410 41132 35420 41188
rect 35476 41132 35644 41188
rect 35700 41132 35710 41188
rect 38098 41132 38108 41188
rect 38164 41132 38892 41188
rect 38948 41132 38958 41188
rect 42690 41132 42700 41188
rect 42756 41132 44380 41188
rect 44436 41132 44446 41188
rect 55122 41132 55132 41188
rect 55188 41132 56140 41188
rect 56196 41132 56206 41188
rect 1026 41020 1036 41076
rect 1092 41020 3052 41076
rect 3108 41020 3118 41076
rect 3490 41020 3500 41076
rect 3556 41020 3724 41076
rect 3780 41020 5740 41076
rect 5796 41020 5806 41076
rect 6290 41020 6300 41076
rect 6356 41020 6860 41076
rect 6916 41020 6926 41076
rect 8194 41020 8204 41076
rect 8260 41020 8988 41076
rect 9044 41020 9548 41076
rect 9604 41020 10668 41076
rect 10724 41020 10734 41076
rect 26338 41020 26348 41076
rect 26404 41020 27356 41076
rect 27412 41020 27422 41076
rect 28690 41020 28700 41076
rect 28756 41020 29932 41076
rect 29988 41020 31500 41076
rect 31556 41020 31566 41076
rect 33842 41020 33852 41076
rect 33908 41020 35532 41076
rect 35588 41020 35598 41076
rect 39106 41020 39116 41076
rect 39172 41020 39676 41076
rect 39732 41020 40124 41076
rect 40180 41020 40190 41076
rect 43250 41020 43260 41076
rect 43316 41020 45388 41076
rect 45444 41020 45454 41076
rect 46834 41020 46844 41076
rect 46900 41020 47740 41076
rect 47796 41020 47806 41076
rect 52098 41020 52108 41076
rect 52164 41020 52444 41076
rect 52500 41020 53788 41076
rect 53844 41020 53854 41076
rect 55234 41020 55244 41076
rect 55300 41020 56252 41076
rect 56308 41020 56318 41076
rect 39116 40964 39172 41020
rect 7970 40908 7980 40964
rect 8036 40908 9660 40964
rect 9716 40908 10780 40964
rect 10836 40908 10846 40964
rect 14690 40908 14700 40964
rect 14756 40908 15148 40964
rect 15204 40908 15820 40964
rect 15876 40908 15886 40964
rect 16044 40908 19628 40964
rect 19684 40908 20860 40964
rect 20916 40908 21644 40964
rect 21700 40908 21710 40964
rect 22194 40908 22204 40964
rect 22260 40908 22988 40964
rect 23044 40908 23054 40964
rect 25890 40908 25900 40964
rect 25956 40908 27244 40964
rect 27300 40908 27310 40964
rect 34066 40908 34076 40964
rect 34132 40908 34748 40964
rect 34804 40908 34814 40964
rect 38322 40908 38332 40964
rect 38388 40908 39172 40964
rect 39554 40908 39564 40964
rect 39620 40908 40012 40964
rect 40068 40908 40078 40964
rect 41570 40908 41580 40964
rect 41636 40908 41916 40964
rect 41972 40908 46396 40964
rect 46452 40908 46462 40964
rect 46722 40908 46732 40964
rect 46788 40908 47404 40964
rect 47460 40908 48076 40964
rect 48132 40908 48142 40964
rect 49858 40908 49868 40964
rect 49924 40908 51548 40964
rect 51604 40908 51772 40964
rect 51828 40908 52668 40964
rect 52724 40908 52734 40964
rect 54338 40908 54348 40964
rect 54404 40908 55468 40964
rect 55524 40908 56364 40964
rect 56420 40908 56430 40964
rect 4946 40796 4956 40852
rect 5012 40796 9996 40852
rect 10052 40796 10062 40852
rect 16044 40740 16100 40908
rect 43586 40796 43596 40852
rect 43652 40796 44940 40852
rect 44996 40796 47516 40852
rect 47572 40796 47582 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 5730 40684 5740 40740
rect 5796 40684 6300 40740
rect 6356 40684 6748 40740
rect 6804 40684 7532 40740
rect 7588 40684 8204 40740
rect 8260 40684 16100 40740
rect 36418 40684 36428 40740
rect 36484 40684 38668 40740
rect 44706 40684 44716 40740
rect 44772 40684 46060 40740
rect 46116 40684 46284 40740
rect 46340 40684 46844 40740
rect 46900 40684 50428 40740
rect 52322 40684 52332 40740
rect 52388 40684 52892 40740
rect 52948 40684 52958 40740
rect 55458 40684 55468 40740
rect 55524 40684 56028 40740
rect 56084 40684 56094 40740
rect 38612 40628 38668 40684
rect 50372 40628 50428 40684
rect 3154 40572 3164 40628
rect 3220 40572 26796 40628
rect 26852 40572 26862 40628
rect 35298 40572 35308 40628
rect 35364 40572 36204 40628
rect 36260 40572 36876 40628
rect 36932 40572 36942 40628
rect 38612 40572 39116 40628
rect 39172 40572 39182 40628
rect 42914 40572 42924 40628
rect 42980 40572 44604 40628
rect 44660 40572 44670 40628
rect 46620 40572 47964 40628
rect 48020 40572 48030 40628
rect 48178 40572 48188 40628
rect 48244 40572 48748 40628
rect 48804 40572 49756 40628
rect 49812 40572 49822 40628
rect 50372 40572 51884 40628
rect 51940 40572 51950 40628
rect 52518 40572 52556 40628
rect 52612 40572 53116 40628
rect 53172 40572 53182 40628
rect 46620 40516 46676 40572
rect 6514 40460 6524 40516
rect 6580 40460 6972 40516
rect 7028 40460 7644 40516
rect 7700 40460 7710 40516
rect 8082 40460 8092 40516
rect 8148 40460 8764 40516
rect 8820 40460 10220 40516
rect 10276 40460 11340 40516
rect 11396 40460 11406 40516
rect 16044 40460 17612 40516
rect 17668 40460 17678 40516
rect 18844 40460 19404 40516
rect 19460 40460 20524 40516
rect 20580 40460 20590 40516
rect 28812 40460 29708 40516
rect 29764 40460 29774 40516
rect 33842 40460 33852 40516
rect 33908 40460 34076 40516
rect 34132 40460 38220 40516
rect 38276 40460 38286 40516
rect 43138 40460 43148 40516
rect 43204 40460 44492 40516
rect 44548 40460 46620 40516
rect 46676 40460 46686 40516
rect 47730 40460 47740 40516
rect 47796 40460 49532 40516
rect 49588 40460 49598 40516
rect 52210 40460 52220 40516
rect 52276 40460 53116 40516
rect 53172 40460 53182 40516
rect 55122 40460 55132 40516
rect 55188 40460 55692 40516
rect 55748 40460 55758 40516
rect 16044 40404 16100 40460
rect 18844 40404 18900 40460
rect 28812 40404 28868 40460
rect 5852 40348 7308 40404
rect 7364 40348 7374 40404
rect 15138 40348 15148 40404
rect 15204 40348 16044 40404
rect 16100 40348 16110 40404
rect 16370 40348 16380 40404
rect 16436 40348 17724 40404
rect 17780 40348 18844 40404
rect 18900 40348 18910 40404
rect 19282 40348 19292 40404
rect 19348 40348 20300 40404
rect 20356 40348 20860 40404
rect 20916 40348 21868 40404
rect 21924 40348 21934 40404
rect 23538 40348 23548 40404
rect 23604 40348 24332 40404
rect 24388 40348 24398 40404
rect 27458 40348 27468 40404
rect 27524 40348 28364 40404
rect 28420 40348 28812 40404
rect 28868 40348 28878 40404
rect 29138 40348 29148 40404
rect 29204 40348 30156 40404
rect 30212 40348 30492 40404
rect 30548 40348 30558 40404
rect 33618 40348 33628 40404
rect 33684 40348 34300 40404
rect 34356 40348 35644 40404
rect 35700 40348 35710 40404
rect 41570 40348 41580 40404
rect 41636 40348 42252 40404
rect 42308 40348 42318 40404
rect 46386 40348 46396 40404
rect 46452 40348 47404 40404
rect 47460 40348 47470 40404
rect 48514 40348 48524 40404
rect 48580 40348 50092 40404
rect 50148 40348 50764 40404
rect 50820 40348 50830 40404
rect 51090 40348 51100 40404
rect 51156 40348 51436 40404
rect 51492 40348 51502 40404
rect 52098 40348 52108 40404
rect 52164 40348 52500 40404
rect 53190 40348 53228 40404
rect 53284 40348 53294 40404
rect 55010 40348 55020 40404
rect 55076 40348 55356 40404
rect 55412 40348 55804 40404
rect 55860 40348 55870 40404
rect 5852 40292 5908 40348
rect 52444 40292 52500 40348
rect 5394 40236 5404 40292
rect 5460 40236 5852 40292
rect 5908 40236 5918 40292
rect 7858 40236 7868 40292
rect 7924 40236 8428 40292
rect 8484 40236 8494 40292
rect 12348 40236 13020 40292
rect 13076 40236 13692 40292
rect 13748 40236 14140 40292
rect 14196 40236 14206 40292
rect 18162 40236 18172 40292
rect 18228 40236 18732 40292
rect 18788 40236 22764 40292
rect 22820 40236 22830 40292
rect 27682 40236 27692 40292
rect 27748 40236 29036 40292
rect 29092 40236 29596 40292
rect 29652 40236 29662 40292
rect 35522 40236 35532 40292
rect 35588 40236 36540 40292
rect 36596 40236 36606 40292
rect 52434 40236 52444 40292
rect 52500 40236 52510 40292
rect 12348 40180 12404 40236
rect 7970 40124 7980 40180
rect 8036 40124 11564 40180
rect 11620 40124 12348 40180
rect 12404 40124 12414 40180
rect 12786 40124 12796 40180
rect 12852 40124 13804 40180
rect 13860 40124 14476 40180
rect 14532 40124 14542 40180
rect 16034 40124 16044 40180
rect 16100 40124 16940 40180
rect 16996 40124 17006 40180
rect 35074 40124 35084 40180
rect 35140 40124 35644 40180
rect 35700 40124 37324 40180
rect 37380 40124 37390 40180
rect 52434 40124 52444 40180
rect 52500 40124 52556 40180
rect 52612 40124 52622 40180
rect 56466 40124 56476 40180
rect 56532 40124 56868 40180
rect 56812 40068 56868 40124
rect 7522 40012 7532 40068
rect 7588 40012 8316 40068
rect 8372 40012 8382 40068
rect 11106 40012 11116 40068
rect 11172 40012 12124 40068
rect 12180 40012 12190 40068
rect 14578 40012 14588 40068
rect 14644 40012 21868 40068
rect 21924 40012 21934 40068
rect 36642 40012 36652 40068
rect 36708 40012 42812 40068
rect 42868 40012 42878 40068
rect 52434 40012 52444 40068
rect 52500 40012 53452 40068
rect 53508 40012 53518 40068
rect 53676 40012 53788 40068
rect 53844 40012 53854 40068
rect 56802 40012 56812 40068
rect 56868 40012 56878 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 53676 39956 53732 40012
rect 12562 39900 12572 39956
rect 12628 39900 13916 39956
rect 13972 39900 14140 39956
rect 14196 39900 14206 39956
rect 39330 39900 39340 39956
rect 39396 39900 53732 39956
rect 53862 39900 53900 39956
rect 53956 39900 53966 39956
rect 4022 39788 4060 39844
rect 4116 39788 4126 39844
rect 8418 39788 8428 39844
rect 8484 39788 9772 39844
rect 9828 39788 9838 39844
rect 37762 39788 37772 39844
rect 37828 39788 38332 39844
rect 38388 39788 38398 39844
rect 56690 39788 56700 39844
rect 56756 39788 57036 39844
rect 57092 39788 57102 39844
rect 200 39732 800 39760
rect 200 39676 1932 39732
rect 1988 39676 1998 39732
rect 7746 39676 7756 39732
rect 7812 39676 8652 39732
rect 8708 39676 8718 39732
rect 18946 39676 18956 39732
rect 19012 39676 20524 39732
rect 20580 39676 20590 39732
rect 20962 39676 20972 39732
rect 21028 39676 22092 39732
rect 22148 39676 22158 39732
rect 36530 39676 36540 39732
rect 36596 39676 38668 39732
rect 38724 39676 38734 39732
rect 38994 39676 39004 39732
rect 39060 39676 40460 39732
rect 40516 39676 41692 39732
rect 41748 39676 41758 39732
rect 43250 39676 43260 39732
rect 43316 39676 43372 39732
rect 43428 39676 43438 39732
rect 54198 39676 54236 39732
rect 54292 39676 54302 39732
rect 55906 39676 55916 39732
rect 55972 39676 56140 39732
rect 56196 39676 56206 39732
rect 200 39648 800 39676
rect 4386 39564 4396 39620
rect 4452 39564 5964 39620
rect 6020 39564 6030 39620
rect 19954 39564 19964 39620
rect 20020 39564 21084 39620
rect 21140 39564 21150 39620
rect 32946 39564 32956 39620
rect 33012 39564 40908 39620
rect 40964 39564 40974 39620
rect 42130 39564 42140 39620
rect 42196 39564 49084 39620
rect 49140 39564 50876 39620
rect 50932 39564 50942 39620
rect 51202 39564 51212 39620
rect 51268 39564 52108 39620
rect 52164 39564 52174 39620
rect 55234 39564 55244 39620
rect 55300 39564 57092 39620
rect 57670 39564 57708 39620
rect 57764 39564 57774 39620
rect 57036 39508 57092 39564
rect 8082 39452 8092 39508
rect 8148 39452 10668 39508
rect 10724 39452 17164 39508
rect 17220 39452 17230 39508
rect 19394 39452 19404 39508
rect 19460 39452 20188 39508
rect 20244 39452 20254 39508
rect 31378 39452 31388 39508
rect 31444 39452 31612 39508
rect 31668 39452 32844 39508
rect 32900 39452 32910 39508
rect 35634 39452 35644 39508
rect 35700 39452 36652 39508
rect 36708 39452 36718 39508
rect 37762 39452 37772 39508
rect 37828 39452 38556 39508
rect 38612 39452 40012 39508
rect 40068 39452 40078 39508
rect 42802 39452 42812 39508
rect 42868 39452 43260 39508
rect 43316 39452 43820 39508
rect 43876 39452 44044 39508
rect 44100 39452 44110 39508
rect 44370 39452 44380 39508
rect 44436 39452 54460 39508
rect 54516 39452 54526 39508
rect 54898 39452 54908 39508
rect 54964 39452 55804 39508
rect 55860 39452 55870 39508
rect 57026 39452 57036 39508
rect 57092 39452 57102 39508
rect 8530 39340 8540 39396
rect 8596 39340 11116 39396
rect 11172 39340 14028 39396
rect 14084 39340 14364 39396
rect 14420 39340 14430 39396
rect 16930 39340 16940 39396
rect 16996 39340 18060 39396
rect 18116 39340 19964 39396
rect 20020 39340 20030 39396
rect 21298 39340 21308 39396
rect 21364 39340 21532 39396
rect 21588 39340 22204 39396
rect 22260 39340 22652 39396
rect 22708 39340 23212 39396
rect 23268 39340 23278 39396
rect 24658 39340 24668 39396
rect 24724 39340 25228 39396
rect 25284 39340 25788 39396
rect 25844 39340 25854 39396
rect 27906 39340 27916 39396
rect 27972 39340 29708 39396
rect 29764 39340 29774 39396
rect 35074 39340 35084 39396
rect 35140 39340 37548 39396
rect 37604 39340 37884 39396
rect 37940 39340 37950 39396
rect 38434 39340 38444 39396
rect 38500 39340 39900 39396
rect 39956 39340 45276 39396
rect 45332 39340 45500 39396
rect 45556 39340 45566 39396
rect 46610 39340 46620 39396
rect 46676 39340 48524 39396
rect 48580 39340 48590 39396
rect 51426 39340 51436 39396
rect 51492 39340 53788 39396
rect 53844 39340 53854 39396
rect 56354 39340 56364 39396
rect 56420 39340 57596 39396
rect 57652 39340 57662 39396
rect 37884 39284 37940 39340
rect 13010 39228 13020 39284
rect 13076 39228 14476 39284
rect 14532 39228 16044 39284
rect 16100 39228 16110 39284
rect 29474 39228 29484 39284
rect 29540 39228 30044 39284
rect 30100 39228 30604 39284
rect 30660 39228 31164 39284
rect 31220 39228 31230 39284
rect 31938 39228 31948 39284
rect 32004 39228 35644 39284
rect 35700 39228 35710 39284
rect 37884 39228 39004 39284
rect 39060 39228 40572 39284
rect 40628 39228 40638 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 14886 39116 14924 39172
rect 14980 39116 14990 39172
rect 21074 39116 21084 39172
rect 21140 39116 21756 39172
rect 21812 39116 21822 39172
rect 30258 39116 30268 39172
rect 30324 39116 49532 39172
rect 49588 39116 49598 39172
rect 52322 39116 52332 39172
rect 52388 39116 53564 39172
rect 53620 39116 53676 39172
rect 53732 39116 53742 39172
rect 56130 39116 56140 39172
rect 56196 39116 57596 39172
rect 57652 39116 57662 39172
rect 3714 39004 3724 39060
rect 3780 39004 4732 39060
rect 4788 39004 4798 39060
rect 5394 39004 5404 39060
rect 5460 39004 5470 39060
rect 32274 39004 32284 39060
rect 32340 39004 33628 39060
rect 33684 39004 33694 39060
rect 38322 39004 38332 39060
rect 38388 39004 43148 39060
rect 43204 39004 44492 39060
rect 44548 39004 50988 39060
rect 51044 39004 51054 39060
rect 52098 39004 52108 39060
rect 52164 39004 53452 39060
rect 53508 39004 53518 39060
rect 54114 39004 54124 39060
rect 54180 39004 54460 39060
rect 54516 39004 54526 39060
rect 55010 39004 55020 39060
rect 55076 39004 57372 39060
rect 57428 39004 57438 39060
rect 5404 38836 5460 39004
rect 12114 38892 12124 38948
rect 12180 38892 12460 38948
rect 12516 38892 14924 38948
rect 14980 38892 17948 38948
rect 18004 38892 18014 38948
rect 20402 38892 20412 38948
rect 20468 38892 20860 38948
rect 20916 38892 21756 38948
rect 21812 38892 22988 38948
rect 23044 38892 28140 38948
rect 28196 38892 28206 38948
rect 41990 38892 42028 38948
rect 42084 38892 42094 38948
rect 45714 38892 45724 38948
rect 45780 38892 46508 38948
rect 46564 38892 46574 38948
rect 47282 38892 47292 38948
rect 47348 38892 51436 38948
rect 51492 38892 51502 38948
rect 51920 38892 51996 38948
rect 52052 38892 55244 38948
rect 55300 38892 55310 38948
rect 55682 38892 55692 38948
rect 55748 38892 57708 38948
rect 57764 38892 57774 38948
rect 3910 38780 3948 38836
rect 4004 38780 4014 38836
rect 4274 38780 4284 38836
rect 4340 38780 4620 38836
rect 4676 38780 6412 38836
rect 6468 38780 6478 38836
rect 13010 38780 13020 38836
rect 13076 38780 14868 38836
rect 15586 38780 15596 38836
rect 15652 38780 16044 38836
rect 16100 38780 16110 38836
rect 16594 38780 16604 38836
rect 16660 38780 17724 38836
rect 17780 38780 17790 38836
rect 24220 38780 24332 38836
rect 24388 38780 24398 38836
rect 30034 38780 30044 38836
rect 30100 38780 30380 38836
rect 30436 38780 30446 38836
rect 36754 38780 36764 38836
rect 36820 38780 37660 38836
rect 37716 38780 37726 38836
rect 41570 38780 41580 38836
rect 41636 38780 42476 38836
rect 42532 38780 42542 38836
rect 50530 38780 50540 38836
rect 50596 38780 53676 38836
rect 53732 38780 57484 38836
rect 57540 38780 57550 38836
rect 4386 38668 4396 38724
rect 4452 38668 5236 38724
rect 5180 38612 5236 38668
rect 5852 38612 5908 38780
rect 14812 38724 14868 38780
rect 6626 38668 6636 38724
rect 6692 38668 8092 38724
rect 8148 38668 8158 38724
rect 8978 38668 8988 38724
rect 9044 38668 9996 38724
rect 10052 38668 10332 38724
rect 10388 38668 10556 38724
rect 10612 38668 10622 38724
rect 11330 38668 11340 38724
rect 11396 38668 13916 38724
rect 13972 38668 13982 38724
rect 14812 38668 17164 38724
rect 17220 38668 17230 38724
rect 21196 38668 22204 38724
rect 22260 38668 22270 38724
rect 14812 38612 14868 38668
rect 21196 38612 21252 38668
rect 24220 38612 24276 38780
rect 26338 38668 26348 38724
rect 26404 38668 27020 38724
rect 27076 38668 28252 38724
rect 28308 38668 28318 38724
rect 33730 38668 33740 38724
rect 33796 38668 34188 38724
rect 34244 38668 37436 38724
rect 37492 38668 37502 38724
rect 38546 38668 38556 38724
rect 38612 38668 39228 38724
rect 39284 38668 39294 38724
rect 41906 38668 41916 38724
rect 41972 38668 42588 38724
rect 42644 38668 42654 38724
rect 52546 38668 52556 38724
rect 52612 38668 54908 38724
rect 54964 38668 54974 38724
rect 3938 38556 3948 38612
rect 4004 38556 4060 38612
rect 4116 38556 4126 38612
rect 4834 38556 4844 38612
rect 4900 38556 5180 38612
rect 5236 38556 5246 38612
rect 5842 38556 5852 38612
rect 5908 38556 5918 38612
rect 6738 38556 6748 38612
rect 6804 38556 7868 38612
rect 7924 38556 8652 38612
rect 8708 38556 8718 38612
rect 14802 38556 14812 38612
rect 14868 38556 14878 38612
rect 15138 38556 15148 38612
rect 15204 38556 15242 38612
rect 16930 38556 16940 38612
rect 16996 38556 19852 38612
rect 19908 38556 19918 38612
rect 21186 38556 21196 38612
rect 21252 38556 21262 38612
rect 23762 38556 23772 38612
rect 23828 38556 24276 38612
rect 24434 38556 24444 38612
rect 24500 38556 24780 38612
rect 24836 38556 25452 38612
rect 25508 38556 27804 38612
rect 27860 38556 27870 38612
rect 33954 38556 33964 38612
rect 34020 38556 55804 38612
rect 55860 38556 56252 38612
rect 56308 38556 56318 38612
rect 10210 38444 10220 38500
rect 10276 38444 11676 38500
rect 11732 38444 11742 38500
rect 15026 38444 15036 38500
rect 15092 38444 16156 38500
rect 16212 38444 16492 38500
rect 16548 38444 17388 38500
rect 17444 38444 19180 38500
rect 19236 38444 19740 38500
rect 19796 38444 19806 38500
rect 41682 38444 41692 38500
rect 41748 38444 42028 38500
rect 42084 38444 42094 38500
rect 45602 38444 45612 38500
rect 45668 38444 47068 38500
rect 47124 38444 47134 38500
rect 49522 38444 49532 38500
rect 49588 38444 57820 38500
rect 57876 38444 58604 38500
rect 58660 38444 58670 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 47068 38388 47124 38444
rect 14018 38332 14028 38388
rect 14084 38332 15148 38388
rect 15204 38332 15484 38388
rect 15540 38332 15550 38388
rect 17714 38332 17724 38388
rect 17780 38332 18732 38388
rect 18788 38332 19516 38388
rect 19572 38332 19582 38388
rect 20850 38332 20860 38388
rect 20916 38332 21980 38388
rect 22036 38332 22046 38388
rect 47068 38332 50204 38388
rect 50260 38332 50270 38388
rect 53330 38332 53340 38388
rect 53396 38332 53564 38388
rect 53620 38332 57932 38388
rect 57988 38332 57998 38388
rect 3938 38220 3948 38276
rect 4004 38220 4172 38276
rect 4228 38220 4732 38276
rect 4788 38220 10220 38276
rect 10276 38220 15148 38276
rect 16594 38220 16604 38276
rect 16660 38220 25340 38276
rect 25396 38220 25900 38276
rect 25956 38220 25966 38276
rect 36194 38220 36204 38276
rect 36260 38220 36764 38276
rect 36820 38220 36830 38276
rect 40786 38220 40796 38276
rect 40852 38220 49868 38276
rect 49924 38220 49934 38276
rect 52770 38220 52780 38276
rect 52836 38220 54012 38276
rect 54068 38220 54078 38276
rect 54646 38220 54684 38276
rect 54740 38220 54750 38276
rect 15092 38164 15148 38220
rect 4946 38108 4956 38164
rect 5012 38108 5628 38164
rect 5684 38108 5694 38164
rect 10546 38108 10556 38164
rect 10612 38108 11172 38164
rect 15092 38108 23212 38164
rect 23268 38108 23996 38164
rect 24052 38108 24062 38164
rect 33730 38108 33740 38164
rect 33796 38108 34076 38164
rect 34132 38108 34860 38164
rect 34916 38108 34926 38164
rect 43362 38108 43372 38164
rect 43428 38108 44716 38164
rect 44772 38108 44782 38164
rect 50372 38108 53452 38164
rect 53508 38108 58156 38164
rect 58212 38108 58222 38164
rect 11116 38052 11172 38108
rect 50372 38052 50428 38108
rect 3602 37996 3612 38052
rect 3668 37996 4620 38052
rect 4676 37996 4686 38052
rect 8866 37996 8876 38052
rect 8932 37996 9660 38052
rect 9716 37996 9726 38052
rect 10882 37996 10892 38052
rect 10948 37996 10958 38052
rect 11106 37996 11116 38052
rect 11172 37996 16604 38052
rect 16660 37996 16670 38052
rect 17602 37996 17612 38052
rect 17668 37996 18956 38052
rect 19012 37996 19022 38052
rect 24658 37996 24668 38052
rect 24724 37996 25900 38052
rect 25956 37996 26908 38052
rect 26964 37996 26974 38052
rect 28354 37996 28364 38052
rect 28420 37996 28812 38052
rect 28868 37996 29036 38052
rect 29092 37996 29102 38052
rect 30146 37996 30156 38052
rect 30212 37996 30716 38052
rect 30772 37996 30782 38052
rect 34262 37996 34300 38052
rect 34356 37996 34366 38052
rect 37762 37996 37772 38052
rect 37828 37996 38332 38052
rect 38388 37996 38398 38052
rect 44044 37996 50428 38052
rect 52322 37996 52332 38052
rect 52388 37996 52892 38052
rect 52948 37996 52958 38052
rect 54898 37996 54908 38052
rect 54964 37996 57596 38052
rect 57652 37996 57662 38052
rect 10892 37940 10948 37996
rect 44044 37940 44100 37996
rect 4274 37884 4284 37940
rect 4340 37884 4508 37940
rect 4564 37884 5964 37940
rect 6020 37884 6030 37940
rect 10892 37884 11228 37940
rect 11284 37884 15148 37940
rect 15250 37884 15260 37940
rect 15316 37884 16044 37940
rect 16100 37884 20860 37940
rect 20916 37884 20926 37940
rect 31042 37884 31052 37940
rect 31108 37884 31836 37940
rect 31892 37884 31902 37940
rect 34850 37884 34860 37940
rect 34916 37884 35644 37940
rect 35700 37884 35710 37940
rect 36530 37884 36540 37940
rect 36596 37884 37212 37940
rect 37268 37884 39004 37940
rect 39060 37884 39070 37940
rect 41430 37884 41468 37940
rect 41524 37884 44044 37940
rect 44100 37884 44110 37940
rect 44370 37884 44380 37940
rect 44436 37884 45500 37940
rect 45556 37884 45724 37940
rect 45780 37884 45790 37940
rect 45948 37884 48748 37940
rect 48804 37884 48814 37940
rect 55010 37884 55020 37940
rect 55076 37884 56924 37940
rect 56980 37884 56990 37940
rect 15092 37828 15148 37884
rect 38332 37828 38388 37884
rect 45948 37828 46004 37884
rect 4386 37772 4396 37828
rect 4452 37772 4956 37828
rect 5012 37772 6188 37828
rect 6244 37772 12348 37828
rect 12404 37772 12414 37828
rect 15092 37772 15932 37828
rect 15988 37772 15998 37828
rect 16146 37772 16156 37828
rect 16212 37772 16604 37828
rect 16660 37772 16670 37828
rect 20066 37772 20076 37828
rect 20132 37772 21532 37828
rect 21588 37772 22204 37828
rect 22260 37772 22270 37828
rect 29698 37772 29708 37828
rect 29764 37772 31500 37828
rect 31556 37772 31566 37828
rect 35074 37772 35084 37828
rect 35140 37772 36876 37828
rect 36932 37772 36942 37828
rect 38322 37772 38332 37828
rect 38388 37772 38398 37828
rect 44146 37772 44156 37828
rect 44212 37772 44492 37828
rect 44548 37772 46004 37828
rect 46834 37772 46844 37828
rect 46900 37772 48300 37828
rect 48356 37772 48366 37828
rect 50978 37772 50988 37828
rect 51044 37772 51212 37828
rect 51268 37772 51278 37828
rect 54786 37772 54796 37828
rect 54852 37772 56140 37828
rect 56196 37772 56206 37828
rect 4162 37660 4172 37716
rect 4228 37660 9100 37716
rect 9156 37660 9884 37716
rect 9940 37660 10892 37716
rect 10948 37660 10958 37716
rect 12226 37660 12236 37716
rect 12292 37660 12908 37716
rect 12964 37660 15260 37716
rect 15316 37660 15326 37716
rect 30818 37660 30828 37716
rect 30884 37660 31724 37716
rect 31780 37660 31790 37716
rect 35970 37660 35980 37716
rect 36036 37660 36204 37716
rect 36260 37660 36988 37716
rect 37044 37660 37054 37716
rect 40786 37660 40796 37716
rect 40852 37660 45612 37716
rect 45668 37660 45678 37716
rect 51090 37660 51100 37716
rect 51156 37660 51324 37716
rect 51380 37660 51884 37716
rect 51940 37660 52780 37716
rect 52836 37660 52846 37716
rect 53750 37660 53788 37716
rect 53844 37660 53854 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 11106 37548 11116 37604
rect 11172 37548 12460 37604
rect 12516 37548 12526 37604
rect 43138 37548 43148 37604
rect 43204 37548 44044 37604
rect 44100 37548 44110 37604
rect 50988 37548 58716 37604
rect 58772 37548 58782 37604
rect 50988 37492 51044 37548
rect 7858 37436 7868 37492
rect 7924 37436 7934 37492
rect 11554 37436 11564 37492
rect 11620 37436 11676 37492
rect 11732 37436 11742 37492
rect 12002 37436 12012 37492
rect 12068 37436 14364 37492
rect 14420 37436 14812 37492
rect 14868 37436 14878 37492
rect 15092 37436 16380 37492
rect 16436 37436 16446 37492
rect 18162 37436 18172 37492
rect 18228 37436 18620 37492
rect 18676 37436 18686 37492
rect 27346 37436 27356 37492
rect 27412 37436 29932 37492
rect 29988 37436 29998 37492
rect 32946 37436 32956 37492
rect 33012 37436 33516 37492
rect 33572 37436 33582 37492
rect 39554 37436 39564 37492
rect 39620 37436 40124 37492
rect 40180 37436 41468 37492
rect 41524 37436 41534 37492
rect 46050 37436 46060 37492
rect 46116 37436 51044 37492
rect 7868 37268 7924 37436
rect 15092 37380 15148 37436
rect 11442 37324 11452 37380
rect 11508 37324 13804 37380
rect 13860 37324 14588 37380
rect 14644 37324 15148 37380
rect 15586 37324 15596 37380
rect 15652 37324 18060 37380
rect 18116 37324 18126 37380
rect 18722 37324 18732 37380
rect 18788 37324 21532 37380
rect 21588 37324 22652 37380
rect 22708 37324 23436 37380
rect 23492 37324 23502 37380
rect 24770 37324 24780 37380
rect 24836 37324 25788 37380
rect 25844 37324 28028 37380
rect 28084 37324 28094 37380
rect 31154 37324 31164 37380
rect 31220 37324 32396 37380
rect 32452 37324 32620 37380
rect 32676 37324 32686 37380
rect 40898 37324 40908 37380
rect 40964 37324 41692 37380
rect 41748 37324 42028 37380
rect 42084 37324 43036 37380
rect 43092 37324 46396 37380
rect 46452 37324 46462 37380
rect 47506 37324 47516 37380
rect 47572 37324 52164 37380
rect 52322 37324 52332 37380
rect 52388 37324 53228 37380
rect 53284 37324 53564 37380
rect 53620 37324 53630 37380
rect 52108 37268 52164 37324
rect 7186 37212 7196 37268
rect 7252 37212 7924 37268
rect 13122 37212 13132 37268
rect 13188 37212 14924 37268
rect 14980 37212 15148 37268
rect 15204 37212 16044 37268
rect 16100 37212 16110 37268
rect 19058 37212 19068 37268
rect 19124 37212 19964 37268
rect 20020 37212 20030 37268
rect 29698 37212 29708 37268
rect 29764 37212 30828 37268
rect 30884 37212 30894 37268
rect 31826 37212 31836 37268
rect 31892 37212 32732 37268
rect 32788 37212 33628 37268
rect 33684 37212 33694 37268
rect 34402 37212 34412 37268
rect 34468 37212 39900 37268
rect 39956 37212 40460 37268
rect 40516 37212 40526 37268
rect 41234 37212 41244 37268
rect 41300 37212 41916 37268
rect 41972 37212 42476 37268
rect 42532 37212 42812 37268
rect 42868 37212 42878 37268
rect 43922 37212 43932 37268
rect 43988 37212 45276 37268
rect 45332 37212 46284 37268
rect 46340 37212 46350 37268
rect 48402 37212 48412 37268
rect 48468 37212 50540 37268
rect 50596 37212 50606 37268
rect 52098 37212 52108 37268
rect 52164 37212 53004 37268
rect 53060 37212 53070 37268
rect 55794 37212 55804 37268
rect 55860 37212 58268 37268
rect 58324 37212 58334 37268
rect 55804 37156 55860 37212
rect 4610 37100 4620 37156
rect 4676 37100 5180 37156
rect 5236 37100 5628 37156
rect 5684 37100 6300 37156
rect 6356 37100 14252 37156
rect 14308 37100 14318 37156
rect 17714 37100 17724 37156
rect 17780 37100 18620 37156
rect 18676 37100 18686 37156
rect 29474 37100 29484 37156
rect 29540 37100 31052 37156
rect 31108 37100 31118 37156
rect 32050 37100 32060 37156
rect 32116 37100 32126 37156
rect 39666 37100 39676 37156
rect 39732 37100 40796 37156
rect 40852 37100 40862 37156
rect 42018 37100 42028 37156
rect 42084 37100 43260 37156
rect 43316 37100 43326 37156
rect 44146 37100 44156 37156
rect 44212 37100 46620 37156
rect 46676 37100 46686 37156
rect 51174 37100 51212 37156
rect 51268 37100 51278 37156
rect 54460 37100 55860 37156
rect 56578 37100 56588 37156
rect 56644 37100 57484 37156
rect 57540 37100 57550 37156
rect 12898 36988 12908 37044
rect 12964 36988 13356 37044
rect 13412 36988 13422 37044
rect 14466 36988 14476 37044
rect 14532 36988 18172 37044
rect 18228 36988 18238 37044
rect 20850 36988 20860 37044
rect 20916 36988 21756 37044
rect 21812 36988 21822 37044
rect 6626 36876 6636 36932
rect 6692 36876 6972 36932
rect 7028 36876 7308 36932
rect 7364 36876 7374 36932
rect 8642 36876 8652 36932
rect 8708 36876 9548 36932
rect 9604 36876 9614 36932
rect 13234 36876 13244 36932
rect 13300 36876 15260 36932
rect 15316 36876 15326 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 8418 36764 8428 36820
rect 8484 36764 9324 36820
rect 9380 36764 10332 36820
rect 10388 36764 10398 36820
rect 16930 36764 16940 36820
rect 16996 36764 17164 36820
rect 17220 36764 18172 36820
rect 18228 36764 18238 36820
rect 13906 36652 13916 36708
rect 13972 36652 15148 36708
rect 15204 36652 15280 36708
rect 20738 36652 20748 36708
rect 20804 36652 20814 36708
rect 20748 36596 20804 36652
rect 14578 36540 14588 36596
rect 14644 36540 15372 36596
rect 15428 36540 15596 36596
rect 15652 36540 15820 36596
rect 15876 36540 15886 36596
rect 20514 36540 20524 36596
rect 20580 36540 20804 36596
rect 32060 36484 32116 37100
rect 54460 37044 54516 37100
rect 59200 37044 59800 37072
rect 35746 36988 35756 37044
rect 35812 36988 36204 37044
rect 36260 36988 36764 37044
rect 36820 36988 38780 37044
rect 38836 36988 38846 37044
rect 43362 36988 43372 37044
rect 43428 36988 44268 37044
rect 44324 36988 44604 37044
rect 44660 36988 44670 37044
rect 46162 36988 46172 37044
rect 46228 36988 47180 37044
rect 47236 36988 47246 37044
rect 48514 36988 48524 37044
rect 48580 36988 54516 37044
rect 55682 36988 55692 37044
rect 55748 36988 59800 37044
rect 59200 36960 59800 36988
rect 38994 36876 39004 36932
rect 39060 36876 48188 36932
rect 48244 36876 48254 36932
rect 52994 36876 53004 36932
rect 53060 36876 53788 36932
rect 53844 36876 53854 36932
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 36978 36764 36988 36820
rect 37044 36764 37436 36820
rect 37492 36764 54124 36820
rect 54180 36764 54190 36820
rect 38658 36652 38668 36708
rect 38724 36652 41860 36708
rect 45042 36652 45052 36708
rect 45108 36652 45500 36708
rect 45556 36652 45566 36708
rect 47282 36652 47292 36708
rect 47348 36652 48524 36708
rect 48580 36652 48590 36708
rect 49634 36652 49644 36708
rect 49700 36652 49710 36708
rect 52434 36652 52444 36708
rect 52500 36652 52510 36708
rect 41804 36596 41860 36652
rect 49644 36596 49700 36652
rect 52444 36596 52500 36652
rect 33170 36540 33180 36596
rect 33236 36540 40572 36596
rect 40628 36540 41580 36596
rect 41636 36540 41646 36596
rect 41804 36540 49700 36596
rect 52210 36540 52220 36596
rect 52276 36540 52500 36596
rect 52658 36540 52668 36596
rect 52724 36540 53956 36596
rect 53900 36484 53956 36540
rect 9762 36428 9772 36484
rect 9828 36428 11900 36484
rect 11956 36428 13468 36484
rect 13524 36428 14812 36484
rect 14868 36428 14878 36484
rect 15138 36428 15148 36484
rect 15204 36428 16044 36484
rect 16100 36428 16110 36484
rect 17042 36428 17052 36484
rect 17108 36428 17948 36484
rect 18004 36428 18014 36484
rect 32060 36428 32172 36484
rect 32228 36428 32238 36484
rect 32722 36428 32732 36484
rect 32788 36428 33628 36484
rect 33684 36428 38556 36484
rect 38612 36428 38622 36484
rect 38770 36428 38780 36484
rect 38836 36428 39676 36484
rect 39732 36428 39742 36484
rect 44482 36428 44492 36484
rect 44548 36428 45276 36484
rect 45332 36428 45836 36484
rect 45892 36428 45902 36484
rect 52098 36428 52108 36484
rect 52164 36428 53340 36484
rect 53396 36428 53406 36484
rect 53890 36428 53900 36484
rect 53956 36428 55468 36484
rect 55524 36428 55534 36484
rect 33180 36372 33236 36428
rect 11526 36316 11564 36372
rect 11620 36316 11630 36372
rect 14690 36316 14700 36372
rect 14756 36316 20412 36372
rect 20468 36316 21644 36372
rect 21700 36316 21710 36372
rect 24546 36316 24556 36372
rect 24612 36316 26068 36372
rect 33170 36316 33180 36372
rect 33236 36316 33246 36372
rect 37986 36316 37996 36372
rect 38052 36316 38220 36372
rect 38276 36316 40572 36372
rect 40628 36316 44156 36372
rect 44212 36316 44222 36372
rect 44594 36316 44604 36372
rect 44660 36316 47292 36372
rect 47348 36316 48188 36372
rect 48244 36316 49756 36372
rect 49812 36316 49822 36372
rect 52434 36316 52444 36372
rect 52500 36316 53676 36372
rect 53732 36316 53742 36372
rect 56802 36316 56812 36372
rect 56868 36316 58156 36372
rect 58212 36316 58222 36372
rect 26012 36260 26068 36316
rect 6290 36204 6300 36260
rect 6356 36204 6972 36260
rect 7028 36204 7252 36260
rect 9426 36204 9436 36260
rect 9492 36204 10220 36260
rect 10276 36204 10668 36260
rect 10724 36204 10734 36260
rect 12898 36204 12908 36260
rect 12964 36204 14028 36260
rect 14084 36204 14588 36260
rect 14644 36204 14654 36260
rect 16482 36204 16492 36260
rect 16548 36204 17276 36260
rect 17332 36204 17724 36260
rect 17780 36204 20244 36260
rect 24098 36204 24108 36260
rect 24164 36204 25676 36260
rect 25732 36204 25742 36260
rect 26002 36204 26012 36260
rect 26068 36204 26684 36260
rect 26740 36204 26750 36260
rect 30706 36204 30716 36260
rect 30772 36204 31276 36260
rect 31332 36204 31342 36260
rect 38658 36204 38668 36260
rect 38724 36204 39116 36260
rect 39172 36204 40348 36260
rect 40404 36204 40414 36260
rect 42466 36204 42476 36260
rect 42532 36204 43260 36260
rect 43316 36204 43326 36260
rect 45154 36204 45164 36260
rect 45220 36204 45948 36260
rect 46004 36204 46014 36260
rect 53330 36204 53340 36260
rect 53396 36204 55132 36260
rect 55188 36204 55198 36260
rect 7196 36036 7252 36204
rect 20188 36148 20244 36204
rect 20188 36092 24892 36148
rect 24948 36092 24958 36148
rect 57250 36092 57260 36148
rect 57316 36092 57820 36148
rect 57876 36092 57886 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 7186 35980 7196 36036
rect 7252 35980 9548 36036
rect 9604 35980 9996 36036
rect 10052 35980 10062 36036
rect 30482 35980 30492 36036
rect 30548 35980 31948 36036
rect 32004 35980 32396 36036
rect 32452 35980 32462 36036
rect 34150 35980 34188 36036
rect 34244 35980 34254 36036
rect 34636 35980 37268 36036
rect 38546 35980 38556 36036
rect 38612 35980 44380 36036
rect 44436 35980 44446 36036
rect 46396 35980 47180 36036
rect 47236 35980 47246 36036
rect 3332 35868 26796 35924
rect 26852 35868 26862 35924
rect 31826 35868 31836 35924
rect 31892 35868 33068 35924
rect 33124 35868 33134 35924
rect 3332 35812 3388 35868
rect 2930 35756 2940 35812
rect 2996 35756 3388 35812
rect 9650 35756 9660 35812
rect 9716 35756 11228 35812
rect 11284 35756 11788 35812
rect 11844 35756 11854 35812
rect 24882 35756 24892 35812
rect 24948 35756 27356 35812
rect 27412 35756 28364 35812
rect 28420 35756 28430 35812
rect 34636 35700 34692 35980
rect 37212 35924 37268 35980
rect 46396 35924 46452 35980
rect 36306 35868 36316 35924
rect 36372 35868 36988 35924
rect 37044 35868 37054 35924
rect 37212 35868 46452 35924
rect 46722 35868 46732 35924
rect 46788 35868 51660 35924
rect 51716 35868 52668 35924
rect 52724 35868 52734 35924
rect 53778 35868 53788 35924
rect 53844 35868 54012 35924
rect 54068 35868 54078 35924
rect 36418 35756 36428 35812
rect 36484 35756 37436 35812
rect 37492 35756 37772 35812
rect 37828 35756 38220 35812
rect 38276 35756 38286 35812
rect 43362 35756 43372 35812
rect 43428 35756 43708 35812
rect 43764 35756 44604 35812
rect 44660 35756 45164 35812
rect 45220 35756 45230 35812
rect 50530 35756 50540 35812
rect 50596 35756 51548 35812
rect 51604 35756 51614 35812
rect 51874 35756 51884 35812
rect 51940 35756 56588 35812
rect 56644 35756 56654 35812
rect 7298 35644 7308 35700
rect 7364 35644 8652 35700
rect 8708 35644 8718 35700
rect 16706 35644 16716 35700
rect 16772 35644 27468 35700
rect 27524 35644 27534 35700
rect 30492 35644 34692 35700
rect 35298 35644 35308 35700
rect 35364 35644 35374 35700
rect 37090 35644 37100 35700
rect 37156 35644 38108 35700
rect 38164 35644 38444 35700
rect 38500 35644 38510 35700
rect 38882 35644 38892 35700
rect 38948 35644 39564 35700
rect 39620 35644 39630 35700
rect 49746 35644 49756 35700
rect 49812 35644 50204 35700
rect 50260 35644 50428 35700
rect 50484 35644 50494 35700
rect 30492 35588 30548 35644
rect 35308 35588 35364 35644
rect 51884 35588 51940 35756
rect 56242 35644 56252 35700
rect 56308 35644 57036 35700
rect 57092 35644 57708 35700
rect 57764 35644 57774 35700
rect 7746 35532 7756 35588
rect 7812 35532 9324 35588
rect 9380 35532 9390 35588
rect 13234 35532 13244 35588
rect 13300 35532 14252 35588
rect 14308 35532 14318 35588
rect 18274 35532 18284 35588
rect 18340 35532 18956 35588
rect 19012 35532 19292 35588
rect 19348 35532 19358 35588
rect 30482 35532 30492 35588
rect 30548 35532 30558 35588
rect 31490 35532 31500 35588
rect 31556 35532 32788 35588
rect 34738 35532 34748 35588
rect 34804 35532 37436 35588
rect 37492 35532 37502 35588
rect 38658 35532 38668 35588
rect 38724 35532 39788 35588
rect 39844 35532 41020 35588
rect 41076 35532 41468 35588
rect 41524 35532 41534 35588
rect 43698 35532 43708 35588
rect 43764 35532 44492 35588
rect 44548 35532 44558 35588
rect 47170 35532 47180 35588
rect 47236 35532 49532 35588
rect 49588 35532 49598 35588
rect 49970 35532 49980 35588
rect 50036 35532 51940 35588
rect 52210 35532 52220 35588
rect 52276 35532 53228 35588
rect 53284 35532 55580 35588
rect 55636 35532 56028 35588
rect 56084 35532 56094 35588
rect 32732 35476 32788 35532
rect 41468 35476 41524 35532
rect 2258 35420 2268 35476
rect 2324 35420 9884 35476
rect 9940 35420 9950 35476
rect 18386 35420 18396 35476
rect 18452 35420 18844 35476
rect 18900 35420 18910 35476
rect 29698 35420 29708 35476
rect 29764 35420 31612 35476
rect 31668 35420 31678 35476
rect 32722 35420 32732 35476
rect 32788 35420 34972 35476
rect 35028 35420 35038 35476
rect 41468 35420 46060 35476
rect 46116 35420 53452 35476
rect 53508 35420 53518 35476
rect 55458 35420 55468 35476
rect 55524 35420 56252 35476
rect 56308 35420 57484 35476
rect 57540 35420 57550 35476
rect 10210 35308 10220 35364
rect 10276 35308 11004 35364
rect 11060 35308 11340 35364
rect 11396 35308 20300 35364
rect 20356 35308 20860 35364
rect 20916 35308 20926 35364
rect 30034 35308 30044 35364
rect 30100 35308 30604 35364
rect 30660 35308 30670 35364
rect 41458 35308 41468 35364
rect 41524 35308 42924 35364
rect 42980 35308 42990 35364
rect 51986 35308 51996 35364
rect 52052 35308 52108 35364
rect 52164 35308 52174 35364
rect 54786 35308 54796 35364
rect 54852 35308 56028 35364
rect 56084 35308 56094 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 39890 35196 39900 35252
rect 39956 35196 41916 35252
rect 41972 35196 41982 35252
rect 46834 35196 46844 35252
rect 46900 35196 48412 35252
rect 48468 35196 52556 35252
rect 52612 35196 52622 35252
rect 4834 35084 4844 35140
rect 4900 35084 8876 35140
rect 8932 35084 9996 35140
rect 10052 35084 10062 35140
rect 20402 35084 20412 35140
rect 20468 35084 21868 35140
rect 21924 35084 21934 35140
rect 50866 35084 50876 35140
rect 50932 35084 51996 35140
rect 52052 35084 52062 35140
rect 4946 34972 4956 35028
rect 5012 34972 6188 35028
rect 6244 34972 6254 35028
rect 7186 34972 7196 35028
rect 7252 34972 9100 35028
rect 9156 34972 24108 35028
rect 24164 34972 24332 35028
rect 24388 34972 24398 35028
rect 55122 34972 55132 35028
rect 55188 34972 55692 35028
rect 55748 34972 55758 35028
rect 56914 34972 56924 35028
rect 56980 34972 58044 35028
rect 58100 34972 58110 35028
rect 2258 34860 2268 34916
rect 2324 34860 2828 34916
rect 2884 34860 3500 34916
rect 3556 34860 3566 34916
rect 6262 34860 6300 34916
rect 6356 34860 6366 34916
rect 10658 34860 10668 34916
rect 10724 34860 11340 34916
rect 11396 34860 11406 34916
rect 11554 34860 11564 34916
rect 11620 34860 12012 34916
rect 12068 34860 12078 34916
rect 12786 34860 12796 34916
rect 12852 34860 13692 34916
rect 13748 34860 13758 34916
rect 14802 34860 14812 34916
rect 14868 34860 15148 34916
rect 15204 34860 16492 34916
rect 16548 34860 16558 34916
rect 21074 34860 21084 34916
rect 21140 34860 23212 34916
rect 23268 34860 23772 34916
rect 23828 34860 25564 34916
rect 25620 34860 27804 34916
rect 27860 34860 27870 34916
rect 39218 34860 39228 34916
rect 39284 34860 40236 34916
rect 40292 34860 40302 34916
rect 48738 34860 48748 34916
rect 48804 34860 51996 34916
rect 52052 34860 52062 34916
rect 53778 34860 53788 34916
rect 53844 34860 54460 34916
rect 54516 34860 55356 34916
rect 55412 34860 55422 34916
rect 55580 34860 55804 34916
rect 55860 34860 55870 34916
rect 13234 34748 13244 34804
rect 13300 34748 13804 34804
rect 13860 34748 13870 34804
rect 15026 34748 15036 34804
rect 15092 34748 15932 34804
rect 15988 34748 15998 34804
rect 20514 34748 20524 34804
rect 20580 34748 21980 34804
rect 22036 34748 22428 34804
rect 22484 34748 23660 34804
rect 23716 34748 24780 34804
rect 24836 34748 24846 34804
rect 37538 34748 37548 34804
rect 37604 34748 39004 34804
rect 39060 34748 39070 34804
rect 15036 34692 15092 34748
rect 39228 34692 39284 34860
rect 55580 34804 55636 34860
rect 41234 34748 41244 34804
rect 41300 34748 41580 34804
rect 41636 34748 41646 34804
rect 44370 34748 44380 34804
rect 44436 34748 44492 34804
rect 44548 34748 44558 34804
rect 48626 34748 48636 34804
rect 48692 34748 48972 34804
rect 49028 34748 49038 34804
rect 50372 34748 51324 34804
rect 51380 34748 53340 34804
rect 53396 34748 53564 34804
rect 53620 34748 53630 34804
rect 55570 34748 55580 34804
rect 55636 34748 55646 34804
rect 56578 34748 56588 34804
rect 56644 34748 58268 34804
rect 58324 34748 58334 34804
rect 50372 34692 50428 34748
rect 4050 34636 4060 34692
rect 4116 34636 4732 34692
rect 4788 34636 4956 34692
rect 5012 34636 5022 34692
rect 13570 34636 13580 34692
rect 13636 34636 15092 34692
rect 19282 34636 19292 34692
rect 19348 34636 21420 34692
rect 21476 34636 21644 34692
rect 21700 34636 21710 34692
rect 31826 34636 31836 34692
rect 31892 34636 32396 34692
rect 32452 34636 32462 34692
rect 33730 34636 33740 34692
rect 33796 34636 34412 34692
rect 34468 34636 34478 34692
rect 36978 34636 36988 34692
rect 37044 34636 39284 34692
rect 42242 34636 42252 34692
rect 42308 34636 43932 34692
rect 43988 34636 45612 34692
rect 45668 34636 45678 34692
rect 47842 34636 47852 34692
rect 47908 34636 50428 34692
rect 52882 34636 52892 34692
rect 52948 34636 54684 34692
rect 54740 34636 54750 34692
rect 55682 34636 55692 34692
rect 55748 34636 58044 34692
rect 58100 34636 58940 34692
rect 58996 34636 59006 34692
rect 33740 34580 33796 34636
rect 30930 34524 30940 34580
rect 30996 34524 31724 34580
rect 31780 34524 33796 34580
rect 36082 34524 36092 34580
rect 36148 34524 37548 34580
rect 37604 34524 37614 34580
rect 38994 34524 39004 34580
rect 39060 34524 39340 34580
rect 39396 34524 40348 34580
rect 40404 34524 40414 34580
rect 45154 34524 45164 34580
rect 45220 34524 46844 34580
rect 46900 34524 46910 34580
rect 53890 34524 53900 34580
rect 53956 34524 56252 34580
rect 56308 34524 56318 34580
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 9762 34412 9772 34468
rect 9828 34412 9884 34468
rect 9940 34412 12012 34468
rect 12068 34412 12078 34468
rect 45042 34412 45052 34468
rect 45108 34412 47292 34468
rect 47348 34412 47358 34468
rect 51986 34412 51996 34468
rect 52052 34412 53900 34468
rect 53956 34412 53966 34468
rect 200 34356 800 34384
rect 200 34300 1932 34356
rect 1988 34300 1998 34356
rect 6626 34300 6636 34356
rect 6692 34300 6972 34356
rect 7028 34300 8428 34356
rect 8484 34300 8494 34356
rect 8978 34300 8988 34356
rect 9044 34300 11004 34356
rect 11060 34300 11070 34356
rect 16594 34300 16604 34356
rect 16660 34300 18844 34356
rect 18900 34300 19180 34356
rect 19236 34300 21420 34356
rect 21476 34300 21486 34356
rect 31154 34300 31164 34356
rect 31220 34300 32284 34356
rect 32340 34300 32350 34356
rect 43026 34300 43036 34356
rect 43092 34300 43484 34356
rect 43540 34300 46396 34356
rect 46452 34300 46462 34356
rect 47618 34300 47628 34356
rect 47684 34300 48636 34356
rect 48692 34300 52332 34356
rect 52388 34300 52398 34356
rect 52556 34300 55132 34356
rect 55188 34300 55198 34356
rect 200 34272 800 34300
rect 52556 34244 52612 34300
rect 7186 34188 7196 34244
rect 7252 34188 7980 34244
rect 8036 34188 8046 34244
rect 9090 34188 9100 34244
rect 9156 34188 9660 34244
rect 9716 34188 9726 34244
rect 11218 34188 11228 34244
rect 11284 34188 11900 34244
rect 11956 34188 11966 34244
rect 18162 34188 18172 34244
rect 18228 34188 26348 34244
rect 26404 34188 27020 34244
rect 27076 34188 27086 34244
rect 40002 34188 40012 34244
rect 40068 34188 41244 34244
rect 41300 34188 41310 34244
rect 43922 34188 43932 34244
rect 43988 34188 49308 34244
rect 49364 34188 49644 34244
rect 49700 34188 49710 34244
rect 50204 34188 50652 34244
rect 50708 34188 50988 34244
rect 51044 34188 51884 34244
rect 51940 34188 52612 34244
rect 52770 34188 52780 34244
rect 52836 34188 55580 34244
rect 55636 34188 55646 34244
rect 50204 34132 50260 34188
rect 7410 34076 7420 34132
rect 7476 34076 16884 34132
rect 21746 34076 21756 34132
rect 21812 34076 26124 34132
rect 26180 34076 26190 34132
rect 30146 34076 30156 34132
rect 30212 34076 30828 34132
rect 30884 34076 30894 34132
rect 43586 34076 43596 34132
rect 43652 34076 46284 34132
rect 46340 34076 46350 34132
rect 46834 34076 46844 34132
rect 46900 34076 50204 34132
rect 50260 34076 50270 34132
rect 53106 34076 53116 34132
rect 53172 34076 54684 34132
rect 54740 34076 56140 34132
rect 56196 34076 56206 34132
rect 56550 34076 56588 34132
rect 56644 34076 56654 34132
rect 16828 34020 16884 34076
rect 6066 33964 6076 34020
rect 6132 33964 7756 34020
rect 7812 33964 7822 34020
rect 11218 33964 11228 34020
rect 11284 33964 13244 34020
rect 13300 33964 13310 34020
rect 14802 33964 14812 34020
rect 14868 33964 15036 34020
rect 15092 33964 15102 34020
rect 15810 33964 15820 34020
rect 15876 33964 16604 34020
rect 16660 33964 16670 34020
rect 16828 33964 24556 34020
rect 24612 33964 24622 34020
rect 43250 33964 43260 34020
rect 43316 33964 44940 34020
rect 44996 33964 45052 34020
rect 45108 33964 48524 34020
rect 48580 33964 48590 34020
rect 49410 33964 49420 34020
rect 49476 33964 58044 34020
rect 58100 33964 58110 34020
rect 7298 33852 7308 33908
rect 7364 33852 8540 33908
rect 8596 33852 8606 33908
rect 12898 33852 12908 33908
rect 12964 33852 13356 33908
rect 13412 33852 14252 33908
rect 14308 33852 15932 33908
rect 15988 33852 15998 33908
rect 36306 33852 36316 33908
rect 36372 33852 36764 33908
rect 36820 33852 39900 33908
rect 39956 33852 40460 33908
rect 40516 33852 40526 33908
rect 44258 33852 44268 33908
rect 44324 33852 47740 33908
rect 47796 33852 53508 33908
rect 54898 33852 54908 33908
rect 54964 33852 55244 33908
rect 55300 33852 55310 33908
rect 8978 33740 8988 33796
rect 9044 33740 11788 33796
rect 11844 33740 11854 33796
rect 12226 33740 12236 33796
rect 12292 33740 17612 33796
rect 17668 33740 18060 33796
rect 18116 33740 19292 33796
rect 19348 33740 19740 33796
rect 19796 33740 19806 33796
rect 47618 33740 47628 33796
rect 47684 33740 47964 33796
rect 48020 33740 48030 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 53452 33684 53508 33852
rect 53666 33740 53676 33796
rect 53732 33740 55468 33796
rect 55524 33740 55534 33796
rect 5842 33628 5852 33684
rect 5908 33628 11788 33684
rect 11844 33628 11854 33684
rect 12002 33628 12012 33684
rect 12068 33628 15932 33684
rect 15988 33628 15998 33684
rect 35532 33628 35644 33684
rect 35700 33628 35710 33684
rect 35858 33628 35868 33684
rect 35924 33628 36316 33684
rect 36372 33628 37772 33684
rect 37828 33628 38108 33684
rect 38164 33628 38174 33684
rect 40226 33628 40236 33684
rect 40292 33628 42028 33684
rect 42084 33628 42094 33684
rect 43810 33628 43820 33684
rect 43876 33628 44156 33684
rect 44212 33628 45164 33684
rect 45220 33628 45230 33684
rect 45490 33628 45500 33684
rect 45556 33628 48188 33684
rect 48244 33628 48254 33684
rect 50988 33628 51716 33684
rect 53452 33628 55804 33684
rect 55860 33628 55870 33684
rect 35532 33572 35588 33628
rect 50988 33572 51044 33628
rect 51660 33572 51716 33628
rect 6290 33516 6300 33572
rect 6356 33516 7868 33572
rect 7924 33516 9100 33572
rect 9156 33516 9166 33572
rect 14914 33516 14924 33572
rect 14980 33516 15820 33572
rect 15876 33516 15886 33572
rect 24322 33516 24332 33572
rect 24388 33516 25116 33572
rect 25172 33516 26908 33572
rect 26964 33516 26974 33572
rect 29474 33516 29484 33572
rect 29540 33516 29932 33572
rect 29988 33516 30604 33572
rect 30660 33516 30670 33572
rect 33730 33516 33740 33572
rect 33796 33516 34972 33572
rect 35028 33516 35038 33572
rect 35298 33516 35308 33572
rect 35364 33516 35588 33572
rect 38434 33516 38444 33572
rect 38500 33516 40572 33572
rect 40628 33516 51044 33572
rect 51202 33516 51212 33572
rect 51268 33516 51436 33572
rect 51492 33516 51502 33572
rect 51660 33516 52724 33572
rect 52882 33516 52892 33572
rect 52948 33516 53564 33572
rect 53620 33516 56476 33572
rect 56532 33516 56542 33572
rect 52668 33460 52724 33516
rect 4498 33404 4508 33460
rect 4564 33404 5068 33460
rect 5124 33404 7308 33460
rect 7364 33404 7374 33460
rect 8306 33404 8316 33460
rect 8372 33404 10108 33460
rect 10164 33404 10174 33460
rect 16034 33404 16044 33460
rect 16100 33404 22540 33460
rect 22596 33404 22606 33460
rect 27010 33404 27020 33460
rect 27076 33404 27356 33460
rect 27412 33404 28812 33460
rect 28868 33404 29708 33460
rect 29764 33404 30716 33460
rect 30772 33404 30782 33460
rect 45378 33404 45388 33460
rect 45444 33404 45948 33460
rect 46004 33404 46620 33460
rect 46676 33404 46686 33460
rect 49858 33404 49868 33460
rect 49924 33404 51548 33460
rect 51604 33404 51614 33460
rect 52668 33404 54348 33460
rect 54404 33404 57260 33460
rect 57316 33404 57326 33460
rect 6738 33292 6748 33348
rect 6804 33292 9212 33348
rect 9268 33292 9278 33348
rect 26562 33292 26572 33348
rect 26628 33292 27580 33348
rect 27636 33292 27646 33348
rect 28018 33292 28028 33348
rect 28084 33292 28476 33348
rect 28532 33292 28542 33348
rect 32498 33292 32508 33348
rect 32564 33292 33292 33348
rect 33348 33292 33358 33348
rect 33506 33292 33516 33348
rect 33572 33292 34636 33348
rect 34692 33292 34702 33348
rect 40002 33292 40012 33348
rect 40068 33292 41580 33348
rect 41636 33292 41646 33348
rect 42018 33292 42028 33348
rect 42084 33292 44156 33348
rect 44212 33292 47292 33348
rect 47348 33292 47358 33348
rect 50950 33292 50988 33348
rect 51044 33292 51054 33348
rect 54002 33292 54012 33348
rect 54068 33292 57932 33348
rect 57988 33292 57998 33348
rect 11890 33180 11900 33236
rect 11956 33180 12460 33236
rect 12516 33180 13580 33236
rect 13636 33180 13646 33236
rect 22082 33180 22092 33236
rect 22148 33180 24444 33236
rect 24500 33180 24510 33236
rect 39778 33180 39788 33236
rect 39844 33180 41020 33236
rect 41076 33180 41086 33236
rect 41234 33180 41244 33236
rect 41300 33180 41916 33236
rect 41972 33180 43764 33236
rect 48066 33180 48076 33236
rect 48132 33180 51212 33236
rect 51268 33180 51278 33236
rect 52668 33180 53564 33236
rect 53620 33180 54572 33236
rect 54628 33180 54638 33236
rect 55906 33180 55916 33236
rect 55972 33180 56924 33236
rect 56980 33180 58716 33236
rect 58772 33180 58782 33236
rect 43708 33124 43764 33180
rect 52668 33124 52724 33180
rect 7186 33068 7196 33124
rect 7252 33068 7980 33124
rect 8036 33068 8046 33124
rect 8194 33068 8204 33124
rect 8260 33068 8428 33124
rect 8484 33068 8494 33124
rect 12338 33068 12348 33124
rect 12404 33068 12908 33124
rect 12964 33068 13692 33124
rect 13748 33068 13758 33124
rect 16594 33068 16604 33124
rect 16660 33068 17724 33124
rect 17780 33068 17790 33124
rect 18610 33068 18620 33124
rect 18676 33068 19180 33124
rect 19236 33068 22988 33124
rect 23044 33068 23054 33124
rect 30258 33068 30268 33124
rect 30324 33068 30828 33124
rect 30884 33068 30894 33124
rect 32386 33068 32396 33124
rect 32452 33068 33628 33124
rect 33684 33068 33852 33124
rect 33908 33068 33918 33124
rect 36866 33068 36876 33124
rect 36932 33068 39228 33124
rect 39284 33068 39294 33124
rect 40786 33068 40796 33124
rect 40852 33068 43260 33124
rect 43316 33068 43326 33124
rect 43698 33068 43708 33124
rect 43764 33068 49868 33124
rect 49924 33068 49934 33124
rect 50372 33068 50988 33124
rect 51044 33068 52332 33124
rect 52388 33068 52398 33124
rect 52658 33068 52668 33124
rect 52724 33068 52734 33124
rect 53106 33068 53116 33124
rect 53172 33068 53340 33124
rect 53396 33068 53406 33124
rect 50372 33012 50428 33068
rect 5730 32956 5740 33012
rect 5796 32956 9660 33012
rect 9716 32956 9726 33012
rect 22866 32956 22876 33012
rect 22932 32956 23884 33012
rect 23940 32956 26012 33012
rect 26068 32956 26572 33012
rect 26628 32956 26638 33012
rect 37538 32956 37548 33012
rect 37604 32956 38556 33012
rect 38612 32956 47068 33012
rect 47124 32956 47852 33012
rect 47908 32956 48524 33012
rect 48580 32956 48590 33012
rect 49970 32956 49980 33012
rect 50036 32956 50428 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 53116 32900 53172 33068
rect 39666 32844 39676 32900
rect 39732 32844 40908 32900
rect 40964 32844 41692 32900
rect 41748 32844 41758 32900
rect 42578 32844 42588 32900
rect 42644 32844 42924 32900
rect 42980 32844 42990 32900
rect 44482 32844 44492 32900
rect 44548 32844 46508 32900
rect 46564 32844 46574 32900
rect 47142 32844 47180 32900
rect 47236 32844 47246 32900
rect 52322 32844 52332 32900
rect 52388 32844 53172 32900
rect 42588 32788 42644 32844
rect 11666 32732 11676 32788
rect 11732 32732 29372 32788
rect 29428 32732 29438 32788
rect 39442 32732 39452 32788
rect 39508 32732 42644 32788
rect 47012 32732 50428 32788
rect 50754 32732 50764 32788
rect 50820 32732 51660 32788
rect 51716 32732 51726 32788
rect 53414 32732 53452 32788
rect 53508 32732 53518 32788
rect 47012 32676 47068 32732
rect 6514 32620 6524 32676
rect 6580 32620 8764 32676
rect 8820 32620 9772 32676
rect 9828 32620 9838 32676
rect 14018 32620 14028 32676
rect 14084 32620 15036 32676
rect 15092 32620 16492 32676
rect 16548 32620 16558 32676
rect 20626 32620 20636 32676
rect 20692 32620 20860 32676
rect 20916 32620 21532 32676
rect 21588 32620 21756 32676
rect 21812 32620 21822 32676
rect 24210 32620 24220 32676
rect 24276 32620 27356 32676
rect 27412 32620 27422 32676
rect 37426 32620 37436 32676
rect 37492 32620 38444 32676
rect 38500 32620 38510 32676
rect 39452 32620 47068 32676
rect 50372 32620 50428 32732
rect 50484 32620 51772 32676
rect 51828 32620 57932 32676
rect 57988 32620 57998 32676
rect 1586 32508 1596 32564
rect 1652 32508 3836 32564
rect 3892 32508 10108 32564
rect 10164 32508 10174 32564
rect 12450 32508 12460 32564
rect 12516 32508 13468 32564
rect 13524 32508 13534 32564
rect 13682 32508 13692 32564
rect 13748 32508 16156 32564
rect 16212 32508 16222 32564
rect 16370 32508 16380 32564
rect 16436 32508 17724 32564
rect 17780 32508 17790 32564
rect 18050 32508 18060 32564
rect 18116 32508 20524 32564
rect 20580 32508 23772 32564
rect 23828 32508 23838 32564
rect 26114 32508 26124 32564
rect 26180 32508 26796 32564
rect 26852 32508 26862 32564
rect 34066 32508 34076 32564
rect 34132 32508 35532 32564
rect 35588 32508 36092 32564
rect 36148 32508 36158 32564
rect 36418 32508 36428 32564
rect 36484 32508 38892 32564
rect 38948 32508 38958 32564
rect 16380 32452 16436 32508
rect 39452 32452 39508 32620
rect 39666 32508 39676 32564
rect 39732 32508 42252 32564
rect 42308 32508 43036 32564
rect 43092 32508 43102 32564
rect 44258 32508 44268 32564
rect 44324 32508 45612 32564
rect 45668 32508 45678 32564
rect 47282 32508 47292 32564
rect 47348 32508 47516 32564
rect 47572 32508 47582 32564
rect 50166 32508 50204 32564
rect 50260 32508 56588 32564
rect 56644 32508 56654 32564
rect 57138 32508 57148 32564
rect 57204 32508 57820 32564
rect 57876 32508 58716 32564
rect 58772 32508 58782 32564
rect 47516 32452 47572 32508
rect 2482 32396 2492 32452
rect 2548 32396 4284 32452
rect 4340 32396 4350 32452
rect 5170 32396 5180 32452
rect 5236 32396 5404 32452
rect 5460 32396 5852 32452
rect 5908 32396 5918 32452
rect 8642 32396 8652 32452
rect 8708 32396 10892 32452
rect 10948 32396 10958 32452
rect 12674 32396 12684 32452
rect 12740 32396 14140 32452
rect 14196 32396 14476 32452
rect 14532 32396 14542 32452
rect 14914 32396 14924 32452
rect 14980 32396 16436 32452
rect 29922 32396 29932 32452
rect 29988 32396 30492 32452
rect 30548 32396 30558 32452
rect 32834 32396 32844 32452
rect 32900 32396 33740 32452
rect 33796 32396 34188 32452
rect 34244 32396 34254 32452
rect 38098 32396 38108 32452
rect 38164 32396 39508 32452
rect 40450 32396 40460 32452
rect 40516 32396 41468 32452
rect 41524 32396 44492 32452
rect 44548 32396 44828 32452
rect 44884 32396 44894 32452
rect 47516 32396 52332 32452
rect 52388 32396 52398 32452
rect 53666 32396 53676 32452
rect 53732 32396 56812 32452
rect 56868 32396 56878 32452
rect 5618 32284 5628 32340
rect 5684 32284 6300 32340
rect 6356 32284 6366 32340
rect 11732 32284 17500 32340
rect 17556 32284 17566 32340
rect 21298 32284 21308 32340
rect 21364 32284 22652 32340
rect 22708 32284 23100 32340
rect 23156 32284 23772 32340
rect 23828 32284 24780 32340
rect 24836 32284 24846 32340
rect 43810 32284 43820 32340
rect 43876 32284 44604 32340
rect 44660 32284 44670 32340
rect 47954 32284 47964 32340
rect 48020 32284 49532 32340
rect 49588 32284 49598 32340
rect 49970 32284 49980 32340
rect 50036 32284 50764 32340
rect 50820 32284 50830 32340
rect 11732 32228 11788 32284
rect 5618 32172 5628 32228
rect 5684 32172 11788 32228
rect 16146 32172 16156 32228
rect 16212 32172 22036 32228
rect 22194 32172 22204 32228
rect 22260 32172 22270 32228
rect 42578 32172 42588 32228
rect 42644 32172 43036 32228
rect 43092 32172 51044 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 5058 32060 5068 32116
rect 5124 32060 5740 32116
rect 5796 32060 6188 32116
rect 6244 32060 6254 32116
rect 8418 32060 8428 32116
rect 8484 32060 17276 32116
rect 17332 32060 17342 32116
rect 21980 32004 22036 32172
rect 22204 32116 22260 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 22204 32060 23100 32116
rect 23156 32060 23166 32116
rect 36194 32060 36204 32116
rect 36260 32060 36988 32116
rect 37044 32060 37054 32116
rect 41570 32060 41580 32116
rect 41636 32060 43372 32116
rect 43428 32060 43438 32116
rect 45042 32060 45052 32116
rect 45108 32060 45118 32116
rect 46274 32060 46284 32116
rect 46340 32060 48636 32116
rect 48692 32060 48702 32116
rect 49606 32060 49644 32116
rect 49700 32060 49710 32116
rect 45052 32004 45108 32060
rect 50988 32004 51044 32172
rect 53974 32060 54012 32116
rect 54068 32060 54078 32116
rect 54562 32060 54572 32116
rect 54628 32060 57148 32116
rect 57204 32060 57214 32116
rect 4834 31948 4844 32004
rect 4900 31948 5292 32004
rect 5348 31948 6076 32004
rect 6132 31948 6748 32004
rect 6804 31948 6814 32004
rect 10210 31948 10220 32004
rect 10276 31948 10724 32004
rect 14130 31948 14140 32004
rect 14196 31948 16156 32004
rect 16212 31948 16222 32004
rect 16380 31948 16492 32004
rect 16548 31948 17276 32004
rect 17332 31948 18060 32004
rect 18116 31948 19628 32004
rect 19684 31948 19694 32004
rect 21980 31948 25340 32004
rect 25396 31948 26012 32004
rect 26068 31948 26684 32004
rect 26740 31948 27692 32004
rect 27748 31948 27758 32004
rect 32946 31948 32956 32004
rect 33012 31948 34524 32004
rect 34580 31948 34590 32004
rect 35858 31948 35868 32004
rect 35924 31948 36428 32004
rect 36484 31948 36494 32004
rect 41906 31948 41916 32004
rect 41972 31948 42700 32004
rect 42756 31948 42766 32004
rect 42924 31948 43708 32004
rect 43764 31948 44492 32004
rect 44548 31948 44558 32004
rect 45052 31948 45276 32004
rect 45332 31948 45342 32004
rect 45714 31948 45724 32004
rect 45780 31948 46508 32004
rect 46564 31948 49980 32004
rect 50036 31948 50046 32004
rect 50978 31948 50988 32004
rect 51044 31948 52108 32004
rect 52164 31948 52174 32004
rect 52434 31948 52444 32004
rect 52500 31948 53340 32004
rect 53396 31948 53406 32004
rect 53666 31948 53676 32004
rect 53732 31948 56140 32004
rect 56196 31948 56206 32004
rect 10668 31892 10724 31948
rect 8530 31836 8540 31892
rect 8596 31836 10332 31892
rect 10388 31836 10398 31892
rect 10658 31836 10668 31892
rect 10724 31836 10734 31892
rect 12338 31836 12348 31892
rect 12404 31836 12796 31892
rect 12852 31836 13356 31892
rect 13412 31836 13916 31892
rect 13972 31836 13982 31892
rect 14700 31780 14756 31948
rect 16380 31892 16436 31948
rect 42924 31892 42980 31948
rect 16034 31836 16044 31892
rect 16100 31836 16436 31892
rect 19394 31836 19404 31892
rect 19460 31836 20188 31892
rect 20244 31836 20254 31892
rect 21746 31836 21756 31892
rect 21812 31836 22540 31892
rect 22596 31836 23660 31892
rect 23716 31836 24444 31892
rect 24500 31836 24510 31892
rect 31378 31836 31388 31892
rect 31444 31836 31948 31892
rect 32004 31836 32014 31892
rect 36530 31836 36540 31892
rect 36596 31836 36988 31892
rect 37044 31836 37054 31892
rect 38546 31836 38556 31892
rect 38612 31836 42980 31892
rect 43138 31836 43148 31892
rect 43204 31836 44044 31892
rect 44100 31836 45052 31892
rect 45108 31836 45118 31892
rect 45490 31836 45500 31892
rect 45556 31836 46284 31892
rect 46340 31836 46956 31892
rect 47012 31836 47022 31892
rect 47394 31836 47404 31892
rect 47460 31836 47964 31892
rect 48020 31836 48412 31892
rect 48468 31836 48478 31892
rect 48626 31836 48636 31892
rect 48692 31836 49756 31892
rect 49812 31836 51268 31892
rect 51426 31836 51436 31892
rect 51492 31836 55244 31892
rect 55300 31836 57372 31892
rect 57428 31836 57438 31892
rect 51212 31780 51268 31836
rect 3378 31724 3388 31780
rect 3444 31724 10388 31780
rect 14690 31724 14700 31780
rect 14756 31724 14766 31780
rect 21858 31724 21868 31780
rect 21924 31724 22428 31780
rect 22484 31724 22494 31780
rect 23202 31724 23212 31780
rect 23268 31724 23996 31780
rect 24052 31724 24668 31780
rect 24724 31724 24734 31780
rect 33730 31724 33740 31780
rect 33796 31724 34860 31780
rect 34916 31724 34926 31780
rect 35746 31724 35756 31780
rect 35812 31724 37436 31780
rect 37492 31724 37502 31780
rect 38434 31724 38444 31780
rect 38500 31724 40124 31780
rect 40180 31724 41468 31780
rect 41524 31724 41534 31780
rect 43026 31724 43036 31780
rect 43092 31724 43484 31780
rect 43540 31724 44156 31780
rect 44212 31724 44222 31780
rect 46834 31724 46844 31780
rect 46900 31724 47740 31780
rect 47796 31724 47806 31780
rect 48850 31724 48860 31780
rect 48916 31724 49308 31780
rect 49364 31724 49374 31780
rect 51202 31724 51212 31780
rect 51268 31724 51278 31780
rect 51660 31724 52220 31780
rect 52276 31724 52668 31780
rect 52724 31724 52734 31780
rect 53890 31724 53900 31780
rect 53956 31724 56476 31780
rect 56532 31724 56542 31780
rect 56802 31724 56812 31780
rect 56868 31724 57484 31780
rect 57540 31724 57550 31780
rect 10332 31668 10388 31724
rect 51660 31668 51716 31724
rect 59200 31668 59800 31696
rect 4162 31612 4172 31668
rect 4228 31612 6524 31668
rect 6580 31612 6590 31668
rect 6850 31612 6860 31668
rect 6916 31612 7532 31668
rect 7588 31612 8428 31668
rect 8484 31612 8494 31668
rect 10322 31612 10332 31668
rect 10388 31612 10398 31668
rect 19394 31612 19404 31668
rect 19460 31612 20076 31668
rect 20132 31612 20142 31668
rect 42690 31612 42700 31668
rect 42756 31612 43820 31668
rect 43876 31612 43886 31668
rect 44044 31612 49980 31668
rect 50036 31612 50046 31668
rect 50194 31612 50204 31668
rect 50260 31612 51716 31668
rect 53666 31612 53676 31668
rect 53732 31612 53770 31668
rect 56018 31612 56028 31668
rect 56084 31612 59800 31668
rect 44044 31556 44100 31612
rect 59200 31584 59800 31612
rect 2342 31500 2380 31556
rect 2436 31500 2446 31556
rect 2818 31500 2828 31556
rect 2884 31500 3500 31556
rect 3556 31500 4844 31556
rect 4900 31500 4910 31556
rect 5730 31500 5740 31556
rect 5796 31500 6412 31556
rect 6468 31500 6478 31556
rect 10434 31500 10444 31556
rect 10500 31500 10780 31556
rect 10836 31500 10846 31556
rect 16594 31500 16604 31556
rect 16660 31500 17948 31556
rect 18004 31500 18508 31556
rect 18564 31500 18574 31556
rect 34962 31500 34972 31556
rect 35028 31500 35420 31556
rect 35476 31500 35486 31556
rect 36306 31500 36316 31556
rect 36372 31500 37660 31556
rect 37716 31500 37726 31556
rect 38658 31500 38668 31556
rect 38724 31500 38780 31556
rect 38836 31500 38846 31556
rect 40898 31500 40908 31556
rect 40964 31500 43260 31556
rect 43316 31500 44100 31556
rect 44258 31500 44268 31556
rect 44324 31500 45948 31556
rect 46004 31500 46014 31556
rect 46722 31500 46732 31556
rect 46788 31500 47068 31556
rect 47124 31500 47134 31556
rect 47506 31500 47516 31556
rect 47572 31500 48524 31556
rect 48580 31500 48590 31556
rect 49746 31500 49756 31556
rect 49812 31500 51044 31556
rect 51202 31500 51212 31556
rect 51268 31500 53452 31556
rect 53508 31500 57820 31556
rect 57876 31500 57886 31556
rect 50988 31444 51044 31500
rect 2258 31388 2268 31444
rect 2324 31388 5068 31444
rect 5124 31388 5134 31444
rect 7746 31388 7756 31444
rect 7812 31388 8316 31444
rect 8372 31388 8382 31444
rect 10098 31388 10108 31444
rect 10164 31388 15036 31444
rect 15092 31388 15102 31444
rect 22978 31388 22988 31444
rect 23044 31388 27020 31444
rect 27076 31388 27086 31444
rect 35522 31388 35532 31444
rect 35588 31388 35756 31444
rect 35812 31388 35822 31444
rect 36530 31388 36540 31444
rect 36596 31388 37996 31444
rect 38052 31388 38062 31444
rect 43922 31388 43932 31444
rect 43988 31388 48300 31444
rect 48356 31388 48366 31444
rect 50988 31388 53452 31444
rect 53508 31388 53676 31444
rect 53732 31388 53742 31444
rect 54898 31388 54908 31444
rect 54964 31388 58492 31444
rect 58548 31388 58558 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 35756 31332 35812 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 3938 31276 3948 31332
rect 4004 31276 15148 31332
rect 21634 31276 21644 31332
rect 21700 31276 22204 31332
rect 22260 31276 23660 31332
rect 23716 31276 23884 31332
rect 23940 31276 24220 31332
rect 24276 31276 24780 31332
rect 24836 31276 24846 31332
rect 31154 31276 31164 31332
rect 31220 31276 31230 31332
rect 35756 31276 38556 31332
rect 38612 31276 38622 31332
rect 42018 31276 42028 31332
rect 42084 31276 45892 31332
rect 46274 31276 46284 31332
rect 46340 31276 50316 31332
rect 50372 31276 50382 31332
rect 51426 31276 51436 31332
rect 51492 31276 51996 31332
rect 52052 31276 53004 31332
rect 53060 31276 53070 31332
rect 15092 31220 15148 31276
rect 3826 31164 3836 31220
rect 3892 31164 4620 31220
rect 4676 31164 4686 31220
rect 4834 31164 4844 31220
rect 4900 31164 10892 31220
rect 10948 31164 10958 31220
rect 15092 31164 29484 31220
rect 29540 31164 29550 31220
rect 4620 31108 4676 31164
rect 4620 31052 5852 31108
rect 5908 31052 5918 31108
rect 7522 31052 7532 31108
rect 7588 31052 8316 31108
rect 8372 31052 8382 31108
rect 11106 31052 11116 31108
rect 11172 31052 12684 31108
rect 12740 31052 12750 31108
rect 19394 31052 19404 31108
rect 19460 31052 19964 31108
rect 20020 31052 20030 31108
rect 24882 31052 24892 31108
rect 24948 31052 26236 31108
rect 26292 31052 26302 31108
rect 8082 30940 8092 30996
rect 8148 30940 8652 30996
rect 8708 30940 8718 30996
rect 12226 30940 12236 30996
rect 12292 30940 13020 30996
rect 13076 30940 13692 30996
rect 13748 30940 13758 30996
rect 19506 30940 19516 30996
rect 19572 30940 19852 30996
rect 19908 30940 19918 30996
rect 20066 30940 20076 30996
rect 20132 30940 22540 30996
rect 22596 30940 22606 30996
rect 24546 30940 24556 30996
rect 24612 30940 25564 30996
rect 25620 30940 25630 30996
rect 31164 30884 31220 31276
rect 45836 31220 45892 31276
rect 31490 31164 31500 31220
rect 31556 31164 31948 31220
rect 32004 31164 32732 31220
rect 32788 31164 33180 31220
rect 33236 31164 33246 31220
rect 40898 31164 40908 31220
rect 40964 31164 44268 31220
rect 44324 31164 44334 31220
rect 44930 31164 44940 31220
rect 44996 31164 45388 31220
rect 45444 31164 45454 31220
rect 45826 31164 45836 31220
rect 45892 31164 50428 31220
rect 50484 31164 51548 31220
rect 51604 31164 51614 31220
rect 53078 31164 53116 31220
rect 53172 31164 53182 31220
rect 55318 31164 55356 31220
rect 55412 31164 55422 31220
rect 31378 31052 31388 31108
rect 31444 31052 33628 31108
rect 33684 31052 33694 31108
rect 39778 31052 39788 31108
rect 39844 31052 40796 31108
rect 40852 31052 43148 31108
rect 43204 31052 43214 31108
rect 44818 31052 44828 31108
rect 44884 31052 47516 31108
rect 47572 31052 47582 31108
rect 48290 31052 48300 31108
rect 48356 31052 50540 31108
rect 50596 31052 52332 31108
rect 52388 31052 52398 31108
rect 34290 30940 34300 30996
rect 34356 30940 35308 30996
rect 35364 30940 35644 30996
rect 35700 30940 35710 30996
rect 43026 30940 43036 30996
rect 43092 30940 43820 30996
rect 43876 30940 43886 30996
rect 47618 30940 47628 30996
rect 47684 30940 50876 30996
rect 50932 30940 55916 30996
rect 55972 30940 57596 30996
rect 57652 30940 57662 30996
rect 6962 30828 6972 30884
rect 7028 30828 7532 30884
rect 7588 30828 7598 30884
rect 8418 30828 8428 30884
rect 8484 30828 9884 30884
rect 9940 30828 9950 30884
rect 10546 30828 10556 30884
rect 10612 30828 10668 30884
rect 10724 30828 10734 30884
rect 11778 30828 11788 30884
rect 11844 30828 16044 30884
rect 16100 30828 26796 30884
rect 26852 30828 26862 30884
rect 31164 30828 31276 30884
rect 31332 30828 31342 30884
rect 34178 30828 34188 30884
rect 34244 30828 34748 30884
rect 34804 30828 34972 30884
rect 35028 30828 35038 30884
rect 42578 30828 42588 30884
rect 42644 30828 43148 30884
rect 43204 30828 46284 30884
rect 46340 30828 46956 30884
rect 47012 30828 47022 30884
rect 47954 30828 47964 30884
rect 48020 30828 54124 30884
rect 54180 30828 54190 30884
rect 7532 30772 7588 30828
rect 3826 30716 3836 30772
rect 3892 30716 4172 30772
rect 4228 30716 4900 30772
rect 7532 30716 8092 30772
rect 8148 30716 9660 30772
rect 9716 30716 10220 30772
rect 10276 30716 10286 30772
rect 11442 30716 11452 30772
rect 11508 30716 11788 30772
rect 11844 30716 11854 30772
rect 19618 30716 19628 30772
rect 19684 30716 22540 30772
rect 22596 30716 22606 30772
rect 35410 30716 35420 30772
rect 35476 30716 38668 30772
rect 38724 30716 38734 30772
rect 42130 30716 42140 30772
rect 42196 30716 48188 30772
rect 48244 30716 48254 30772
rect 50866 30716 50876 30772
rect 50932 30716 51660 30772
rect 51716 30716 51726 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 4844 30548 4900 30716
rect 7522 30604 7532 30660
rect 7588 30604 8540 30660
rect 8596 30604 8876 30660
rect 8932 30604 8942 30660
rect 10882 30604 10892 30660
rect 10948 30604 12012 30660
rect 12068 30604 12078 30660
rect 38658 30604 38668 30660
rect 38724 30604 39900 30660
rect 39956 30604 41468 30660
rect 41524 30604 41534 30660
rect 42914 30604 42924 30660
rect 42980 30604 43932 30660
rect 43988 30604 43998 30660
rect 44594 30604 44604 30660
rect 44660 30604 45164 30660
rect 45220 30604 45230 30660
rect 49970 30604 49980 30660
rect 50036 30604 56588 30660
rect 56644 30604 56700 30660
rect 56756 30604 56766 30660
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 4844 30492 11284 30548
rect 12114 30492 12124 30548
rect 12180 30492 15372 30548
rect 15428 30492 15438 30548
rect 22082 30492 22092 30548
rect 22148 30492 22764 30548
rect 22820 30492 22830 30548
rect 38406 30492 38444 30548
rect 38500 30492 38510 30548
rect 38612 30492 43596 30548
rect 43652 30492 43662 30548
rect 49970 30492 49980 30548
rect 50036 30492 54236 30548
rect 54292 30492 54302 30548
rect 5282 30380 5292 30436
rect 5348 30380 5740 30436
rect 5796 30380 5806 30436
rect 6178 30380 6188 30436
rect 6244 30380 6636 30436
rect 6692 30380 7756 30436
rect 7812 30380 7822 30436
rect 11228 30324 11284 30492
rect 38612 30436 38668 30492
rect 15092 30380 29932 30436
rect 29988 30380 29998 30436
rect 30146 30380 30156 30436
rect 30212 30380 31500 30436
rect 31556 30380 31566 30436
rect 32834 30380 32844 30436
rect 32900 30380 33516 30436
rect 33572 30380 38668 30436
rect 39676 30380 47292 30436
rect 47348 30380 47358 30436
rect 47964 30380 50204 30436
rect 50260 30380 50270 30436
rect 50362 30380 50372 30436
rect 50428 30380 52164 30436
rect 52546 30380 52556 30436
rect 52612 30380 54796 30436
rect 54852 30380 54862 30436
rect 15092 30324 15148 30380
rect 39676 30324 39732 30380
rect 5954 30268 5964 30324
rect 6020 30268 6748 30324
rect 6804 30268 6814 30324
rect 7410 30268 7420 30324
rect 7476 30268 8316 30324
rect 8372 30268 9100 30324
rect 9156 30268 10780 30324
rect 10836 30268 10846 30324
rect 11228 30268 15148 30324
rect 17714 30268 17724 30324
rect 17780 30268 18396 30324
rect 18452 30268 18462 30324
rect 18610 30268 18620 30324
rect 18676 30268 18956 30324
rect 19012 30268 19022 30324
rect 19730 30268 19740 30324
rect 19796 30268 19964 30324
rect 20020 30268 20030 30324
rect 20290 30268 20300 30324
rect 20356 30268 20860 30324
rect 20916 30268 21980 30324
rect 22036 30268 23212 30324
rect 23268 30268 23278 30324
rect 34738 30268 34748 30324
rect 34804 30268 38892 30324
rect 38948 30268 39732 30324
rect 42242 30268 42252 30324
rect 42308 30268 42476 30324
rect 42532 30268 42542 30324
rect 45714 30268 45724 30324
rect 45780 30268 47068 30324
rect 47124 30268 47134 30324
rect 47964 30212 48020 30380
rect 52108 30324 52164 30380
rect 48178 30268 48188 30324
rect 48244 30268 48804 30324
rect 49522 30268 49532 30324
rect 49588 30268 50428 30324
rect 50484 30268 50494 30324
rect 52108 30268 53788 30324
rect 53844 30268 53854 30324
rect 57474 30268 57484 30324
rect 57540 30268 57550 30324
rect 24434 30156 24444 30212
rect 24500 30156 24780 30212
rect 24836 30156 24846 30212
rect 28130 30156 28140 30212
rect 28196 30156 28700 30212
rect 28756 30156 29932 30212
rect 29988 30156 30716 30212
rect 30772 30156 30782 30212
rect 30930 30156 30940 30212
rect 30996 30156 32284 30212
rect 32340 30156 35756 30212
rect 35812 30156 35822 30212
rect 40422 30156 40460 30212
rect 40516 30156 40526 30212
rect 40786 30156 40796 30212
rect 40852 30156 46172 30212
rect 46228 30156 46238 30212
rect 46732 30156 48020 30212
rect 48748 30212 48804 30268
rect 57484 30212 57540 30268
rect 48748 30156 51996 30212
rect 52052 30156 54684 30212
rect 54740 30156 54750 30212
rect 55132 30156 57540 30212
rect 46732 30100 46788 30156
rect 3714 30044 3724 30100
rect 3780 30044 6412 30100
rect 6468 30044 6478 30100
rect 6626 30044 6636 30100
rect 6692 30044 7084 30100
rect 7140 30044 7150 30100
rect 11106 30044 11116 30100
rect 11172 30044 11676 30100
rect 11732 30044 11742 30100
rect 14130 30044 14140 30100
rect 14196 30044 15148 30100
rect 15204 30044 15214 30100
rect 18694 30044 18732 30100
rect 18788 30044 18798 30100
rect 29586 30044 29596 30100
rect 29652 30044 30828 30100
rect 30884 30044 30894 30100
rect 33842 30044 33852 30100
rect 33908 30044 34188 30100
rect 34244 30044 34254 30100
rect 34402 30044 34412 30100
rect 34468 30044 35084 30100
rect 35140 30044 35150 30100
rect 35634 30044 35644 30100
rect 35700 30044 36652 30100
rect 36708 30044 41244 30100
rect 41300 30044 41310 30100
rect 42130 30044 42140 30100
rect 42196 30044 43596 30100
rect 43652 30044 43820 30100
rect 43876 30044 43886 30100
rect 44044 30044 45500 30100
rect 45556 30044 46788 30100
rect 51090 30044 51100 30100
rect 51156 30044 52444 30100
rect 52500 30044 52510 30100
rect 44044 29988 44100 30044
rect 55132 29988 55188 30156
rect 55542 30044 55580 30100
rect 55636 30044 55646 30100
rect 56578 30044 56588 30100
rect 56644 30044 56700 30100
rect 56756 30044 56766 30100
rect 3826 29932 3836 29988
rect 3892 29932 5068 29988
rect 5124 29932 5134 29988
rect 5590 29932 5628 29988
rect 5684 29932 5694 29988
rect 5954 29932 5964 29988
rect 6020 29932 6300 29988
rect 6356 29932 6366 29988
rect 7634 29932 7644 29988
rect 7700 29932 8652 29988
rect 8708 29932 8718 29988
rect 9538 29932 9548 29988
rect 9604 29932 10892 29988
rect 10948 29932 10958 29988
rect 12674 29932 12684 29988
rect 12740 29932 17276 29988
rect 17332 29932 18060 29988
rect 18116 29932 18396 29988
rect 18452 29932 18462 29988
rect 28466 29932 28476 29988
rect 28532 29932 30716 29988
rect 30772 29932 30782 29988
rect 31826 29932 31836 29988
rect 31892 29932 33180 29988
rect 33236 29932 33246 29988
rect 34514 29932 34524 29988
rect 34580 29932 38108 29988
rect 38164 29932 38174 29988
rect 38434 29932 38444 29988
rect 38500 29932 39116 29988
rect 39172 29932 40796 29988
rect 40852 29932 40862 29988
rect 42578 29932 42588 29988
rect 42644 29932 44100 29988
rect 45378 29932 45388 29988
rect 45444 29932 46396 29988
rect 46452 29932 46462 29988
rect 50372 29932 53340 29988
rect 53396 29932 53406 29988
rect 54674 29932 54684 29988
rect 54740 29932 55132 29988
rect 55188 29932 55198 29988
rect 4946 29820 4956 29876
rect 5012 29820 5516 29876
rect 5572 29820 10444 29876
rect 10500 29820 13468 29876
rect 13524 29820 13534 29876
rect 14354 29820 14364 29876
rect 14420 29820 14476 29876
rect 14532 29820 15260 29876
rect 15316 29820 15326 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 31836 29764 31892 29932
rect 50372 29876 50428 29932
rect 33730 29820 33740 29876
rect 33796 29820 35644 29876
rect 35700 29820 35710 29876
rect 36530 29820 36540 29876
rect 36596 29820 40012 29876
rect 40068 29820 40078 29876
rect 40562 29820 40572 29876
rect 40628 29820 43036 29876
rect 43092 29820 43102 29876
rect 44034 29820 44044 29876
rect 44100 29820 44156 29876
rect 44212 29820 44940 29876
rect 44996 29820 45006 29876
rect 47506 29820 47516 29876
rect 47572 29820 50428 29876
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 8614 29708 8652 29764
rect 8708 29708 9884 29764
rect 9940 29708 9950 29764
rect 11890 29708 11900 29764
rect 11956 29708 12908 29764
rect 12964 29708 12974 29764
rect 28802 29708 28812 29764
rect 28868 29708 30716 29764
rect 30772 29708 31892 29764
rect 37202 29708 37212 29764
rect 37268 29708 39340 29764
rect 39396 29708 39406 29764
rect 40674 29708 40684 29764
rect 40740 29708 43484 29764
rect 43540 29708 43550 29764
rect 44044 29708 50204 29764
rect 50260 29708 50270 29764
rect 52322 29708 52332 29764
rect 52388 29708 55580 29764
rect 55636 29708 55646 29764
rect 2146 29596 2156 29652
rect 2212 29596 3388 29652
rect 3444 29596 4620 29652
rect 4676 29596 4686 29652
rect 8418 29596 8428 29652
rect 8484 29596 9548 29652
rect 9604 29596 9614 29652
rect 11218 29596 11228 29652
rect 11284 29596 11564 29652
rect 11620 29596 11630 29652
rect 20962 29596 20972 29652
rect 21028 29596 21868 29652
rect 21924 29596 21934 29652
rect 23538 29596 23548 29652
rect 23604 29596 25900 29652
rect 25956 29596 26236 29652
rect 26292 29596 26302 29652
rect 29474 29596 29484 29652
rect 29540 29596 30492 29652
rect 30548 29596 30558 29652
rect 36754 29596 36764 29652
rect 36820 29596 37772 29652
rect 37828 29596 38332 29652
rect 38388 29596 39004 29652
rect 39060 29596 39070 29652
rect 41682 29596 41692 29652
rect 41748 29596 43820 29652
rect 43876 29596 43886 29652
rect 44044 29540 44100 29708
rect 47170 29596 47180 29652
rect 47236 29596 47964 29652
rect 48020 29596 48748 29652
rect 48804 29596 48814 29652
rect 4834 29484 4844 29540
rect 4900 29484 5628 29540
rect 5684 29484 5694 29540
rect 7074 29484 7084 29540
rect 7140 29484 7532 29540
rect 7588 29484 7598 29540
rect 10994 29484 11004 29540
rect 11060 29484 11070 29540
rect 15810 29484 15820 29540
rect 15876 29484 16492 29540
rect 16548 29484 16828 29540
rect 16884 29484 27580 29540
rect 27636 29484 27916 29540
rect 27972 29484 27982 29540
rect 37874 29484 37884 29540
rect 37940 29484 38220 29540
rect 38276 29484 41580 29540
rect 41636 29484 41646 29540
rect 42354 29484 42364 29540
rect 42420 29484 42812 29540
rect 42868 29484 44100 29540
rect 48066 29484 48076 29540
rect 48132 29484 49980 29540
rect 50036 29484 50046 29540
rect 50866 29484 50876 29540
rect 50932 29484 51772 29540
rect 51828 29484 51838 29540
rect 56476 29484 58828 29540
rect 58884 29484 59500 29540
rect 59556 29484 59566 29540
rect 11004 29428 11060 29484
rect 56476 29428 56532 29484
rect 6178 29372 6188 29428
rect 6244 29372 6972 29428
rect 7028 29372 7308 29428
rect 7364 29372 7374 29428
rect 10434 29372 10444 29428
rect 10500 29372 11564 29428
rect 11620 29372 11630 29428
rect 12226 29372 12236 29428
rect 12292 29372 14252 29428
rect 14308 29372 14588 29428
rect 14644 29372 16268 29428
rect 16324 29372 16334 29428
rect 17266 29372 17276 29428
rect 17332 29372 17836 29428
rect 17892 29372 18620 29428
rect 18676 29372 19628 29428
rect 19684 29372 20412 29428
rect 20468 29372 20478 29428
rect 20738 29372 20748 29428
rect 20804 29372 21196 29428
rect 21252 29372 21262 29428
rect 23650 29372 23660 29428
rect 23716 29372 24332 29428
rect 24388 29372 24556 29428
rect 24612 29372 24622 29428
rect 24770 29372 24780 29428
rect 24836 29372 25564 29428
rect 25620 29372 25630 29428
rect 26002 29372 26012 29428
rect 26068 29372 26684 29428
rect 26740 29372 26750 29428
rect 41906 29372 41916 29428
rect 41972 29372 44492 29428
rect 44548 29372 44558 29428
rect 48738 29372 48748 29428
rect 48804 29372 49756 29428
rect 49812 29372 49822 29428
rect 50194 29372 50204 29428
rect 50260 29372 54908 29428
rect 54964 29372 54974 29428
rect 55122 29372 55132 29428
rect 55188 29372 55198 29428
rect 55458 29372 55468 29428
rect 55524 29372 56028 29428
rect 56084 29372 56094 29428
rect 56466 29372 56476 29428
rect 56532 29372 56542 29428
rect 56690 29372 56700 29428
rect 56756 29372 57260 29428
rect 57316 29372 59164 29428
rect 59220 29372 59230 29428
rect 55132 29316 55188 29372
rect 4162 29260 4172 29316
rect 4228 29260 4396 29316
rect 4452 29260 5852 29316
rect 5908 29260 6076 29316
rect 6132 29260 6142 29316
rect 6514 29260 6524 29316
rect 6580 29260 6636 29316
rect 6692 29260 6702 29316
rect 7158 29260 7196 29316
rect 7252 29260 7262 29316
rect 10994 29260 11004 29316
rect 11060 29260 12684 29316
rect 12740 29260 12750 29316
rect 12898 29260 12908 29316
rect 12964 29260 15596 29316
rect 15652 29260 21532 29316
rect 21588 29260 22428 29316
rect 22484 29260 22494 29316
rect 22754 29260 22764 29316
rect 22820 29260 24108 29316
rect 24164 29260 24892 29316
rect 24948 29260 24958 29316
rect 36530 29260 36540 29316
rect 36596 29260 47180 29316
rect 47236 29260 47246 29316
rect 47506 29260 47516 29316
rect 47572 29260 51324 29316
rect 51380 29260 51390 29316
rect 52434 29260 52444 29316
rect 52500 29260 53564 29316
rect 53620 29260 53630 29316
rect 55132 29260 55804 29316
rect 55860 29260 55870 29316
rect 12908 29204 12964 29260
rect 9538 29148 9548 29204
rect 9604 29148 9996 29204
rect 10052 29148 10780 29204
rect 10836 29148 12964 29204
rect 15698 29148 15708 29204
rect 15764 29148 16380 29204
rect 16436 29148 19628 29204
rect 19684 29148 19694 29204
rect 30258 29148 30268 29204
rect 30324 29148 31724 29204
rect 31780 29148 36092 29204
rect 36148 29148 36158 29204
rect 40786 29148 40796 29204
rect 40852 29148 41468 29204
rect 41524 29148 41692 29204
rect 41748 29148 41758 29204
rect 42690 29148 42700 29204
rect 42756 29148 43260 29204
rect 43316 29148 43596 29204
rect 43652 29148 43662 29204
rect 48626 29148 48636 29204
rect 48692 29148 49980 29204
rect 50036 29148 50046 29204
rect 51202 29148 51212 29204
rect 51268 29148 51436 29204
rect 51492 29148 51502 29204
rect 55570 29148 55580 29204
rect 55636 29148 56140 29204
rect 56196 29148 56206 29204
rect 5058 29036 5068 29092
rect 5124 29036 7420 29092
rect 7476 29036 7486 29092
rect 10434 29036 10444 29092
rect 10500 29036 20132 29092
rect 21858 29036 21868 29092
rect 21924 29036 33180 29092
rect 33236 29036 33246 29092
rect 36978 29036 36988 29092
rect 37044 29036 40572 29092
rect 40628 29036 40638 29092
rect 42354 29036 42364 29092
rect 42420 29036 42812 29092
rect 42868 29036 42878 29092
rect 46722 29036 46732 29092
rect 46788 29036 49644 29092
rect 49700 29036 49868 29092
rect 49924 29036 54684 29092
rect 54740 29036 54750 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 20076 28980 20132 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 6514 28924 6524 28980
rect 6580 28924 16604 28980
rect 16660 28924 16670 28980
rect 20076 28924 25116 28980
rect 25172 28924 25182 28980
rect 32498 28924 32508 28980
rect 32564 28924 34748 28980
rect 34804 28924 34814 28980
rect 37986 28924 37996 28980
rect 38052 28924 38556 28980
rect 38612 28924 38622 28980
rect 40786 28924 40796 28980
rect 40852 28924 41356 28980
rect 41412 28924 41422 28980
rect 44118 28924 44156 28980
rect 44212 28924 44222 28980
rect 48514 28924 48524 28980
rect 48580 28924 50988 28980
rect 51044 28924 51054 28980
rect 53004 28924 56028 28980
rect 56084 28924 56094 28980
rect 53004 28868 53060 28924
rect 3714 28812 3724 28868
rect 3780 28812 8428 28868
rect 8484 28812 8494 28868
rect 12002 28812 12012 28868
rect 12068 28812 12572 28868
rect 12628 28812 12638 28868
rect 15092 28812 16940 28868
rect 16996 28812 17006 28868
rect 22642 28812 22652 28868
rect 22708 28812 23660 28868
rect 23716 28812 27356 28868
rect 27412 28812 28588 28868
rect 28644 28812 28654 28868
rect 29698 28812 29708 28868
rect 29764 28812 31276 28868
rect 31332 28812 31342 28868
rect 32274 28812 32284 28868
rect 32340 28812 33068 28868
rect 33124 28812 33134 28868
rect 35074 28812 35084 28868
rect 35140 28812 38668 28868
rect 39330 28812 39340 28868
rect 39396 28812 45388 28868
rect 45444 28812 45454 28868
rect 47394 28812 47404 28868
rect 47460 28812 48860 28868
rect 48916 28812 48926 28868
rect 49868 28812 53060 28868
rect 53218 28812 53228 28868
rect 53284 28812 56756 28868
rect 15092 28756 15148 28812
rect 38612 28756 38668 28812
rect 49868 28756 49924 28812
rect 56700 28756 56756 28812
rect 7298 28700 7308 28756
rect 7364 28700 7402 28756
rect 9090 28700 9100 28756
rect 9156 28700 9996 28756
rect 10052 28700 11340 28756
rect 11396 28700 11406 28756
rect 13458 28700 13468 28756
rect 13524 28700 14252 28756
rect 14308 28700 15148 28756
rect 18162 28700 18172 28756
rect 18228 28700 21532 28756
rect 21588 28700 21598 28756
rect 21746 28700 21756 28756
rect 21812 28700 23100 28756
rect 23156 28700 23772 28756
rect 23828 28700 23838 28756
rect 27906 28700 27916 28756
rect 27972 28700 28700 28756
rect 28756 28700 28766 28756
rect 32162 28700 32172 28756
rect 32228 28700 33964 28756
rect 34020 28700 34030 28756
rect 34524 28700 35196 28756
rect 35252 28700 35644 28756
rect 35700 28700 36092 28756
rect 36148 28700 36540 28756
rect 36596 28700 36606 28756
rect 36754 28700 36764 28756
rect 36820 28700 37548 28756
rect 37604 28700 37614 28756
rect 38612 28700 39228 28756
rect 39284 28700 39564 28756
rect 39620 28700 39630 28756
rect 48850 28700 48860 28756
rect 48916 28700 49924 28756
rect 50082 28700 50092 28756
rect 50148 28700 55916 28756
rect 55972 28700 55982 28756
rect 56690 28700 56700 28756
rect 56756 28700 58044 28756
rect 58100 28700 59052 28756
rect 59108 28700 59118 28756
rect 34524 28644 34580 28700
rect 7196 28588 8428 28644
rect 8484 28588 8494 28644
rect 8642 28588 8652 28644
rect 8708 28588 10052 28644
rect 10210 28588 10220 28644
rect 10276 28588 11228 28644
rect 11284 28588 15484 28644
rect 15540 28588 15550 28644
rect 16034 28588 16044 28644
rect 16100 28588 18508 28644
rect 18564 28588 18574 28644
rect 20962 28588 20972 28644
rect 21028 28588 21588 28644
rect 23090 28588 23100 28644
rect 23156 28588 24668 28644
rect 24724 28588 24734 28644
rect 26674 28588 26684 28644
rect 26740 28588 28028 28644
rect 28084 28588 28094 28644
rect 30594 28588 30604 28644
rect 30660 28588 31052 28644
rect 31108 28588 31118 28644
rect 33506 28588 33516 28644
rect 33572 28588 34580 28644
rect 34738 28588 34748 28644
rect 34804 28588 35868 28644
rect 35924 28588 35934 28644
rect 36530 28588 36540 28644
rect 36596 28588 36606 28644
rect 38546 28588 38556 28644
rect 38612 28588 39676 28644
rect 39732 28588 40572 28644
rect 40628 28588 41804 28644
rect 41860 28588 41870 28644
rect 43586 28588 43596 28644
rect 43652 28588 44380 28644
rect 44436 28588 48300 28644
rect 48356 28588 48366 28644
rect 48626 28588 48636 28644
rect 48692 28588 48702 28644
rect 49970 28588 49980 28644
rect 50036 28588 50652 28644
rect 50708 28588 51660 28644
rect 51716 28588 51726 28644
rect 51986 28588 51996 28644
rect 52052 28588 52164 28644
rect 55346 28588 55356 28644
rect 55412 28588 57652 28644
rect 7196 28532 7252 28588
rect 9996 28532 10052 28588
rect 21532 28532 21588 28588
rect 7186 28476 7196 28532
rect 7252 28476 7262 28532
rect 9996 28476 11676 28532
rect 11732 28476 11742 28532
rect 21532 28476 22092 28532
rect 22148 28476 22540 28532
rect 22596 28476 22606 28532
rect 26338 28476 26348 28532
rect 26404 28476 27356 28532
rect 27412 28476 27422 28532
rect 29362 28476 29372 28532
rect 29428 28476 30268 28532
rect 30324 28476 31276 28532
rect 31332 28476 32172 28532
rect 32228 28476 32238 28532
rect 34514 28476 34524 28532
rect 34580 28476 35084 28532
rect 35140 28476 35150 28532
rect 36540 28420 36596 28588
rect 48636 28532 48692 28588
rect 52108 28532 52164 28588
rect 38612 28476 41580 28532
rect 41636 28476 41646 28532
rect 48626 28476 48636 28532
rect 48692 28476 49644 28532
rect 49700 28476 49710 28532
rect 51090 28476 51100 28532
rect 51156 28476 52052 28532
rect 52108 28476 54292 28532
rect 6066 28364 6076 28420
rect 6132 28364 7084 28420
rect 7140 28364 7150 28420
rect 9090 28364 9100 28420
rect 9156 28364 10108 28420
rect 10164 28364 12348 28420
rect 12404 28364 12414 28420
rect 14354 28364 14364 28420
rect 14420 28364 18060 28420
rect 18116 28364 18126 28420
rect 21410 28364 21420 28420
rect 21476 28364 23436 28420
rect 23492 28364 23502 28420
rect 25218 28364 25228 28420
rect 25284 28364 25900 28420
rect 25956 28364 26460 28420
rect 26516 28364 27132 28420
rect 27188 28364 27198 28420
rect 29586 28364 29596 28420
rect 29652 28364 31500 28420
rect 31556 28364 31566 28420
rect 35858 28364 35868 28420
rect 35924 28364 36596 28420
rect 38546 28364 38556 28420
rect 38612 28364 38668 28476
rect 50866 28364 50876 28420
rect 50932 28364 51772 28420
rect 51828 28364 51838 28420
rect 200 28308 800 28336
rect 12348 28308 12404 28364
rect 51996 28308 52052 28476
rect 54236 28420 54292 28476
rect 57596 28420 57652 28588
rect 52658 28364 52668 28420
rect 52724 28364 53564 28420
rect 53620 28364 53630 28420
rect 54236 28364 57148 28420
rect 57204 28364 57214 28420
rect 57586 28364 57596 28420
rect 57652 28364 57662 28420
rect 200 28252 1932 28308
rect 1988 28252 1998 28308
rect 3938 28252 3948 28308
rect 4004 28252 6300 28308
rect 6356 28252 6366 28308
rect 6626 28252 6636 28308
rect 6692 28252 9324 28308
rect 9380 28252 9390 28308
rect 9734 28252 9772 28308
rect 9828 28252 9838 28308
rect 12348 28252 14700 28308
rect 14756 28252 14766 28308
rect 15474 28252 15484 28308
rect 15540 28252 17724 28308
rect 17780 28252 18844 28308
rect 18900 28252 19292 28308
rect 19348 28252 19358 28308
rect 22194 28252 22204 28308
rect 22260 28252 23660 28308
rect 23716 28252 23726 28308
rect 29250 28252 29260 28308
rect 29316 28252 33628 28308
rect 33684 28252 33694 28308
rect 40114 28252 40124 28308
rect 40180 28252 40348 28308
rect 40404 28252 40414 28308
rect 43586 28252 43596 28308
rect 43652 28252 49868 28308
rect 49924 28252 50428 28308
rect 51986 28252 51996 28308
rect 52052 28252 52062 28308
rect 52770 28252 52780 28308
rect 52836 28252 53116 28308
rect 53172 28252 53182 28308
rect 54338 28252 54348 28308
rect 54404 28252 54460 28308
rect 54516 28252 54526 28308
rect 56214 28252 56252 28308
rect 56308 28252 56318 28308
rect 200 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 5180 28140 10780 28196
rect 10836 28140 10846 28196
rect 11442 28140 11452 28196
rect 11508 28140 13132 28196
rect 13188 28140 13198 28196
rect 14018 28140 14028 28196
rect 14084 28140 15820 28196
rect 15876 28140 15886 28196
rect 25330 28140 25340 28196
rect 25396 28140 25900 28196
rect 25956 28140 25966 28196
rect 33618 28140 33628 28196
rect 33684 28140 38444 28196
rect 38500 28140 40572 28196
rect 40628 28140 40638 28196
rect 40796 28140 48300 28196
rect 48356 28140 48366 28196
rect 48962 28140 48972 28196
rect 49028 28140 49420 28196
rect 49476 28140 49486 28196
rect 5180 28084 5236 28140
rect 40796 28084 40852 28140
rect 50372 28084 50428 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 51202 28140 51212 28196
rect 51268 28140 55804 28196
rect 55860 28140 55870 28196
rect 2370 28028 2380 28084
rect 2436 28028 2716 28084
rect 2772 28028 3724 28084
rect 3780 28028 3790 28084
rect 4834 28028 4844 28084
rect 4900 28028 5180 28084
rect 5236 28028 5246 28084
rect 6514 28028 6524 28084
rect 6580 28028 10220 28084
rect 10276 28028 10286 28084
rect 10658 28028 10668 28084
rect 10724 28028 14364 28084
rect 14420 28028 14430 28084
rect 16258 28028 16268 28084
rect 16324 28028 16940 28084
rect 16996 28028 17006 28084
rect 17948 28028 18396 28084
rect 18452 28028 19404 28084
rect 19460 28028 20636 28084
rect 20692 28028 20702 28084
rect 31042 28028 31052 28084
rect 31108 28028 31724 28084
rect 31780 28028 31790 28084
rect 32386 28028 32396 28084
rect 32452 28028 32620 28084
rect 32676 28028 33852 28084
rect 33908 28028 33918 28084
rect 34066 28028 34076 28084
rect 34132 28028 34170 28084
rect 37874 28028 37884 28084
rect 37940 28028 38444 28084
rect 38500 28028 38510 28084
rect 38658 28028 38668 28084
rect 38724 28028 39228 28084
rect 39284 28028 40852 28084
rect 41570 28028 41580 28084
rect 41636 28028 42252 28084
rect 42308 28028 42318 28084
rect 42700 28028 48076 28084
rect 48132 28028 48142 28084
rect 48402 28028 48412 28084
rect 48468 28028 49868 28084
rect 49924 28028 50092 28084
rect 50148 28028 50158 28084
rect 50372 28028 54460 28084
rect 54516 28028 55132 28084
rect 55188 28028 55198 28084
rect 56018 28028 56028 28084
rect 56084 28028 56812 28084
rect 56868 28028 56878 28084
rect 57138 28028 57148 28084
rect 57204 28028 57876 28084
rect 6524 27972 6580 28028
rect 17948 27972 18004 28028
rect 3154 27916 3164 27972
rect 3220 27916 6580 27972
rect 6636 27916 12012 27972
rect 12068 27916 12908 27972
rect 12964 27916 12974 27972
rect 13244 27916 15708 27972
rect 15764 27916 15774 27972
rect 16716 27916 18004 27972
rect 18162 27916 18172 27972
rect 18228 27916 22316 27972
rect 22372 27916 22764 27972
rect 22820 27916 22830 27972
rect 27234 27916 27244 27972
rect 27300 27916 28252 27972
rect 28308 27916 28318 27972
rect 34626 27916 34636 27972
rect 34692 27916 34972 27972
rect 35028 27916 35532 27972
rect 35588 27916 35756 27972
rect 35812 27916 39116 27972
rect 39172 27916 39182 27972
rect 40534 27916 40572 27972
rect 40628 27916 40638 27972
rect 6636 27860 6692 27916
rect 7868 27860 7924 27916
rect 13244 27860 13300 27916
rect 16716 27860 16772 27916
rect 42700 27860 42756 28028
rect 48412 27972 48468 28028
rect 56028 27972 56084 28028
rect 57820 27972 57876 28028
rect 44818 27916 44828 27972
rect 44884 27916 45164 27972
rect 45220 27916 45724 27972
rect 45780 27916 45790 27972
rect 46722 27916 46732 27972
rect 46788 27916 48468 27972
rect 50194 27916 50204 27972
rect 50260 27916 50764 27972
rect 50820 27916 50830 27972
rect 51874 27916 51884 27972
rect 51940 27916 54236 27972
rect 54292 27916 54302 27972
rect 54674 27916 54684 27972
rect 54740 27916 56084 27972
rect 56578 27916 56588 27972
rect 56644 27916 57484 27972
rect 57540 27916 57550 27972
rect 57810 27916 57820 27972
rect 57876 27916 58492 27972
rect 58548 27916 58558 27972
rect 3938 27804 3948 27860
rect 4004 27804 6692 27860
rect 6850 27804 6860 27860
rect 6916 27804 7196 27860
rect 7252 27804 7262 27860
rect 7410 27804 7420 27860
rect 7476 27804 7514 27860
rect 7858 27804 7868 27860
rect 7924 27804 7934 27860
rect 8092 27804 8764 27860
rect 8820 27804 10444 27860
rect 10500 27804 10510 27860
rect 12226 27804 12236 27860
rect 12292 27804 13020 27860
rect 13076 27804 13086 27860
rect 13234 27804 13244 27860
rect 13300 27804 13310 27860
rect 14242 27804 14252 27860
rect 14308 27804 14588 27860
rect 14644 27804 14654 27860
rect 15250 27804 15260 27860
rect 15316 27804 16716 27860
rect 16772 27804 16782 27860
rect 17042 27804 17052 27860
rect 17108 27804 18620 27860
rect 18676 27804 18686 27860
rect 19282 27804 19292 27860
rect 19348 27804 19740 27860
rect 19796 27804 19806 27860
rect 21634 27804 21644 27860
rect 21700 27804 24556 27860
rect 24612 27804 24622 27860
rect 36754 27804 36764 27860
rect 36820 27804 37436 27860
rect 37492 27804 37502 27860
rect 38658 27804 38668 27860
rect 38724 27804 42756 27860
rect 42914 27804 42924 27860
rect 42980 27804 47292 27860
rect 47348 27804 47740 27860
rect 47796 27804 47806 27860
rect 49634 27804 49644 27860
rect 49700 27804 50316 27860
rect 50372 27804 50382 27860
rect 3948 27748 4004 27804
rect 8092 27748 8148 27804
rect 14252 27748 14308 27804
rect 19292 27748 19348 27804
rect 51884 27748 51940 27916
rect 53106 27804 53116 27860
rect 53172 27804 53900 27860
rect 53956 27804 53966 27860
rect 1698 27692 1708 27748
rect 1764 27692 4004 27748
rect 4274 27692 4284 27748
rect 4340 27692 4396 27748
rect 4452 27692 4462 27748
rect 4946 27692 4956 27748
rect 5012 27692 5852 27748
rect 5908 27692 8148 27748
rect 8306 27692 8316 27748
rect 8372 27692 11788 27748
rect 11844 27692 12796 27748
rect 12852 27692 12862 27748
rect 13122 27692 13132 27748
rect 13188 27692 14308 27748
rect 17154 27692 17164 27748
rect 17220 27692 19348 27748
rect 20626 27692 20636 27748
rect 20692 27692 25004 27748
rect 25060 27692 25340 27748
rect 25396 27692 25406 27748
rect 37538 27692 37548 27748
rect 37604 27692 40908 27748
rect 40964 27692 41244 27748
rect 41300 27692 41310 27748
rect 42242 27692 42252 27748
rect 42308 27692 43596 27748
rect 43652 27692 43662 27748
rect 44706 27692 44716 27748
rect 44772 27692 45948 27748
rect 46004 27692 46014 27748
rect 46946 27692 46956 27748
rect 47012 27692 49308 27748
rect 49364 27692 51940 27748
rect 25340 27636 25396 27692
rect 42252 27636 42308 27692
rect 3602 27580 3612 27636
rect 3668 27580 6300 27636
rect 6356 27580 7420 27636
rect 7476 27580 9436 27636
rect 9492 27580 9502 27636
rect 9650 27580 9660 27636
rect 9716 27580 16044 27636
rect 16100 27580 16110 27636
rect 17714 27580 17724 27636
rect 17780 27580 19180 27636
rect 19236 27580 23100 27636
rect 23156 27580 23166 27636
rect 25340 27580 26460 27636
rect 26516 27580 26526 27636
rect 26786 27580 26796 27636
rect 26852 27580 28700 27636
rect 28756 27580 28766 27636
rect 36194 27580 36204 27636
rect 36260 27580 36764 27636
rect 36820 27580 36830 27636
rect 37202 27580 37212 27636
rect 37268 27580 37772 27636
rect 37828 27580 37838 27636
rect 38546 27580 38556 27636
rect 38612 27580 39788 27636
rect 39844 27580 41132 27636
rect 41188 27580 42308 27636
rect 43026 27580 43036 27636
rect 43092 27580 46844 27636
rect 46900 27580 52108 27636
rect 52164 27580 52174 27636
rect 54226 27580 54236 27636
rect 54292 27580 54348 27636
rect 54404 27580 54414 27636
rect 26852 27524 26908 27580
rect 5170 27468 5180 27524
rect 5236 27468 14028 27524
rect 14084 27468 14094 27524
rect 14354 27468 14364 27524
rect 14420 27468 26236 27524
rect 26292 27468 26908 27524
rect 39106 27468 39116 27524
rect 39172 27468 41468 27524
rect 41524 27468 43540 27524
rect 43670 27468 43708 27524
rect 43764 27468 43774 27524
rect 45378 27468 45388 27524
rect 45444 27468 45948 27524
rect 46004 27468 46014 27524
rect 48850 27468 48860 27524
rect 48916 27468 50204 27524
rect 50260 27468 50270 27524
rect 50642 27468 50652 27524
rect 50708 27468 54348 27524
rect 54404 27468 54414 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 43484 27412 43540 27468
rect 4946 27356 4956 27412
rect 5012 27356 8148 27412
rect 8390 27356 8428 27412
rect 8484 27356 8494 27412
rect 9874 27356 9884 27412
rect 9940 27356 12236 27412
rect 12292 27356 12302 27412
rect 12786 27356 12796 27412
rect 12852 27356 13356 27412
rect 13412 27356 13422 27412
rect 13570 27356 13580 27412
rect 13636 27356 14924 27412
rect 14980 27356 18844 27412
rect 18900 27356 20188 27412
rect 20244 27356 20860 27412
rect 20916 27356 20926 27412
rect 22082 27356 22092 27412
rect 22148 27356 24780 27412
rect 24836 27356 25676 27412
rect 25732 27356 25742 27412
rect 27906 27356 27916 27412
rect 27972 27356 28252 27412
rect 28308 27356 28318 27412
rect 31490 27356 31500 27412
rect 31556 27356 31724 27412
rect 31780 27356 31790 27412
rect 37986 27356 37996 27412
rect 38052 27356 38668 27412
rect 38724 27356 38734 27412
rect 41906 27356 41916 27412
rect 41972 27356 43428 27412
rect 43484 27356 46396 27412
rect 46452 27356 46462 27412
rect 48514 27356 48524 27412
rect 48580 27356 52668 27412
rect 52724 27356 52734 27412
rect 55906 27356 55916 27412
rect 55972 27356 56476 27412
rect 56532 27356 56542 27412
rect 3332 27244 7924 27300
rect 3332 27188 3388 27244
rect 1250 27132 1260 27188
rect 1316 27132 3164 27188
rect 3220 27132 3388 27188
rect 3490 27132 3500 27188
rect 3556 27132 3594 27188
rect 3826 27132 3836 27188
rect 3892 27132 4956 27188
rect 5012 27132 5022 27188
rect 6038 27132 6076 27188
rect 6132 27132 6142 27188
rect 2594 27020 2604 27076
rect 2660 27020 6860 27076
rect 6916 27020 7308 27076
rect 7364 27020 7374 27076
rect 2258 26908 2268 26964
rect 2324 26908 3612 26964
rect 3668 26908 4396 26964
rect 4452 26908 5740 26964
rect 5796 26908 5806 26964
rect 7868 26852 7924 27244
rect 8092 26964 8148 27356
rect 43372 27300 43428 27356
rect 8306 27244 8316 27300
rect 8372 27244 8382 27300
rect 11218 27244 11228 27300
rect 11284 27244 11676 27300
rect 11732 27244 14252 27300
rect 14308 27244 14318 27300
rect 16482 27244 16492 27300
rect 16548 27244 16716 27300
rect 16772 27244 18508 27300
rect 18564 27244 18574 27300
rect 19964 27244 21644 27300
rect 21700 27244 21710 27300
rect 22642 27244 22652 27300
rect 22708 27244 24780 27300
rect 24836 27244 27244 27300
rect 27300 27244 27310 27300
rect 30902 27244 30940 27300
rect 30996 27244 31006 27300
rect 34178 27244 34188 27300
rect 34244 27244 34524 27300
rect 34580 27244 34590 27300
rect 36642 27244 36652 27300
rect 36708 27244 39116 27300
rect 39172 27244 39182 27300
rect 43362 27244 43372 27300
rect 43428 27244 44268 27300
rect 44324 27244 47852 27300
rect 47908 27244 47918 27300
rect 51874 27244 51884 27300
rect 51940 27244 53004 27300
rect 53060 27244 53070 27300
rect 53526 27244 53564 27300
rect 53620 27244 53630 27300
rect 55794 27244 55804 27300
rect 55860 27244 56812 27300
rect 56868 27244 56878 27300
rect 8316 27188 8372 27244
rect 19964 27188 20020 27244
rect 8316 27132 12908 27188
rect 12964 27132 13468 27188
rect 13524 27132 13534 27188
rect 13794 27132 13804 27188
rect 13860 27132 16604 27188
rect 16660 27132 16670 27188
rect 18162 27132 18172 27188
rect 18228 27132 20020 27188
rect 20178 27132 20188 27188
rect 20244 27132 24724 27188
rect 24882 27132 24892 27188
rect 24948 27132 26124 27188
rect 26180 27132 28140 27188
rect 28196 27132 28700 27188
rect 28756 27132 28766 27188
rect 36418 27132 36428 27188
rect 36484 27132 36540 27188
rect 36596 27132 36606 27188
rect 37202 27132 37212 27188
rect 37268 27132 37324 27188
rect 37380 27132 37390 27188
rect 38210 27132 38220 27188
rect 38276 27132 39004 27188
rect 39060 27132 39070 27188
rect 40310 27132 40348 27188
rect 40404 27132 40414 27188
rect 41794 27132 41804 27188
rect 41860 27132 44492 27188
rect 44548 27132 44558 27188
rect 52294 27132 52332 27188
rect 52388 27132 52398 27188
rect 54310 27132 54348 27188
rect 54404 27132 54414 27188
rect 55234 27132 55244 27188
rect 55300 27132 57932 27188
rect 57988 27132 57998 27188
rect 24668 27076 24724 27132
rect 8306 27020 8316 27076
rect 8372 27020 14644 27076
rect 15362 27020 15372 27076
rect 15428 27020 17724 27076
rect 17780 27020 17790 27076
rect 18498 27020 18508 27076
rect 18564 27020 20860 27076
rect 20916 27020 21420 27076
rect 21476 27020 21486 27076
rect 24668 27020 25900 27076
rect 25956 27020 25966 27076
rect 26450 27020 26460 27076
rect 26516 27020 28588 27076
rect 28644 27020 28654 27076
rect 30146 27020 30156 27076
rect 30212 27020 31276 27076
rect 31332 27020 31342 27076
rect 35186 27020 35196 27076
rect 35252 27020 38444 27076
rect 38500 27020 38510 27076
rect 39218 27020 39228 27076
rect 39284 27020 42140 27076
rect 42196 27020 42206 27076
rect 43222 27020 43260 27076
rect 43316 27020 43326 27076
rect 43558 27020 43596 27076
rect 43652 27020 43662 27076
rect 44930 27020 44940 27076
rect 44996 27020 48524 27076
rect 48580 27020 48590 27076
rect 48748 27020 51212 27076
rect 51268 27020 51278 27076
rect 52098 27020 52108 27076
rect 52164 27020 54124 27076
rect 54180 27020 55580 27076
rect 55636 27020 55646 27076
rect 14588 26964 14644 27020
rect 42140 26964 42196 27020
rect 48748 26964 48804 27020
rect 8082 26908 8092 26964
rect 8148 26908 10332 26964
rect 10388 26908 10398 26964
rect 10770 26908 10780 26964
rect 10836 26908 11116 26964
rect 11172 26908 11182 26964
rect 12226 26908 12236 26964
rect 12292 26908 13580 26964
rect 13636 26908 13646 26964
rect 13794 26908 13804 26964
rect 13860 26908 13898 26964
rect 14578 26908 14588 26964
rect 14644 26908 19292 26964
rect 19348 26908 23324 26964
rect 23380 26908 23390 26964
rect 25442 26908 25452 26964
rect 25508 26908 26572 26964
rect 26628 26908 26638 26964
rect 27122 26908 27132 26964
rect 27188 26908 27580 26964
rect 27636 26908 27646 26964
rect 30258 26908 30268 26964
rect 30324 26908 30828 26964
rect 30884 26908 30894 26964
rect 32162 26908 32172 26964
rect 32228 26908 32732 26964
rect 32788 26908 32798 26964
rect 34402 26908 34412 26964
rect 34468 26908 36540 26964
rect 36596 26908 36606 26964
rect 37874 26908 37884 26964
rect 37940 26908 38332 26964
rect 38388 26908 38398 26964
rect 40450 26908 40460 26964
rect 40516 26908 41132 26964
rect 41188 26908 41198 26964
rect 42140 26908 42588 26964
rect 42644 26908 43372 26964
rect 43428 26908 43438 26964
rect 46722 26908 46732 26964
rect 46788 26908 46844 26964
rect 46900 26908 48804 26964
rect 49410 26908 49420 26964
rect 49476 26908 50428 26964
rect 50484 26908 50494 26964
rect 51314 26908 51324 26964
rect 51380 26908 51548 26964
rect 51604 26908 51614 26964
rect 54198 26908 54236 26964
rect 54292 26908 54302 26964
rect 54450 26908 54460 26964
rect 54516 26908 54526 26964
rect 54870 26908 54908 26964
rect 54964 26908 54974 26964
rect 55122 26908 55132 26964
rect 55188 26908 56028 26964
rect 56084 26908 57148 26964
rect 54460 26852 54516 26908
rect 2146 26796 2156 26852
rect 2212 26796 6860 26852
rect 6916 26796 7196 26852
rect 7252 26796 7262 26852
rect 7858 26796 7868 26852
rect 7924 26796 7934 26852
rect 15586 26796 15596 26852
rect 15652 26796 16604 26852
rect 16660 26796 16670 26852
rect 18582 26796 18620 26852
rect 18676 26796 18686 26852
rect 24098 26796 24108 26852
rect 24164 26796 25788 26852
rect 25844 26796 25854 26852
rect 28242 26796 28252 26852
rect 28308 26796 28476 26852
rect 28532 26796 28542 26852
rect 32386 26796 32396 26852
rect 32452 26796 33180 26852
rect 33236 26796 33246 26852
rect 35410 26796 35420 26852
rect 35476 26796 35486 26852
rect 38546 26796 38556 26852
rect 38612 26796 40236 26852
rect 40292 26796 40302 26852
rect 40674 26796 40684 26852
rect 40740 26796 40908 26852
rect 40964 26796 40974 26852
rect 43250 26796 43260 26852
rect 43316 26796 43708 26852
rect 43764 26796 43774 26852
rect 43922 26796 43932 26852
rect 43988 26796 43998 26852
rect 46946 26796 46956 26852
rect 47012 26796 47852 26852
rect 47908 26796 47918 26852
rect 50082 26796 50092 26852
rect 50148 26796 50204 26852
rect 50260 26796 50652 26852
rect 50708 26796 50718 26852
rect 52210 26796 52220 26852
rect 52276 26796 53676 26852
rect 53732 26796 53742 26852
rect 54338 26796 54348 26852
rect 54404 26796 54516 26852
rect 57092 26796 57148 26908
rect 57204 26796 57214 26852
rect 57474 26796 57484 26852
rect 57540 26796 57820 26852
rect 57876 26796 57886 26852
rect 35420 26740 35476 26796
rect 43932 26740 43988 26796
rect 2706 26684 2716 26740
rect 2772 26684 4844 26740
rect 4900 26684 4910 26740
rect 6962 26684 6972 26740
rect 7028 26684 7084 26740
rect 7140 26684 8428 26740
rect 8484 26684 8494 26740
rect 9314 26684 9324 26740
rect 9380 26684 11228 26740
rect 11284 26684 11294 26740
rect 11442 26684 11452 26740
rect 11508 26684 14924 26740
rect 14980 26684 17164 26740
rect 17220 26684 17836 26740
rect 17892 26684 17902 26740
rect 27794 26684 27804 26740
rect 27860 26684 28364 26740
rect 28420 26684 28430 26740
rect 35420 26684 35644 26740
rect 35700 26684 35710 26740
rect 38322 26684 38332 26740
rect 38388 26684 40684 26740
rect 40740 26684 40750 26740
rect 42130 26684 42140 26740
rect 42196 26684 42252 26740
rect 42308 26684 42318 26740
rect 42802 26684 42812 26740
rect 42868 26684 45164 26740
rect 45220 26684 45500 26740
rect 45556 26684 45566 26740
rect 46162 26684 46172 26740
rect 46228 26684 46620 26740
rect 46676 26684 46686 26740
rect 47394 26684 47404 26740
rect 47460 26684 48076 26740
rect 48132 26684 49532 26740
rect 49588 26684 49598 26740
rect 51314 26684 51324 26740
rect 51380 26684 51548 26740
rect 51604 26684 54460 26740
rect 54516 26684 54526 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 3490 26572 3500 26628
rect 3556 26572 4396 26628
rect 4452 26572 7196 26628
rect 7252 26572 7868 26628
rect 7924 26572 7934 26628
rect 8082 26572 8092 26628
rect 8148 26572 10444 26628
rect 10500 26572 10510 26628
rect 10658 26572 10668 26628
rect 10724 26572 12796 26628
rect 12852 26572 12862 26628
rect 35410 26572 35420 26628
rect 35476 26572 35980 26628
rect 36036 26572 36540 26628
rect 36596 26572 36606 26628
rect 40310 26572 40348 26628
rect 40404 26572 40414 26628
rect 41570 26572 41580 26628
rect 41636 26572 42364 26628
rect 42420 26572 42430 26628
rect 43334 26572 43372 26628
rect 43428 26572 43438 26628
rect 43820 26572 44268 26628
rect 44324 26572 49084 26628
rect 49140 26572 49150 26628
rect 51090 26572 51100 26628
rect 51156 26572 57708 26628
rect 57764 26572 57774 26628
rect 7868 26516 7924 26572
rect 43820 26516 43876 26572
rect 3798 26460 3836 26516
rect 3892 26460 3902 26516
rect 5730 26460 5740 26516
rect 5796 26460 6300 26516
rect 6356 26460 6366 26516
rect 6850 26460 6860 26516
rect 6916 26460 7532 26516
rect 7588 26460 7598 26516
rect 7868 26460 8316 26516
rect 8372 26460 8382 26516
rect 8530 26460 8540 26516
rect 8596 26460 9212 26516
rect 9268 26460 9278 26516
rect 12450 26460 12460 26516
rect 12516 26460 12908 26516
rect 12964 26460 12974 26516
rect 13132 26460 24108 26516
rect 24164 26460 24174 26516
rect 25106 26460 25116 26516
rect 25172 26460 27132 26516
rect 27188 26460 27198 26516
rect 28690 26460 28700 26516
rect 28756 26460 28924 26516
rect 28980 26460 28990 26516
rect 35532 26460 38892 26516
rect 38948 26460 38958 26516
rect 40450 26460 40460 26516
rect 40516 26460 41468 26516
rect 41524 26460 41534 26516
rect 41804 26460 43876 26516
rect 44006 26460 44044 26516
rect 44100 26460 44380 26516
rect 44436 26460 44446 26516
rect 44594 26460 44604 26516
rect 44660 26460 46620 26516
rect 46676 26460 50764 26516
rect 50820 26460 50830 26516
rect 13132 26404 13188 26460
rect 35532 26404 35588 26460
rect 41804 26404 41860 26460
rect 5394 26348 5404 26404
rect 5460 26348 13132 26404
rect 13188 26348 13198 26404
rect 14578 26348 14588 26404
rect 14644 26348 15596 26404
rect 15652 26348 15662 26404
rect 16482 26348 16492 26404
rect 16548 26348 20412 26404
rect 20468 26348 20478 26404
rect 23426 26348 23436 26404
rect 23492 26348 24332 26404
rect 24388 26348 24398 26404
rect 26226 26348 26236 26404
rect 26292 26348 29484 26404
rect 29540 26348 29550 26404
rect 32162 26348 32172 26404
rect 32228 26348 32508 26404
rect 32564 26348 32574 26404
rect 35522 26348 35532 26404
rect 35588 26348 35598 26404
rect 36726 26348 36764 26404
rect 36820 26348 36830 26404
rect 37986 26348 37996 26404
rect 38052 26348 38332 26404
rect 38388 26348 38668 26404
rect 38724 26348 38734 26404
rect 41570 26348 41580 26404
rect 41636 26348 41804 26404
rect 41860 26348 41870 26404
rect 42130 26348 42140 26404
rect 42196 26348 43820 26404
rect 43876 26348 43886 26404
rect 44706 26348 44716 26404
rect 44772 26348 45612 26404
rect 45668 26348 46060 26404
rect 46116 26348 46126 26404
rect 47702 26348 47740 26404
rect 47796 26348 47806 26404
rect 49186 26348 49196 26404
rect 49252 26348 50092 26404
rect 50148 26348 50316 26404
rect 50372 26348 50382 26404
rect 51650 26348 51660 26404
rect 51716 26348 53228 26404
rect 53284 26348 53294 26404
rect 1810 26236 1820 26292
rect 1876 26236 5740 26292
rect 5796 26236 6748 26292
rect 6804 26236 6814 26292
rect 7186 26236 7196 26292
rect 7252 26236 7980 26292
rect 8036 26236 8046 26292
rect 8418 26236 8428 26292
rect 8484 26236 10556 26292
rect 10612 26236 10622 26292
rect 11788 26236 14364 26292
rect 14420 26236 14430 26292
rect 17602 26236 17612 26292
rect 17668 26236 19404 26292
rect 19460 26236 19470 26292
rect 20514 26236 20524 26292
rect 20580 26236 22652 26292
rect 22708 26236 24892 26292
rect 24948 26236 24958 26292
rect 25666 26236 25676 26292
rect 25732 26236 26348 26292
rect 26404 26236 26414 26292
rect 27458 26236 27468 26292
rect 27524 26236 28476 26292
rect 28532 26236 28542 26292
rect 31490 26236 31500 26292
rect 31556 26236 32060 26292
rect 32116 26236 35644 26292
rect 35700 26236 35710 26292
rect 36390 26236 36428 26292
rect 36484 26236 36494 26292
rect 39078 26236 39116 26292
rect 39172 26236 39182 26292
rect 40562 26236 40572 26292
rect 40628 26236 47852 26292
rect 47908 26236 48076 26292
rect 48132 26236 49868 26292
rect 49924 26236 50204 26292
rect 50260 26236 50270 26292
rect 51062 26236 51100 26292
rect 51156 26236 51166 26292
rect 54786 26236 54796 26292
rect 54852 26236 54908 26292
rect 54964 26236 54974 26292
rect 8428 26180 8484 26236
rect 11788 26180 11844 26236
rect 2146 26124 2156 26180
rect 2212 26124 6748 26180
rect 6804 26124 6814 26180
rect 7410 26124 7420 26180
rect 7476 26124 8484 26180
rect 11778 26124 11788 26180
rect 11844 26124 11882 26180
rect 12198 26124 12236 26180
rect 12292 26124 12302 26180
rect 14466 26124 14476 26180
rect 14532 26124 17724 26180
rect 17780 26124 17790 26180
rect 18946 26124 18956 26180
rect 19012 26124 24276 26180
rect 26002 26124 26012 26180
rect 26068 26124 26236 26180
rect 26292 26124 26302 26180
rect 28578 26124 28588 26180
rect 28644 26124 29036 26180
rect 29092 26124 29102 26180
rect 31714 26124 31724 26180
rect 31780 26124 31948 26180
rect 32004 26124 32014 26180
rect 32610 26124 32620 26180
rect 32676 26124 33516 26180
rect 33572 26124 33582 26180
rect 33954 26124 33964 26180
rect 34020 26124 34412 26180
rect 34468 26124 37436 26180
rect 37492 26124 37502 26180
rect 37986 26124 37996 26180
rect 38052 26124 40012 26180
rect 40068 26124 40078 26180
rect 40786 26124 40796 26180
rect 40852 26124 41356 26180
rect 41412 26124 41422 26180
rect 41794 26124 41804 26180
rect 41860 26124 46620 26180
rect 46676 26124 46686 26180
rect 48524 26124 51660 26180
rect 51716 26124 51726 26180
rect 51986 26124 51996 26180
rect 52052 26124 53340 26180
rect 53396 26124 53406 26180
rect 54450 26124 54460 26180
rect 54516 26124 56588 26180
rect 56644 26124 56654 26180
rect 24220 26068 24276 26124
rect 40012 26068 40068 26124
rect 2482 26012 2492 26068
rect 2548 26012 8988 26068
rect 9044 26012 9884 26068
rect 9940 26012 9950 26068
rect 10882 26012 10892 26068
rect 10948 26012 15484 26068
rect 15540 26012 15550 26068
rect 16706 26012 16716 26068
rect 16772 26012 18508 26068
rect 18564 26012 20188 26068
rect 20244 26012 20254 26068
rect 24210 26012 24220 26068
rect 24276 26012 26572 26068
rect 26628 26012 30044 26068
rect 30100 26012 30110 26068
rect 33394 26012 33404 26068
rect 33460 26012 36428 26068
rect 36484 26012 36494 26068
rect 37762 26012 37772 26068
rect 37828 26012 39228 26068
rect 39284 26012 39294 26068
rect 40012 26012 42028 26068
rect 42084 26012 42094 26068
rect 42354 26012 42364 26068
rect 42420 26012 44604 26068
rect 44660 26012 44670 26068
rect 45602 26012 45612 26068
rect 45668 26012 48300 26068
rect 48356 26012 48366 26068
rect 16716 25956 16772 26012
rect 6738 25900 6748 25956
rect 6804 25900 7644 25956
rect 7700 25900 7710 25956
rect 7858 25900 7868 25956
rect 7924 25900 8652 25956
rect 8708 25900 9324 25956
rect 9380 25900 9390 25956
rect 9986 25900 9996 25956
rect 10052 25900 11564 25956
rect 11620 25900 11630 25956
rect 11788 25900 13804 25956
rect 13860 25900 13870 25956
rect 14354 25900 14364 25956
rect 14420 25900 16772 25956
rect 17490 25900 17500 25956
rect 17556 25900 23324 25956
rect 23380 25900 23390 25956
rect 27682 25900 27692 25956
rect 27748 25900 28252 25956
rect 28308 25900 28318 25956
rect 31266 25900 31276 25956
rect 31332 25900 31612 25956
rect 31668 25900 32284 25956
rect 32340 25900 32350 25956
rect 37650 25900 37660 25956
rect 37716 25900 38444 25956
rect 38500 25900 38510 25956
rect 39554 25900 39564 25956
rect 39620 25900 46172 25956
rect 46228 25900 46238 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 11788 25844 11844 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 48524 25844 48580 26124
rect 49074 26012 49084 26068
rect 49140 26012 51212 26068
rect 51268 26012 52220 26068
rect 52276 26012 52286 26068
rect 52770 26012 52780 26068
rect 52836 26012 56252 26068
rect 56308 26012 57932 26068
rect 57988 26012 57998 26068
rect 49746 25900 49756 25956
rect 49812 25900 51324 25956
rect 51380 25900 51390 25956
rect 52882 25900 52892 25956
rect 52948 25900 57820 25956
rect 57876 25900 58940 25956
rect 58996 25900 59006 25956
rect 5170 25788 5180 25844
rect 5236 25788 11844 25844
rect 12226 25788 12236 25844
rect 12292 25788 17948 25844
rect 18004 25788 18014 25844
rect 19506 25788 19516 25844
rect 19572 25788 19852 25844
rect 19908 25788 19918 25844
rect 36194 25788 36204 25844
rect 36260 25788 42140 25844
rect 42196 25788 42206 25844
rect 43810 25788 43820 25844
rect 43876 25788 48580 25844
rect 49186 25788 49196 25844
rect 49252 25788 50204 25844
rect 50260 25788 55356 25844
rect 55412 25788 55422 25844
rect 2594 25676 2604 25732
rect 2660 25676 2940 25732
rect 2996 25676 7420 25732
rect 7476 25676 7486 25732
rect 11442 25676 11452 25732
rect 11508 25676 12908 25732
rect 12964 25676 12974 25732
rect 16706 25676 16716 25732
rect 16772 25676 22652 25732
rect 22708 25676 23492 25732
rect 24882 25676 24892 25732
rect 24948 25676 25900 25732
rect 25956 25676 25966 25732
rect 35522 25676 35532 25732
rect 35588 25676 35868 25732
rect 35924 25676 35934 25732
rect 37650 25676 37660 25732
rect 37716 25676 43260 25732
rect 43316 25676 43326 25732
rect 44416 25676 44492 25732
rect 44548 25676 48748 25732
rect 48804 25676 48814 25732
rect 52994 25676 53004 25732
rect 53060 25676 53676 25732
rect 53732 25676 53742 25732
rect 23436 25620 23492 25676
rect 59200 25620 59800 25648
rect 1810 25564 1820 25620
rect 1876 25564 2268 25620
rect 2324 25564 2334 25620
rect 4386 25564 4396 25620
rect 4452 25564 4732 25620
rect 4788 25564 4798 25620
rect 4946 25564 4956 25620
rect 5012 25564 6076 25620
rect 6132 25564 6142 25620
rect 6598 25564 6636 25620
rect 6692 25564 6702 25620
rect 7186 25564 7196 25620
rect 7252 25564 7308 25620
rect 7364 25564 7374 25620
rect 7522 25564 7532 25620
rect 7588 25564 9660 25620
rect 9716 25564 9726 25620
rect 14466 25564 14476 25620
rect 14532 25564 16268 25620
rect 16324 25564 16334 25620
rect 16930 25564 16940 25620
rect 16996 25564 18956 25620
rect 19012 25564 19022 25620
rect 19170 25564 19180 25620
rect 19236 25564 19740 25620
rect 19796 25564 19806 25620
rect 22530 25564 22540 25620
rect 22596 25564 23212 25620
rect 23268 25564 23278 25620
rect 23436 25564 26236 25620
rect 26292 25564 26302 25620
rect 31042 25564 31052 25620
rect 31108 25564 32060 25620
rect 32116 25564 32126 25620
rect 36642 25564 36652 25620
rect 36708 25564 36988 25620
rect 37044 25564 38556 25620
rect 38612 25564 38622 25620
rect 40674 25564 40684 25620
rect 40740 25564 45612 25620
rect 45668 25564 45678 25620
rect 46620 25564 48972 25620
rect 49028 25564 49038 25620
rect 50372 25564 51884 25620
rect 51940 25564 51950 25620
rect 52098 25564 52108 25620
rect 52164 25564 52332 25620
rect 52388 25564 52398 25620
rect 53330 25564 53340 25620
rect 53396 25564 55524 25620
rect 56018 25564 56028 25620
rect 56084 25564 59800 25620
rect 46620 25508 46676 25564
rect 48972 25508 49028 25564
rect 50372 25508 50428 25564
rect 55468 25508 55524 25564
rect 59200 25536 59800 25564
rect 1922 25452 1932 25508
rect 1988 25452 7980 25508
rect 8036 25452 8046 25508
rect 9314 25452 9324 25508
rect 9380 25452 11452 25508
rect 11508 25452 11900 25508
rect 11956 25452 11966 25508
rect 13346 25452 13356 25508
rect 13412 25452 17276 25508
rect 17332 25452 17342 25508
rect 18722 25452 18732 25508
rect 18788 25452 19068 25508
rect 19124 25452 20860 25508
rect 20916 25452 23436 25508
rect 23492 25452 23502 25508
rect 33506 25452 33516 25508
rect 33572 25452 34412 25508
rect 34468 25452 36204 25508
rect 36260 25452 36270 25508
rect 36418 25452 36428 25508
rect 36484 25452 37772 25508
rect 37828 25452 37838 25508
rect 39554 25452 39564 25508
rect 39620 25452 40348 25508
rect 40404 25452 41468 25508
rect 41524 25452 41534 25508
rect 44902 25452 44940 25508
rect 44996 25452 45006 25508
rect 45826 25452 45836 25508
rect 45892 25452 46620 25508
rect 46676 25452 46686 25508
rect 48000 25452 48076 25508
rect 48132 25452 48412 25508
rect 48468 25452 48478 25508
rect 48972 25452 50428 25508
rect 51202 25452 51212 25508
rect 51268 25452 53452 25508
rect 53508 25452 53518 25508
rect 53666 25452 53676 25508
rect 53732 25452 55244 25508
rect 55300 25452 55310 25508
rect 55468 25452 56476 25508
rect 56532 25452 56588 25508
rect 56644 25452 56654 25508
rect 2818 25340 2828 25396
rect 2884 25340 7028 25396
rect 7186 25340 7196 25396
rect 7252 25340 7420 25396
rect 7476 25340 7486 25396
rect 7634 25340 7644 25396
rect 7700 25340 8428 25396
rect 8484 25340 8494 25396
rect 9548 25340 9996 25396
rect 10052 25340 13020 25396
rect 13076 25340 13860 25396
rect 13952 25340 14028 25396
rect 14084 25340 14476 25396
rect 14532 25340 14542 25396
rect 15092 25340 17052 25396
rect 17108 25340 17118 25396
rect 17714 25340 17724 25396
rect 17780 25340 23212 25396
rect 23268 25340 23278 25396
rect 25554 25340 25564 25396
rect 25620 25340 26012 25396
rect 26068 25340 26078 25396
rect 32274 25340 32284 25396
rect 32340 25340 34188 25396
rect 34244 25340 34254 25396
rect 34850 25340 34860 25396
rect 34916 25340 42924 25396
rect 42980 25340 42990 25396
rect 44146 25340 44156 25396
rect 44212 25340 45052 25396
rect 45108 25340 49084 25396
rect 49140 25340 49150 25396
rect 49522 25340 49532 25396
rect 49588 25340 56644 25396
rect 6972 25284 7028 25340
rect 9548 25284 9604 25340
rect 13804 25284 13860 25340
rect 15092 25284 15148 25340
rect 56588 25284 56644 25340
rect 2482 25228 2492 25284
rect 2548 25228 2884 25284
rect 3266 25228 3276 25284
rect 3332 25228 3948 25284
rect 4004 25228 4014 25284
rect 4162 25228 4172 25284
rect 4228 25228 5068 25284
rect 5124 25228 5134 25284
rect 5282 25228 5292 25284
rect 5348 25228 5740 25284
rect 5796 25228 5806 25284
rect 5964 25228 6748 25284
rect 6804 25228 6814 25284
rect 6972 25228 9100 25284
rect 9156 25228 9604 25284
rect 9762 25228 9772 25284
rect 9828 25228 9838 25284
rect 13804 25228 15148 25284
rect 16034 25228 16044 25284
rect 16100 25228 17052 25284
rect 17108 25228 18060 25284
rect 18116 25228 20076 25284
rect 20132 25228 20244 25284
rect 20514 25228 20524 25284
rect 20580 25228 21868 25284
rect 21924 25228 21934 25284
rect 24210 25228 24220 25284
rect 24276 25228 24892 25284
rect 24948 25228 24958 25284
rect 25218 25228 25228 25284
rect 25284 25228 26460 25284
rect 26516 25228 26796 25284
rect 26852 25228 27356 25284
rect 27412 25228 27422 25284
rect 29250 25228 29260 25284
rect 29316 25228 31724 25284
rect 31780 25228 31790 25284
rect 33394 25228 33404 25284
rect 33460 25228 33516 25284
rect 33572 25228 33582 25284
rect 35074 25228 35084 25284
rect 35140 25228 35644 25284
rect 35700 25228 35710 25284
rect 37090 25228 37100 25284
rect 37156 25228 37660 25284
rect 37716 25228 37726 25284
rect 38332 25228 38892 25284
rect 38948 25228 38958 25284
rect 39890 25228 39900 25284
rect 39956 25228 40460 25284
rect 40516 25228 40526 25284
rect 40982 25228 41020 25284
rect 41076 25228 41804 25284
rect 41860 25228 41870 25284
rect 42354 25228 42364 25284
rect 42420 25228 42476 25284
rect 42532 25228 42542 25284
rect 42802 25228 42812 25284
rect 42868 25228 42878 25284
rect 42998 25228 43036 25284
rect 43092 25228 43102 25284
rect 43260 25228 43932 25284
rect 43988 25228 43998 25284
rect 46050 25228 46060 25284
rect 46116 25228 47628 25284
rect 47684 25228 47694 25284
rect 48178 25228 48188 25284
rect 48244 25228 48254 25284
rect 48402 25228 48412 25284
rect 48468 25228 49868 25284
rect 49924 25228 49934 25284
rect 51314 25228 51324 25284
rect 51380 25228 51660 25284
rect 51716 25228 51726 25284
rect 52434 25228 52444 25284
rect 52500 25228 53676 25284
rect 53732 25228 53742 25284
rect 56578 25228 56588 25284
rect 56644 25228 56654 25284
rect 57698 25228 57708 25284
rect 57764 25228 58604 25284
rect 58660 25228 58670 25284
rect 2828 25172 2884 25228
rect 5964 25172 6020 25228
rect 9772 25172 9828 25228
rect 20188 25172 20244 25228
rect 38332 25172 38388 25228
rect 42812 25172 42868 25228
rect 43260 25172 43316 25228
rect 2818 25116 2828 25172
rect 2884 25116 2894 25172
rect 3714 25116 3724 25172
rect 3780 25116 6020 25172
rect 6336 25116 6412 25172
rect 6468 25116 7420 25172
rect 7476 25116 7486 25172
rect 7858 25116 7868 25172
rect 7924 25116 10444 25172
rect 10500 25116 11228 25172
rect 11284 25116 11294 25172
rect 12786 25116 12796 25172
rect 12852 25116 13916 25172
rect 13972 25116 13982 25172
rect 15250 25116 15260 25172
rect 15316 25116 15484 25172
rect 15540 25116 15932 25172
rect 15988 25116 15998 25172
rect 20188 25116 21980 25172
rect 22036 25116 22046 25172
rect 23090 25116 23100 25172
rect 23156 25116 25340 25172
rect 25396 25116 25406 25172
rect 28242 25116 28252 25172
rect 28308 25116 29372 25172
rect 29428 25116 29438 25172
rect 30930 25116 30940 25172
rect 30996 25116 31276 25172
rect 31332 25116 31342 25172
rect 36642 25116 36652 25172
rect 36708 25116 36764 25172
rect 36820 25116 36830 25172
rect 37174 25116 37212 25172
rect 37268 25116 37278 25172
rect 38322 25116 38332 25172
rect 38388 25116 38398 25172
rect 39442 25116 39452 25172
rect 39508 25116 40236 25172
rect 40292 25116 40302 25172
rect 42812 25116 43316 25172
rect 43586 25116 43596 25172
rect 43652 25116 43708 25172
rect 43764 25116 43774 25172
rect 46918 25116 46956 25172
rect 47012 25116 47022 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 48188 25060 48244 25228
rect 48514 25116 48524 25172
rect 48580 25116 49756 25172
rect 49812 25116 49822 25172
rect 54002 25116 54012 25172
rect 54068 25116 54796 25172
rect 54852 25116 54862 25172
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 2706 25004 2716 25060
rect 2772 25004 6076 25060
rect 6132 25004 7308 25060
rect 7364 25004 9772 25060
rect 9828 25004 9838 25060
rect 10098 25004 10108 25060
rect 10164 25004 15148 25060
rect 15204 25004 15708 25060
rect 15764 25004 15774 25060
rect 19282 25004 19292 25060
rect 19348 25004 19460 25060
rect 32498 25004 32508 25060
rect 32564 25004 36988 25060
rect 37044 25004 37324 25060
rect 37380 25004 37390 25060
rect 38612 25004 39228 25060
rect 39284 25004 39340 25060
rect 39396 25004 39406 25060
rect 43026 25004 43036 25060
rect 43092 25004 43372 25060
rect 43428 25004 43438 25060
rect 43596 25004 47404 25060
rect 47460 25004 47470 25060
rect 48188 25004 48972 25060
rect 49028 25004 49038 25060
rect 52322 25004 52332 25060
rect 52388 25004 54124 25060
rect 54180 25004 54190 25060
rect 57446 25004 57484 25060
rect 57540 25004 57550 25060
rect 19404 24948 19460 25004
rect 37324 24948 37380 25004
rect 38612 24948 38668 25004
rect 43596 24948 43652 25004
rect 3602 24892 3612 24948
rect 3668 24892 4284 24948
rect 4340 24892 4350 24948
rect 5058 24892 5068 24948
rect 5124 24892 11452 24948
rect 11508 24892 11518 24948
rect 11890 24892 11900 24948
rect 11956 24892 16380 24948
rect 16436 24892 16446 24948
rect 18946 24892 18956 24948
rect 19012 24892 19180 24948
rect 19236 24892 19246 24948
rect 19404 24892 21644 24948
rect 21700 24892 26068 24948
rect 28578 24892 28588 24948
rect 28644 24892 28924 24948
rect 28980 24892 29932 24948
rect 29988 24892 29998 24948
rect 32946 24892 32956 24948
rect 33012 24892 33404 24948
rect 33460 24892 34300 24948
rect 34356 24892 34366 24948
rect 37324 24892 38668 24948
rect 40898 24892 40908 24948
rect 40964 24892 41580 24948
rect 41636 24892 43652 24948
rect 46610 24892 46620 24948
rect 46676 24892 47964 24948
rect 48020 24892 48030 24948
rect 48178 24892 48188 24948
rect 48244 24892 51212 24948
rect 51268 24892 51278 24948
rect 54002 24892 54012 24948
rect 54068 24892 55692 24948
rect 55748 24892 55758 24948
rect 26012 24836 26068 24892
rect 4162 24780 4172 24836
rect 4228 24780 6076 24836
rect 6132 24780 6142 24836
rect 7270 24780 7308 24836
rect 7364 24780 7374 24836
rect 7522 24780 7532 24836
rect 7588 24780 7644 24836
rect 7700 24780 7710 24836
rect 9762 24780 9772 24836
rect 9828 24780 9884 24836
rect 9940 24780 15036 24836
rect 15092 24780 15102 24836
rect 15698 24780 15708 24836
rect 15764 24780 23100 24836
rect 23156 24780 24332 24836
rect 24388 24780 25564 24836
rect 25620 24780 25630 24836
rect 26002 24780 26012 24836
rect 26068 24780 26460 24836
rect 26516 24780 26526 24836
rect 26852 24780 27244 24836
rect 27300 24780 29484 24836
rect 29540 24780 29550 24836
rect 33730 24780 33740 24836
rect 33796 24780 34412 24836
rect 34468 24780 34636 24836
rect 34692 24780 35980 24836
rect 36036 24780 46732 24836
rect 46788 24780 46798 24836
rect 48066 24780 48076 24836
rect 48132 24780 48636 24836
rect 48692 24780 48702 24836
rect 49084 24780 55804 24836
rect 55860 24780 55870 24836
rect 26460 24724 26516 24780
rect 26852 24724 26908 24780
rect 2482 24668 2492 24724
rect 2548 24668 4284 24724
rect 4340 24668 4350 24724
rect 4806 24668 4844 24724
rect 4900 24668 4910 24724
rect 5506 24668 5516 24724
rect 5572 24668 6972 24724
rect 7028 24668 7038 24724
rect 7186 24668 7196 24724
rect 7252 24668 7756 24724
rect 7812 24668 7822 24724
rect 8418 24668 8428 24724
rect 8484 24668 9212 24724
rect 9268 24668 9278 24724
rect 10434 24668 10444 24724
rect 10500 24668 10892 24724
rect 10948 24668 10958 24724
rect 12786 24668 12796 24724
rect 12852 24668 15260 24724
rect 15316 24668 16716 24724
rect 16772 24668 16782 24724
rect 18162 24668 18172 24724
rect 18228 24668 18396 24724
rect 18452 24668 18462 24724
rect 18722 24668 18732 24724
rect 18788 24668 18956 24724
rect 19012 24668 19022 24724
rect 20850 24668 20860 24724
rect 20916 24668 23548 24724
rect 23604 24668 23614 24724
rect 26460 24668 26908 24724
rect 28242 24668 28252 24724
rect 28308 24668 29148 24724
rect 29204 24668 29214 24724
rect 35634 24668 35644 24724
rect 35700 24668 37548 24724
rect 37604 24668 38108 24724
rect 38164 24668 38174 24724
rect 44080 24668 44156 24724
rect 44212 24668 48860 24724
rect 48916 24668 48926 24724
rect 49084 24612 49140 24780
rect 49634 24668 49644 24724
rect 49700 24668 50316 24724
rect 50372 24668 51100 24724
rect 51156 24668 51166 24724
rect 53106 24668 53116 24724
rect 53172 24668 53564 24724
rect 53620 24668 57260 24724
rect 57316 24668 57326 24724
rect 3938 24556 3948 24612
rect 4004 24556 5964 24612
rect 6020 24556 6030 24612
rect 6290 24556 6300 24612
rect 6356 24556 10108 24612
rect 10164 24556 10174 24612
rect 13458 24556 13468 24612
rect 13524 24556 21028 24612
rect 28802 24556 28812 24612
rect 28868 24556 29260 24612
rect 29316 24556 29326 24612
rect 31154 24556 31164 24612
rect 31220 24556 31612 24612
rect 31668 24556 32172 24612
rect 32228 24556 33180 24612
rect 33236 24556 33246 24612
rect 34738 24556 34748 24612
rect 34804 24556 35532 24612
rect 35588 24556 36876 24612
rect 36932 24556 38780 24612
rect 38836 24556 38846 24612
rect 40124 24556 42812 24612
rect 42868 24556 42878 24612
rect 45154 24556 45164 24612
rect 45220 24556 49140 24612
rect 50754 24556 50764 24612
rect 50820 24556 51884 24612
rect 51940 24556 51950 24612
rect 3378 24444 3388 24500
rect 3444 24444 6188 24500
rect 6244 24444 6254 24500
rect 6412 24444 9324 24500
rect 9380 24444 9390 24500
rect 9986 24444 9996 24500
rect 10052 24444 19068 24500
rect 19124 24444 19134 24500
rect 19478 24444 19516 24500
rect 19572 24444 19582 24500
rect 6412 24388 6468 24444
rect 20972 24388 21028 24556
rect 40124 24500 40180 24556
rect 21634 24444 21644 24500
rect 21700 24444 23660 24500
rect 23716 24444 24332 24500
rect 24388 24444 24398 24500
rect 26114 24444 26124 24500
rect 26180 24444 32060 24500
rect 32116 24444 32126 24500
rect 33506 24444 33516 24500
rect 33572 24444 33852 24500
rect 33908 24444 35756 24500
rect 35812 24444 40180 24500
rect 40338 24444 40348 24500
rect 40404 24444 41916 24500
rect 41972 24444 43484 24500
rect 43540 24444 48076 24500
rect 48132 24444 48142 24500
rect 48290 24444 48300 24500
rect 48356 24444 48636 24500
rect 48692 24444 55132 24500
rect 55188 24444 55198 24500
rect 5954 24332 5964 24388
rect 6020 24332 6468 24388
rect 6626 24332 6636 24388
rect 6692 24332 8540 24388
rect 8596 24332 8606 24388
rect 9090 24332 9100 24388
rect 9156 24332 15260 24388
rect 15316 24332 15326 24388
rect 16034 24332 16044 24388
rect 16100 24332 18172 24388
rect 18228 24332 18238 24388
rect 18834 24332 18844 24388
rect 18900 24332 20300 24388
rect 20356 24332 20366 24388
rect 20972 24332 27020 24388
rect 27076 24332 30380 24388
rect 30436 24332 30446 24388
rect 41010 24332 41020 24388
rect 41076 24332 41804 24388
rect 41860 24332 41870 24388
rect 42354 24332 42364 24388
rect 42420 24332 43596 24388
rect 43652 24332 43662 24388
rect 47170 24332 47180 24388
rect 47236 24332 47740 24388
rect 47796 24332 47806 24388
rect 50306 24332 50316 24388
rect 50372 24332 52332 24388
rect 52388 24332 52398 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 3042 24220 3052 24276
rect 3108 24220 3612 24276
rect 3668 24220 3678 24276
rect 4844 24220 12012 24276
rect 12068 24220 12348 24276
rect 12404 24220 13468 24276
rect 13524 24220 13534 24276
rect 14466 24220 14476 24276
rect 14532 24220 14812 24276
rect 14868 24220 14878 24276
rect 15138 24220 15148 24276
rect 15204 24220 19068 24276
rect 19124 24220 19134 24276
rect 25302 24220 25340 24276
rect 25396 24220 25406 24276
rect 25778 24220 25788 24276
rect 25844 24220 30828 24276
rect 30884 24220 30894 24276
rect 37762 24220 37772 24276
rect 37828 24220 38220 24276
rect 38276 24220 51324 24276
rect 51380 24220 51390 24276
rect 4844 24164 4900 24220
rect 3154 24108 3164 24164
rect 3220 24108 3230 24164
rect 3714 24108 3724 24164
rect 3780 24108 4900 24164
rect 5842 24108 5852 24164
rect 5908 24108 6300 24164
rect 6356 24108 7980 24164
rect 8036 24108 8046 24164
rect 9090 24108 9100 24164
rect 9156 24108 9436 24164
rect 9492 24108 9502 24164
rect 11778 24108 11788 24164
rect 11844 24108 13804 24164
rect 13860 24108 13870 24164
rect 15138 24108 15148 24164
rect 15204 24108 16940 24164
rect 16996 24108 17276 24164
rect 17332 24108 18508 24164
rect 18564 24108 18574 24164
rect 19170 24108 19180 24164
rect 19236 24108 20300 24164
rect 20356 24108 20366 24164
rect 29810 24108 29820 24164
rect 29876 24108 31164 24164
rect 31220 24108 31230 24164
rect 40684 24108 42140 24164
rect 42196 24108 42206 24164
rect 42578 24108 42588 24164
rect 42644 24108 42700 24164
rect 42756 24108 44492 24164
rect 44548 24108 45836 24164
rect 45892 24108 45902 24164
rect 47954 24108 47964 24164
rect 48020 24108 49308 24164
rect 49364 24108 49374 24164
rect 49522 24108 49532 24164
rect 49588 24108 52444 24164
rect 52500 24108 52510 24164
rect 55906 24108 55916 24164
rect 55972 24108 57484 24164
rect 57540 24108 57550 24164
rect 3164 24052 3220 24108
rect 40684 24052 40740 24108
rect 2146 23996 2156 24052
rect 2212 23996 6580 24052
rect 8866 23996 8876 24052
rect 8932 23996 16940 24052
rect 16996 23996 17052 24052
rect 17108 23996 17118 24052
rect 17612 23996 18396 24052
rect 18452 23996 21308 24052
rect 21364 23996 26796 24052
rect 26852 23996 26862 24052
rect 31826 23996 31836 24052
rect 31892 23996 33292 24052
rect 33348 23996 33358 24052
rect 39330 23996 39340 24052
rect 39396 23996 40236 24052
rect 40292 23996 40302 24052
rect 40646 23996 40684 24052
rect 40740 23996 40750 24052
rect 41654 23996 41692 24052
rect 41748 23996 41758 24052
rect 42578 23996 42588 24052
rect 42644 23996 42700 24052
rect 42756 23996 42766 24052
rect 45490 23996 45500 24052
rect 45556 23996 48748 24052
rect 48804 23996 48814 24052
rect 49298 23996 49308 24052
rect 49364 23996 50876 24052
rect 50932 23996 50942 24052
rect 51538 23996 51548 24052
rect 51604 23996 54908 24052
rect 54964 23996 58044 24052
rect 58100 23996 58110 24052
rect 6524 23940 6580 23996
rect 17612 23940 17668 23996
rect 3154 23884 3164 23940
rect 3220 23884 4284 23940
rect 4340 23884 4844 23940
rect 4900 23884 4910 23940
rect 6514 23884 6524 23940
rect 6580 23884 6590 23940
rect 6710 23884 6748 23940
rect 6804 23884 6814 23940
rect 7186 23884 7196 23940
rect 7252 23884 7262 23940
rect 7410 23884 7420 23940
rect 7476 23884 8204 23940
rect 8260 23884 8270 23940
rect 9762 23884 9772 23940
rect 9828 23884 10668 23940
rect 10724 23884 10734 23940
rect 11554 23884 11564 23940
rect 11620 23884 11676 23940
rect 11732 23884 11742 23940
rect 13906 23884 13916 23940
rect 13972 23884 17668 23940
rect 19282 23884 19292 23940
rect 19348 23884 20804 23940
rect 23202 23884 23212 23940
rect 23268 23884 24108 23940
rect 24164 23884 24174 23940
rect 24770 23884 24780 23940
rect 24836 23884 25788 23940
rect 25844 23884 25854 23940
rect 31490 23884 31500 23940
rect 31556 23884 32284 23940
rect 32340 23884 32350 23940
rect 37202 23884 37212 23940
rect 37268 23884 38388 23940
rect 38882 23884 38892 23940
rect 38948 23884 43708 23940
rect 43764 23884 44044 23940
rect 44100 23884 44110 23940
rect 2370 23772 2380 23828
rect 2436 23772 3724 23828
rect 3780 23772 3790 23828
rect 6178 23772 6188 23828
rect 6244 23772 6254 23828
rect 2034 23660 2044 23716
rect 2100 23660 2268 23716
rect 2324 23660 2940 23716
rect 2996 23660 3006 23716
rect 3490 23660 3500 23716
rect 3556 23660 5068 23716
rect 5124 23660 5134 23716
rect 5954 23660 5964 23716
rect 6020 23660 6030 23716
rect 5964 23604 6020 23660
rect 6188 23604 6244 23772
rect 7196 23716 7252 23884
rect 20748 23828 20804 23884
rect 38332 23828 38388 23884
rect 45500 23828 45556 23996
rect 46162 23884 46172 23940
rect 46228 23884 48188 23940
rect 48244 23884 48254 23940
rect 52770 23884 52780 23940
rect 52836 23884 53452 23940
rect 53508 23884 53518 23940
rect 53890 23884 53900 23940
rect 53956 23884 56588 23940
rect 56644 23884 57484 23940
rect 57540 23884 57550 23940
rect 6972 23660 7252 23716
rect 7308 23772 9772 23828
rect 9828 23772 9838 23828
rect 9986 23772 9996 23828
rect 10052 23772 13636 23828
rect 13794 23772 13804 23828
rect 13860 23772 14700 23828
rect 14756 23772 14766 23828
rect 14914 23772 14924 23828
rect 14980 23772 17724 23828
rect 17780 23772 18060 23828
rect 18116 23772 18126 23828
rect 20738 23772 20748 23828
rect 20804 23772 23548 23828
rect 23604 23772 23772 23828
rect 23828 23772 23838 23828
rect 25330 23772 25340 23828
rect 25396 23772 26124 23828
rect 26180 23772 26190 23828
rect 26898 23772 26908 23828
rect 26964 23772 27244 23828
rect 27300 23772 28532 23828
rect 28690 23772 28700 23828
rect 28756 23772 29708 23828
rect 29764 23772 29932 23828
rect 29988 23772 29998 23828
rect 32722 23772 32732 23828
rect 32788 23772 33292 23828
rect 33348 23772 33358 23828
rect 33506 23772 33516 23828
rect 33572 23772 34300 23828
rect 34356 23772 34366 23828
rect 34626 23772 34636 23828
rect 34692 23772 37884 23828
rect 37940 23772 37950 23828
rect 38332 23772 39340 23828
rect 39396 23772 39406 23828
rect 41458 23772 41468 23828
rect 41524 23772 42588 23828
rect 42644 23772 42654 23828
rect 43148 23772 45556 23828
rect 47282 23772 47292 23828
rect 47348 23772 48412 23828
rect 48468 23772 48478 23828
rect 49298 23772 49308 23828
rect 49364 23772 49420 23828
rect 49476 23772 49486 23828
rect 50530 23772 50540 23828
rect 50596 23772 57204 23828
rect 2146 23548 2156 23604
rect 2212 23548 4284 23604
rect 4340 23548 6020 23604
rect 6178 23548 6188 23604
rect 6244 23548 6254 23604
rect 6738 23548 6748 23604
rect 6804 23548 6842 23604
rect 6972 23492 7028 23660
rect 7308 23604 7364 23772
rect 13580 23716 13636 23772
rect 28476 23716 28532 23772
rect 43148 23716 43204 23772
rect 57148 23716 57204 23772
rect 7522 23660 7532 23716
rect 7588 23660 7644 23716
rect 7700 23660 7710 23716
rect 8530 23660 8540 23716
rect 8596 23660 10220 23716
rect 10276 23660 10286 23716
rect 10434 23660 10444 23716
rect 10500 23660 11788 23716
rect 11844 23660 11854 23716
rect 13580 23660 14476 23716
rect 14532 23660 15148 23716
rect 15204 23660 15214 23716
rect 15558 23660 15596 23716
rect 15652 23660 15662 23716
rect 17826 23660 17836 23716
rect 17892 23660 20076 23716
rect 20132 23660 20300 23716
rect 20356 23660 20366 23716
rect 26012 23660 26236 23716
rect 26292 23660 26302 23716
rect 26786 23660 26796 23716
rect 26852 23660 27804 23716
rect 27860 23660 28252 23716
rect 28308 23660 28318 23716
rect 28476 23660 29484 23716
rect 29540 23660 29820 23716
rect 29876 23660 29886 23716
rect 35634 23660 35644 23716
rect 35700 23660 36540 23716
rect 36596 23660 36606 23716
rect 38070 23660 38108 23716
rect 38164 23660 38174 23716
rect 38294 23660 38332 23716
rect 38388 23660 38398 23716
rect 38770 23660 38780 23716
rect 38836 23660 39228 23716
rect 39284 23660 39294 23716
rect 42802 23660 42812 23716
rect 42868 23660 43148 23716
rect 43204 23660 43214 23716
rect 45490 23660 45500 23716
rect 45556 23660 47516 23716
rect 47572 23660 47582 23716
rect 48066 23660 48076 23716
rect 48132 23660 48636 23716
rect 48692 23660 48702 23716
rect 50194 23660 50204 23716
rect 50260 23660 50428 23716
rect 50484 23660 50494 23716
rect 50642 23660 50652 23716
rect 50708 23660 51324 23716
rect 51380 23660 51390 23716
rect 57138 23660 57148 23716
rect 57204 23660 59276 23716
rect 59332 23660 59342 23716
rect 26012 23604 26068 23660
rect 7196 23548 7364 23604
rect 7522 23548 7532 23604
rect 7588 23548 7868 23604
rect 7924 23548 7934 23604
rect 9986 23548 9996 23604
rect 10052 23548 10556 23604
rect 10612 23548 10622 23604
rect 15026 23548 15036 23604
rect 15092 23548 18564 23604
rect 26002 23548 26012 23604
rect 26068 23548 26078 23604
rect 30594 23548 30604 23604
rect 30660 23548 33460 23604
rect 33618 23548 33628 23604
rect 33684 23548 33964 23604
rect 34020 23548 34300 23604
rect 34356 23548 34524 23604
rect 34580 23548 34590 23604
rect 36418 23548 36428 23604
rect 36484 23548 36652 23604
rect 36708 23548 36718 23604
rect 36978 23548 36988 23604
rect 37044 23548 38444 23604
rect 38500 23548 39788 23604
rect 39844 23548 39854 23604
rect 45826 23548 45836 23604
rect 45892 23548 46396 23604
rect 46452 23548 46462 23604
rect 46834 23548 46844 23604
rect 46900 23548 47852 23604
rect 47908 23548 47918 23604
rect 7196 23492 7252 23548
rect 9996 23492 10052 23548
rect 6850 23436 6860 23492
rect 6916 23436 7028 23492
rect 7186 23436 7196 23492
rect 7252 23436 7262 23492
rect 7410 23436 7420 23492
rect 7476 23436 10052 23492
rect 13122 23436 13132 23492
rect 13188 23436 16044 23492
rect 16100 23436 16110 23492
rect 18508 23380 18564 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 33404 23492 33460 23548
rect 49522 23492 49532 23548
rect 49588 23492 49598 23548
rect 50082 23492 50092 23548
rect 50148 23492 50158 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 18918 23436 18956 23492
rect 19012 23436 19022 23492
rect 21746 23436 21756 23492
rect 21812 23436 25676 23492
rect 25732 23436 25742 23492
rect 33404 23436 33684 23492
rect 36306 23436 36316 23492
rect 36372 23436 37772 23492
rect 37828 23436 38668 23492
rect 40338 23436 40348 23492
rect 40404 23436 42476 23492
rect 42532 23436 42542 23492
rect 42690 23436 42700 23492
rect 42756 23436 47180 23492
rect 47236 23436 47246 23492
rect 47842 23436 47852 23492
rect 47908 23436 49084 23492
rect 49140 23436 49150 23492
rect 49298 23436 49308 23492
rect 49364 23436 49374 23492
rect 33628 23380 33684 23436
rect 38612 23380 38668 23436
rect 47852 23380 47908 23436
rect 3938 23324 3948 23380
rect 4004 23324 4014 23380
rect 4498 23324 4508 23380
rect 4564 23324 6076 23380
rect 6132 23324 7532 23380
rect 7588 23324 7598 23380
rect 13430 23324 13468 23380
rect 13524 23324 13534 23380
rect 15138 23324 15148 23380
rect 15204 23324 16716 23380
rect 16772 23324 16782 23380
rect 18508 23324 19516 23380
rect 19572 23324 20076 23380
rect 20132 23324 20142 23380
rect 25778 23324 25788 23380
rect 25844 23324 27916 23380
rect 27972 23324 28812 23380
rect 28868 23324 29484 23380
rect 29540 23324 29550 23380
rect 32610 23324 32620 23380
rect 32676 23324 33068 23380
rect 33124 23324 33134 23380
rect 33618 23324 33628 23380
rect 33684 23324 33694 23380
rect 35746 23324 35756 23380
rect 35812 23324 35822 23380
rect 37874 23324 37884 23380
rect 37940 23324 37950 23380
rect 38612 23324 39900 23380
rect 39956 23324 39966 23380
rect 40898 23324 40908 23380
rect 40964 23324 43036 23380
rect 43092 23324 43102 23380
rect 47282 23324 47292 23380
rect 47348 23324 47908 23380
rect 48514 23324 48524 23380
rect 48580 23324 48636 23380
rect 48692 23324 48702 23380
rect 3948 23268 4004 23324
rect 3948 23212 4396 23268
rect 4452 23212 14588 23268
rect 14644 23212 14654 23268
rect 15250 23212 15260 23268
rect 15316 23212 16044 23268
rect 16100 23212 18060 23268
rect 18116 23212 18126 23268
rect 19058 23212 19068 23268
rect 19124 23212 19516 23268
rect 19572 23212 22316 23268
rect 22372 23212 23436 23268
rect 23492 23212 23502 23268
rect 32386 23212 32396 23268
rect 32452 23212 32844 23268
rect 32900 23212 33404 23268
rect 33460 23212 33516 23268
rect 33572 23212 33582 23268
rect 3490 23100 3500 23156
rect 3556 23100 4060 23156
rect 4116 23100 4126 23156
rect 6626 23100 6636 23156
rect 6692 23100 7308 23156
rect 7364 23100 7374 23156
rect 14802 23100 14812 23156
rect 14868 23100 15148 23156
rect 15204 23100 15214 23156
rect 15698 23100 15708 23156
rect 15764 23100 16716 23156
rect 16772 23100 20636 23156
rect 20692 23100 20702 23156
rect 23212 23100 24892 23156
rect 24948 23100 24958 23156
rect 28438 23100 28476 23156
rect 28532 23100 28542 23156
rect 29026 23100 29036 23156
rect 29092 23100 29932 23156
rect 29988 23100 29998 23156
rect 23212 23044 23268 23100
rect 35756 23044 35812 23324
rect 37884 23268 37940 23324
rect 49308 23268 49364 23436
rect 37884 23212 40124 23268
rect 40180 23212 40190 23268
rect 40338 23212 40348 23268
rect 40404 23212 48188 23268
rect 48244 23212 48254 23268
rect 48972 23212 49364 23268
rect 48972 23156 49028 23212
rect 36082 23100 36092 23156
rect 36148 23100 41580 23156
rect 41636 23100 41646 23156
rect 42438 23100 42476 23156
rect 42532 23100 42542 23156
rect 43474 23100 43484 23156
rect 43540 23100 45052 23156
rect 45108 23100 45118 23156
rect 47394 23100 47404 23156
rect 47460 23100 49028 23156
rect 49532 23044 49588 23492
rect 50092 23436 50204 23492
rect 50260 23436 50270 23492
rect 51538 23436 51548 23492
rect 51604 23436 53676 23492
rect 53732 23436 53742 23492
rect 56914 23436 56924 23492
rect 56980 23436 57484 23492
rect 57540 23436 57550 23492
rect 50082 23324 50092 23380
rect 50148 23324 51100 23380
rect 51156 23324 51166 23380
rect 53442 23324 53452 23380
rect 53508 23324 54236 23380
rect 54292 23324 54302 23380
rect 55206 23324 55244 23380
rect 55300 23324 55310 23380
rect 57362 23324 57372 23380
rect 57428 23324 57708 23380
rect 57764 23324 57774 23380
rect 49746 23212 49756 23268
rect 49812 23212 50036 23268
rect 52406 23212 52444 23268
rect 52500 23212 52510 23268
rect 56018 23212 56028 23268
rect 56084 23212 56476 23268
rect 56532 23212 56542 23268
rect 49980 23156 50036 23212
rect 49980 23100 50204 23156
rect 50260 23100 50270 23156
rect 51314 23100 51324 23156
rect 51380 23100 53060 23156
rect 53442 23100 53452 23156
rect 53508 23100 54572 23156
rect 54628 23100 55580 23156
rect 55636 23100 57484 23156
rect 57540 23100 57550 23156
rect 1810 22988 1820 23044
rect 1876 22988 7196 23044
rect 7252 22988 7262 23044
rect 15586 22988 15596 23044
rect 15652 22988 16492 23044
rect 16548 22988 16558 23044
rect 17686 22988 17724 23044
rect 17780 22988 17790 23044
rect 18498 22988 18508 23044
rect 18564 22988 19404 23044
rect 19460 22988 19470 23044
rect 20402 22988 20412 23044
rect 20468 22988 22204 23044
rect 22260 22988 22270 23044
rect 22754 22988 22764 23044
rect 22820 22988 23212 23044
rect 23268 22988 23278 23044
rect 24210 22988 24220 23044
rect 24276 22988 26348 23044
rect 26404 22988 26414 23044
rect 32274 22988 32284 23044
rect 32340 22988 34636 23044
rect 34692 22988 34702 23044
rect 35532 22988 36988 23044
rect 37044 22988 37054 23044
rect 37874 22988 37884 23044
rect 37940 22988 39004 23044
rect 39060 22988 40684 23044
rect 40740 22988 40750 23044
rect 42130 22988 42140 23044
rect 42196 22988 43820 23044
rect 43876 22988 44380 23044
rect 44436 22988 44446 23044
rect 44818 22988 44828 23044
rect 44884 22988 49308 23044
rect 49364 22988 49374 23044
rect 49522 22988 49532 23044
rect 49588 22988 49598 23044
rect 50054 22988 50092 23044
rect 50148 22988 50158 23044
rect 50530 22988 50540 23044
rect 50596 22988 51884 23044
rect 51940 22988 51950 23044
rect 200 22932 800 22960
rect 20412 22932 20468 22988
rect 35532 22932 35588 22988
rect 53004 22932 53060 23100
rect 53190 22988 53228 23044
rect 53284 22988 53294 23044
rect 55122 22988 55132 23044
rect 55188 22988 55916 23044
rect 55972 22988 55982 23044
rect 56466 22988 56476 23044
rect 56532 22988 58828 23044
rect 58884 22988 58894 23044
rect 200 22876 1932 22932
rect 1988 22876 1998 22932
rect 2258 22876 2268 22932
rect 2324 22876 7420 22932
rect 7476 22876 7486 22932
rect 11778 22876 11788 22932
rect 11844 22876 11900 22932
rect 11956 22876 16548 22932
rect 16930 22876 16940 22932
rect 16996 22876 17612 22932
rect 17668 22876 20468 22932
rect 24322 22876 24332 22932
rect 24388 22876 25788 22932
rect 25844 22876 25854 22932
rect 32050 22876 32060 22932
rect 32116 22876 32956 22932
rect 33012 22876 33022 22932
rect 34514 22876 34524 22932
rect 34580 22876 35532 22932
rect 35588 22876 35598 22932
rect 36754 22876 36764 22932
rect 36820 22876 38556 22932
rect 38612 22876 38622 22932
rect 40114 22876 40124 22932
rect 40180 22876 46508 22932
rect 46564 22876 47068 22932
rect 47124 22876 47134 22932
rect 49568 22876 49644 22932
rect 49700 22876 52332 22932
rect 52388 22876 52398 22932
rect 53004 22876 56924 22932
rect 56980 22876 56990 22932
rect 200 22848 800 22876
rect 16492 22820 16548 22876
rect 4946 22764 4956 22820
rect 5012 22764 9100 22820
rect 9156 22764 9166 22820
rect 10770 22764 10780 22820
rect 10836 22764 12236 22820
rect 12292 22764 12302 22820
rect 16482 22764 16492 22820
rect 16548 22764 21196 22820
rect 21252 22764 23548 22820
rect 23604 22764 25564 22820
rect 25620 22764 25630 22820
rect 25890 22764 25900 22820
rect 25956 22764 26572 22820
rect 26628 22764 26638 22820
rect 36866 22764 36876 22820
rect 36932 22764 43260 22820
rect 43316 22764 43326 22820
rect 46050 22764 46060 22820
rect 46116 22764 47740 22820
rect 47796 22764 47806 22820
rect 49074 22764 49084 22820
rect 49140 22764 49980 22820
rect 50036 22764 57372 22820
rect 57428 22764 57438 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 4844 22652 12684 22708
rect 12740 22652 12750 22708
rect 14242 22652 14252 22708
rect 14308 22652 15372 22708
rect 15428 22652 15596 22708
rect 15652 22652 15662 22708
rect 15810 22652 15820 22708
rect 15876 22652 16604 22708
rect 16660 22652 17276 22708
rect 17332 22652 20860 22708
rect 20916 22652 20926 22708
rect 26422 22652 26460 22708
rect 26516 22652 26526 22708
rect 36950 22652 36988 22708
rect 37044 22652 37054 22708
rect 38098 22652 38108 22708
rect 38164 22652 38444 22708
rect 38500 22652 41692 22708
rect 41748 22652 41758 22708
rect 48178 22652 48188 22708
rect 48244 22652 52108 22708
rect 52164 22652 52174 22708
rect 4844 22596 4900 22652
rect 3602 22540 3612 22596
rect 3668 22540 4900 22596
rect 8530 22540 8540 22596
rect 8596 22540 10220 22596
rect 10276 22540 13468 22596
rect 13524 22540 16940 22596
rect 16996 22540 18956 22596
rect 19012 22540 19022 22596
rect 19170 22540 19180 22596
rect 19236 22540 26124 22596
rect 26180 22540 27020 22596
rect 27076 22540 27086 22596
rect 27234 22540 27244 22596
rect 27300 22540 28252 22596
rect 28308 22540 28700 22596
rect 28756 22540 29372 22596
rect 29428 22540 29932 22596
rect 29988 22540 29998 22596
rect 34738 22540 34748 22596
rect 34804 22540 35756 22596
rect 35812 22540 35822 22596
rect 42578 22540 42588 22596
rect 42644 22540 43708 22596
rect 43764 22540 43774 22596
rect 49746 22540 49756 22596
rect 49812 22540 51212 22596
rect 51268 22540 51278 22596
rect 51426 22540 51436 22596
rect 51492 22540 51548 22596
rect 51604 22540 51614 22596
rect 55430 22540 55468 22596
rect 55524 22540 55534 22596
rect 55682 22540 55692 22596
rect 55748 22540 56588 22596
rect 56644 22540 56654 22596
rect 19180 22484 19236 22540
rect 3714 22428 3724 22484
rect 3780 22428 5852 22484
rect 5908 22428 5918 22484
rect 6738 22428 6748 22484
rect 6804 22428 7084 22484
rect 7140 22428 7150 22484
rect 12562 22428 12572 22484
rect 12628 22428 15036 22484
rect 15092 22428 15102 22484
rect 15260 22428 17724 22484
rect 17780 22428 17790 22484
rect 18694 22428 18732 22484
rect 18788 22428 18798 22484
rect 19058 22428 19068 22484
rect 19124 22428 19236 22484
rect 19394 22428 19404 22484
rect 19460 22428 20636 22484
rect 20692 22428 20702 22484
rect 21074 22428 21084 22484
rect 21140 22428 21644 22484
rect 21700 22428 21710 22484
rect 26562 22428 26572 22484
rect 26628 22428 28140 22484
rect 28196 22428 28206 22484
rect 30706 22428 30716 22484
rect 30772 22428 31388 22484
rect 31444 22428 31892 22484
rect 15260 22372 15316 22428
rect 31836 22372 31892 22428
rect 38612 22372 38668 22484
rect 38724 22428 38734 22484
rect 40198 22428 40236 22484
rect 40292 22428 40302 22484
rect 41906 22428 41916 22484
rect 41972 22428 44380 22484
rect 44436 22428 50652 22484
rect 50708 22428 51996 22484
rect 52052 22428 52062 22484
rect 55766 22428 55804 22484
rect 55860 22428 55870 22484
rect 43372 22372 43428 22428
rect 51212 22372 51268 22428
rect 2370 22316 2380 22372
rect 2436 22316 2828 22372
rect 2884 22316 2894 22372
rect 3938 22316 3948 22372
rect 4004 22316 4956 22372
rect 5012 22316 5022 22372
rect 6290 22316 6300 22372
rect 6356 22316 6412 22372
rect 6468 22316 6478 22372
rect 6626 22316 6636 22372
rect 6692 22316 6972 22372
rect 7028 22316 7038 22372
rect 7410 22316 7420 22372
rect 7476 22316 8428 22372
rect 8484 22316 10332 22372
rect 10388 22316 10398 22372
rect 11106 22316 11116 22372
rect 11172 22316 15316 22372
rect 16482 22316 16492 22372
rect 16548 22316 21868 22372
rect 21924 22316 21934 22372
rect 22866 22316 22876 22372
rect 22932 22316 28588 22372
rect 28644 22316 29596 22372
rect 29652 22316 29662 22372
rect 31826 22316 31836 22372
rect 31892 22316 31902 22372
rect 36418 22316 36428 22372
rect 36484 22316 37660 22372
rect 37716 22316 37726 22372
rect 37874 22316 37884 22372
rect 37940 22316 38668 22372
rect 40002 22316 40012 22372
rect 40068 22316 40348 22372
rect 40404 22316 40908 22372
rect 40964 22316 40974 22372
rect 43362 22316 43372 22372
rect 43428 22316 43438 22372
rect 44482 22316 44492 22372
rect 44548 22316 44558 22372
rect 45490 22316 45500 22372
rect 45556 22316 47292 22372
rect 47348 22316 47358 22372
rect 47618 22316 47628 22372
rect 47684 22316 48636 22372
rect 48692 22316 48702 22372
rect 48962 22316 48972 22372
rect 49028 22316 50316 22372
rect 50372 22316 50382 22372
rect 51202 22316 51212 22372
rect 51268 22316 51278 22372
rect 51426 22316 51436 22372
rect 51492 22316 52332 22372
rect 52388 22316 52556 22372
rect 52612 22316 52622 22372
rect 54674 22316 54684 22372
rect 54740 22316 55020 22372
rect 55076 22316 55086 22372
rect 44492 22260 44548 22316
rect 47628 22260 47684 22316
rect 3042 22204 3052 22260
rect 3108 22204 3836 22260
rect 3892 22204 3902 22260
rect 5842 22204 5852 22260
rect 5908 22204 14252 22260
rect 14308 22204 14318 22260
rect 15026 22204 15036 22260
rect 15092 22204 19628 22260
rect 19684 22204 19694 22260
rect 20626 22204 20636 22260
rect 20692 22204 21756 22260
rect 21812 22204 24276 22260
rect 25890 22204 25900 22260
rect 25956 22204 25966 22260
rect 28802 22204 28812 22260
rect 28868 22204 30156 22260
rect 30212 22204 30604 22260
rect 30660 22204 30670 22260
rect 33478 22204 33516 22260
rect 33572 22204 33582 22260
rect 36642 22204 36652 22260
rect 36708 22204 37996 22260
rect 38052 22204 38062 22260
rect 38480 22204 38556 22260
rect 38612 22204 40460 22260
rect 40516 22204 41132 22260
rect 41188 22204 41198 22260
rect 41468 22204 44716 22260
rect 44772 22204 44782 22260
rect 45266 22204 45276 22260
rect 45332 22204 45836 22260
rect 45892 22204 46620 22260
rect 46676 22204 46686 22260
rect 47058 22204 47068 22260
rect 47124 22204 47684 22260
rect 48402 22204 48412 22260
rect 48468 22204 48524 22260
rect 48580 22204 48590 22260
rect 49298 22204 49308 22260
rect 49364 22204 50540 22260
rect 50596 22204 50606 22260
rect 50754 22204 50764 22260
rect 50820 22204 52444 22260
rect 52500 22204 52780 22260
rect 52836 22204 52846 22260
rect 56886 22204 56924 22260
rect 56980 22204 56990 22260
rect 6738 22092 6748 22148
rect 6804 22092 7644 22148
rect 7700 22092 10108 22148
rect 10164 22092 10174 22148
rect 10434 22092 10444 22148
rect 10500 22092 11228 22148
rect 11284 22092 11294 22148
rect 13906 22092 13916 22148
rect 13972 22092 14588 22148
rect 14644 22092 14654 22148
rect 15698 22092 15708 22148
rect 15764 22092 17108 22148
rect 17826 22092 17836 22148
rect 17892 22092 18508 22148
rect 18564 22092 18574 22148
rect 18722 22092 18732 22148
rect 18788 22092 19180 22148
rect 19236 22092 19246 22148
rect 21298 22092 21308 22148
rect 21364 22092 21980 22148
rect 22036 22092 22046 22148
rect 17052 22036 17108 22092
rect 24220 22036 24276 22204
rect 4172 21980 8988 22036
rect 9044 21980 11116 22036
rect 11172 21980 11182 22036
rect 13234 21980 13244 22036
rect 13300 21980 13636 22036
rect 16034 21980 16044 22036
rect 16100 21980 16828 22036
rect 16884 21980 16894 22036
rect 17052 21980 19180 22036
rect 19236 21980 19246 22036
rect 21858 21980 21868 22036
rect 21924 21980 23660 22036
rect 23716 21980 23726 22036
rect 24210 21980 24220 22036
rect 24276 21980 25676 22036
rect 25732 21980 25742 22036
rect 4172 21924 4228 21980
rect 13580 21924 13636 21980
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 4162 21868 4172 21924
rect 4228 21868 4238 21924
rect 5842 21868 5852 21924
rect 5908 21868 8092 21924
rect 8148 21868 8158 21924
rect 9202 21868 9212 21924
rect 9268 21868 9772 21924
rect 9828 21868 9838 21924
rect 10770 21868 10780 21924
rect 10836 21868 13356 21924
rect 13412 21868 13422 21924
rect 13580 21868 15372 21924
rect 15428 21868 15820 21924
rect 15876 21868 15886 21924
rect 23314 21868 23324 21924
rect 23380 21868 24108 21924
rect 24164 21868 24174 21924
rect 25900 21812 25956 22204
rect 41468 22148 41524 22204
rect 48412 22148 48468 22204
rect 32834 22092 32844 22148
rect 32900 22092 33180 22148
rect 33236 22092 35644 22148
rect 35700 22092 36204 22148
rect 36260 22092 37436 22148
rect 37492 22092 37502 22148
rect 37986 22092 37996 22148
rect 38052 22092 38108 22148
rect 38164 22092 38174 22148
rect 39442 22092 39452 22148
rect 39508 22092 40012 22148
rect 40068 22092 40078 22148
rect 40226 22092 40236 22148
rect 40292 22092 41524 22148
rect 41682 22092 41692 22148
rect 41748 22092 48468 22148
rect 49718 22092 49756 22148
rect 49812 22092 49822 22148
rect 50082 22092 50092 22148
rect 50148 22092 50428 22148
rect 50484 22092 50494 22148
rect 51202 22092 51212 22148
rect 51268 22092 53788 22148
rect 53844 22092 53854 22148
rect 55682 22092 55692 22148
rect 55748 22092 56700 22148
rect 56756 22092 56766 22148
rect 32050 21980 32060 22036
rect 32116 21980 32732 22036
rect 32788 21980 34972 22036
rect 35028 21980 35038 22036
rect 37996 21924 38052 22092
rect 38322 21980 38332 22036
rect 38388 21980 45276 22036
rect 45332 21980 45342 22036
rect 47170 21980 47180 22036
rect 47236 21980 48188 22036
rect 48244 21980 48254 22036
rect 50978 21980 50988 22036
rect 51044 21980 51436 22036
rect 51492 21980 51502 22036
rect 51650 21980 51660 22036
rect 51716 21980 51754 22036
rect 51986 21980 51996 22036
rect 52052 21980 52090 22036
rect 52220 21980 55916 22036
rect 55972 21980 57372 22036
rect 57428 21980 59052 22036
rect 59108 21980 59118 22036
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 51996 21924 52052 21980
rect 27794 21868 27804 21924
rect 27860 21868 27870 21924
rect 34066 21868 34076 21924
rect 34132 21868 34524 21924
rect 34580 21868 34590 21924
rect 37324 21868 38052 21924
rect 40534 21868 40572 21924
rect 40628 21868 40638 21924
rect 41458 21868 41468 21924
rect 41524 21868 41692 21924
rect 41748 21868 41758 21924
rect 44706 21868 44716 21924
rect 44772 21868 45948 21924
rect 46004 21868 46014 21924
rect 46386 21868 46396 21924
rect 46452 21868 47068 21924
rect 48178 21868 48188 21924
rect 48244 21868 49420 21924
rect 49476 21868 49486 21924
rect 51090 21868 51100 21924
rect 51156 21868 52052 21924
rect 27804 21812 27860 21868
rect 37324 21812 37380 21868
rect 47012 21812 47068 21868
rect 52220 21812 52276 21980
rect 7970 21756 7980 21812
rect 8036 21756 8316 21812
rect 8372 21756 8382 21812
rect 14130 21756 14140 21812
rect 14196 21756 17500 21812
rect 17556 21756 17566 21812
rect 18162 21756 18172 21812
rect 18228 21756 18732 21812
rect 18788 21756 18798 21812
rect 20066 21756 20076 21812
rect 20132 21756 23884 21812
rect 23940 21756 23950 21812
rect 24406 21756 24444 21812
rect 24500 21756 24510 21812
rect 25900 21756 26012 21812
rect 26068 21756 26078 21812
rect 26450 21756 26460 21812
rect 26516 21756 27860 21812
rect 28466 21756 28476 21812
rect 28532 21756 30828 21812
rect 30884 21756 30894 21812
rect 31266 21756 31276 21812
rect 31332 21756 32732 21812
rect 32788 21756 32798 21812
rect 35942 21756 35980 21812
rect 36036 21756 36046 21812
rect 36642 21756 36652 21812
rect 36708 21756 37380 21812
rect 37538 21756 37548 21812
rect 37604 21756 41916 21812
rect 41972 21756 44156 21812
rect 44212 21756 44222 21812
rect 47012 21756 47404 21812
rect 47460 21756 47470 21812
rect 48290 21756 48300 21812
rect 48356 21756 49644 21812
rect 49700 21756 49710 21812
rect 50530 21756 50540 21812
rect 50596 21756 50988 21812
rect 51044 21756 51054 21812
rect 51762 21756 51772 21812
rect 51828 21756 52276 21812
rect 52332 21868 54236 21924
rect 54292 21868 54302 21924
rect 52332 21700 52388 21868
rect 1586 21644 1596 21700
rect 1652 21644 2828 21700
rect 2884 21644 3164 21700
rect 3220 21644 3230 21700
rect 6402 21644 6412 21700
rect 6468 21644 12908 21700
rect 12964 21644 12974 21700
rect 15092 21644 15708 21700
rect 15764 21644 15774 21700
rect 17042 21644 17052 21700
rect 17108 21644 18060 21700
rect 18116 21644 18126 21700
rect 18498 21644 18508 21700
rect 18564 21644 21308 21700
rect 21364 21644 21374 21700
rect 21634 21644 21644 21700
rect 21700 21644 22092 21700
rect 22148 21644 22158 21700
rect 22278 21644 22316 21700
rect 22372 21644 22382 21700
rect 23650 21644 23660 21700
rect 23716 21644 26684 21700
rect 26740 21644 27804 21700
rect 27860 21644 27870 21700
rect 30006 21644 30044 21700
rect 30100 21644 30110 21700
rect 33394 21644 33404 21700
rect 33460 21644 34076 21700
rect 34132 21644 37100 21700
rect 37156 21644 37166 21700
rect 37772 21644 38108 21700
rect 38164 21644 38174 21700
rect 42578 21644 42588 21700
rect 42644 21644 44156 21700
rect 44212 21644 44222 21700
rect 47012 21644 47740 21700
rect 47796 21644 47806 21700
rect 47954 21644 47964 21700
rect 48020 21644 52388 21700
rect 53218 21644 53228 21700
rect 53284 21644 55244 21700
rect 55300 21644 56364 21700
rect 56420 21644 56430 21700
rect 15092 21588 15148 21644
rect 37772 21588 37828 21644
rect 47012 21588 47068 21644
rect 2706 21532 2716 21588
rect 2772 21532 3276 21588
rect 3332 21532 4508 21588
rect 4564 21532 4574 21588
rect 7186 21532 7196 21588
rect 7252 21532 7262 21588
rect 7858 21532 7868 21588
rect 7924 21532 7980 21588
rect 8036 21532 8046 21588
rect 8866 21532 8876 21588
rect 8932 21532 12124 21588
rect 12180 21532 12190 21588
rect 13346 21532 13356 21588
rect 13412 21532 14700 21588
rect 14756 21532 15148 21588
rect 15362 21532 15372 21588
rect 15428 21532 16156 21588
rect 16212 21532 16940 21588
rect 16996 21532 19404 21588
rect 19460 21532 20524 21588
rect 20580 21532 20590 21588
rect 22754 21532 22764 21588
rect 22820 21532 23324 21588
rect 23380 21532 23390 21588
rect 24322 21532 24332 21588
rect 24388 21532 24444 21588
rect 24500 21532 24510 21588
rect 26562 21532 26572 21588
rect 26628 21532 27580 21588
rect 27636 21532 27646 21588
rect 28914 21532 28924 21588
rect 28980 21532 29260 21588
rect 29316 21532 31276 21588
rect 31332 21532 31342 21588
rect 33954 21532 33964 21588
rect 34020 21532 34412 21588
rect 34468 21532 34478 21588
rect 35970 21532 35980 21588
rect 36036 21532 37772 21588
rect 37828 21532 37838 21588
rect 37986 21532 37996 21588
rect 38052 21532 38500 21588
rect 40114 21532 40124 21588
rect 40180 21532 40348 21588
rect 40404 21532 42476 21588
rect 42532 21532 42542 21588
rect 44034 21532 44044 21588
rect 44100 21532 46172 21588
rect 46228 21532 47068 21588
rect 47440 21532 47516 21588
rect 47572 21532 48300 21588
rect 48356 21532 48366 21588
rect 49298 21532 49308 21588
rect 49364 21532 50204 21588
rect 50260 21532 50540 21588
rect 50596 21532 50606 21588
rect 50866 21532 50876 21588
rect 50932 21532 53452 21588
rect 53508 21532 53518 21588
rect 53778 21532 53788 21588
rect 53844 21532 55692 21588
rect 55748 21532 55758 21588
rect 56690 21532 56700 21588
rect 56756 21532 57260 21588
rect 57316 21532 57596 21588
rect 57652 21532 57662 21588
rect 7196 21476 7252 21532
rect 12124 21476 12180 21532
rect 3490 21420 3500 21476
rect 3556 21420 4956 21476
rect 5012 21420 5022 21476
rect 6962 21420 6972 21476
rect 7028 21420 7644 21476
rect 7700 21420 7710 21476
rect 7970 21420 7980 21476
rect 8036 21420 9996 21476
rect 10052 21420 10062 21476
rect 12124 21420 13580 21476
rect 13636 21420 13646 21476
rect 16594 21420 16604 21476
rect 16660 21420 18732 21476
rect 18788 21420 19068 21476
rect 19124 21420 19134 21476
rect 21746 21420 21756 21476
rect 21812 21420 24892 21476
rect 24948 21420 24958 21476
rect 26898 21420 26908 21476
rect 26964 21420 28028 21476
rect 28084 21420 28094 21476
rect 35410 21420 35420 21476
rect 35476 21420 36652 21476
rect 36708 21420 36718 21476
rect 37202 21420 37212 21476
rect 37268 21420 38108 21476
rect 38164 21420 38174 21476
rect 24892 21364 24948 21420
rect 38444 21364 38500 21532
rect 38966 21420 39004 21476
rect 39060 21420 39340 21476
rect 39396 21420 39406 21476
rect 40562 21420 40572 21476
rect 40628 21420 42140 21476
rect 42196 21420 42588 21476
rect 42644 21420 42654 21476
rect 43922 21420 43932 21476
rect 43988 21420 48188 21476
rect 48244 21420 48254 21476
rect 48626 21420 48636 21476
rect 48692 21420 49924 21476
rect 51090 21420 51100 21476
rect 51156 21420 52668 21476
rect 52724 21420 52734 21476
rect 53264 21420 53340 21476
rect 53396 21420 53676 21476
rect 53732 21420 53742 21476
rect 54646 21420 54684 21476
rect 54740 21420 54750 21476
rect 49868 21364 49924 21420
rect 2258 21308 2268 21364
rect 2324 21308 6972 21364
rect 7028 21308 8092 21364
rect 8148 21308 8158 21364
rect 13010 21308 13020 21364
rect 13076 21308 16044 21364
rect 16100 21308 16110 21364
rect 17490 21308 17500 21364
rect 17556 21308 18060 21364
rect 18116 21308 20300 21364
rect 20356 21308 21028 21364
rect 24892 21308 27244 21364
rect 27300 21308 27692 21364
rect 27748 21308 27758 21364
rect 29474 21308 29484 21364
rect 29540 21308 30716 21364
rect 30772 21308 30782 21364
rect 35746 21308 35756 21364
rect 35812 21308 36764 21364
rect 36820 21308 36830 21364
rect 38444 21308 39452 21364
rect 39508 21308 39518 21364
rect 40562 21308 40572 21364
rect 40628 21308 47964 21364
rect 48020 21308 48030 21364
rect 49634 21308 49644 21364
rect 49700 21308 49738 21364
rect 49868 21308 51436 21364
rect 51492 21308 51502 21364
rect 51762 21308 51772 21364
rect 51828 21308 52892 21364
rect 52948 21308 56588 21364
rect 56644 21308 56654 21364
rect 20972 21252 21028 21308
rect 13570 21196 13580 21252
rect 13636 21196 20748 21252
rect 20804 21196 20814 21252
rect 20972 21196 23772 21252
rect 23828 21196 23838 21252
rect 33506 21196 33516 21252
rect 33572 21196 34188 21252
rect 34244 21196 34254 21252
rect 38210 21196 38220 21252
rect 38276 21196 38892 21252
rect 38948 21196 38958 21252
rect 46582 21196 46620 21252
rect 46676 21196 46686 21252
rect 47058 21196 47068 21252
rect 47124 21196 49756 21252
rect 49812 21196 49822 21252
rect 50978 21196 50988 21252
rect 51044 21196 53228 21252
rect 53284 21196 55468 21252
rect 55524 21196 55534 21252
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 12898 21084 12908 21140
rect 12964 21084 15148 21140
rect 15810 21084 15820 21140
rect 15876 21084 18396 21140
rect 18452 21084 22316 21140
rect 22372 21084 22382 21140
rect 38546 21084 38556 21140
rect 38612 21084 53340 21140
rect 53396 21084 53406 21140
rect 54002 21084 54012 21140
rect 54068 21084 54124 21140
rect 54180 21084 54190 21140
rect 15092 21028 15148 21084
rect 4386 20972 4396 21028
rect 4452 20972 5404 21028
rect 5460 20972 10332 21028
rect 10388 20972 13692 21028
rect 13748 20972 13758 21028
rect 15092 20972 15372 21028
rect 15428 20972 23100 21028
rect 23156 20972 23166 21028
rect 35410 20972 35420 21028
rect 35476 20972 35644 21028
rect 35700 20972 35710 21028
rect 35858 20972 35868 21028
rect 35924 20972 37660 21028
rect 37716 20972 37726 21028
rect 40002 20972 40012 21028
rect 40068 20972 40348 21028
rect 40404 20972 40414 21028
rect 41794 20972 41804 21028
rect 41860 20972 42252 21028
rect 42308 20972 42318 21028
rect 44034 20972 44044 21028
rect 44100 20972 44156 21028
rect 44212 20972 44222 21028
rect 45798 20972 45836 21028
rect 45892 20972 45902 21028
rect 46050 20972 46060 21028
rect 46116 20972 49756 21028
rect 49812 20972 49822 21028
rect 50754 20972 50764 21028
rect 50820 20972 51436 21028
rect 51492 20972 57708 21028
rect 57764 20972 57774 21028
rect 58258 20972 58268 21028
rect 58324 20972 58604 21028
rect 58660 20972 58670 21028
rect 12338 20860 12348 20916
rect 12404 20860 13244 20916
rect 13300 20860 13310 20916
rect 16482 20860 16492 20916
rect 16548 20860 17724 20916
rect 17780 20860 17790 20916
rect 18610 20860 18620 20916
rect 18676 20860 19292 20916
rect 19348 20860 19358 20916
rect 20626 20860 20636 20916
rect 20692 20860 22652 20916
rect 22708 20860 22718 20916
rect 25218 20860 25228 20916
rect 25284 20860 25340 20916
rect 25396 20860 25406 20916
rect 26450 20860 26460 20916
rect 26516 20860 28252 20916
rect 28308 20860 28318 20916
rect 32274 20860 32284 20916
rect 32340 20860 33404 20916
rect 33460 20860 33470 20916
rect 34402 20860 34412 20916
rect 34468 20860 36652 20916
rect 36708 20860 36718 20916
rect 39554 20860 39564 20916
rect 39620 20860 41132 20916
rect 41188 20860 42364 20916
rect 42420 20860 42430 20916
rect 43698 20860 43708 20916
rect 43764 20860 45388 20916
rect 45444 20860 45454 20916
rect 45602 20860 45612 20916
rect 45668 20860 46956 20916
rect 47012 20860 51100 20916
rect 51156 20860 51548 20916
rect 51604 20860 51614 20916
rect 52658 20860 52668 20916
rect 52724 20860 57820 20916
rect 57876 20860 57886 20916
rect 2034 20748 2044 20804
rect 2100 20748 6300 20804
rect 6356 20748 6366 20804
rect 6626 20748 6636 20804
rect 6692 20748 8988 20804
rect 9044 20748 9054 20804
rect 10546 20748 10556 20804
rect 10612 20748 14588 20804
rect 14644 20748 14654 20804
rect 15092 20748 27972 20804
rect 28130 20748 28140 20804
rect 28196 20748 30828 20804
rect 30884 20748 30894 20804
rect 38098 20748 38108 20804
rect 38164 20748 40908 20804
rect 40964 20748 40974 20804
rect 41234 20748 41244 20804
rect 41300 20748 41468 20804
rect 41524 20748 41534 20804
rect 42774 20748 42812 20804
rect 42868 20748 42878 20804
rect 43026 20748 43036 20804
rect 43092 20748 43708 20804
rect 43764 20748 43774 20804
rect 45266 20748 45276 20804
rect 45332 20748 46620 20804
rect 46676 20748 48412 20804
rect 48468 20748 51660 20804
rect 51716 20748 51726 20804
rect 51874 20748 51884 20804
rect 51940 20748 53900 20804
rect 53956 20748 54012 20804
rect 54068 20748 54078 20804
rect 55010 20748 55020 20804
rect 55076 20748 57372 20804
rect 57428 20748 57708 20804
rect 57764 20748 57774 20804
rect 15092 20692 15148 20748
rect 27916 20692 27972 20748
rect 1698 20636 1708 20692
rect 1764 20636 3052 20692
rect 3108 20636 3118 20692
rect 4610 20636 4620 20692
rect 4676 20636 14252 20692
rect 14308 20636 15148 20692
rect 19170 20636 19180 20692
rect 19236 20636 19516 20692
rect 19572 20636 21532 20692
rect 21588 20636 23324 20692
rect 23380 20636 23390 20692
rect 24658 20636 24668 20692
rect 24724 20636 25116 20692
rect 25172 20636 25182 20692
rect 27916 20636 29932 20692
rect 29988 20636 29998 20692
rect 31490 20636 31500 20692
rect 31556 20636 36652 20692
rect 36708 20636 36718 20692
rect 38322 20636 38332 20692
rect 38388 20636 38556 20692
rect 38612 20636 38622 20692
rect 39890 20636 39900 20692
rect 39956 20636 40460 20692
rect 40516 20636 41076 20692
rect 42690 20636 42700 20692
rect 42756 20636 43596 20692
rect 43652 20636 44268 20692
rect 44324 20636 44334 20692
rect 47366 20636 47404 20692
rect 47460 20636 47470 20692
rect 48290 20636 48300 20692
rect 48356 20636 55580 20692
rect 55636 20636 55646 20692
rect 39900 20580 39956 20636
rect 41020 20580 41076 20636
rect 3266 20524 3276 20580
rect 3332 20524 6300 20580
rect 6356 20524 6748 20580
rect 6804 20524 6814 20580
rect 7522 20524 7532 20580
rect 7588 20524 7980 20580
rect 8036 20524 8046 20580
rect 8530 20524 8540 20580
rect 8596 20524 12572 20580
rect 12628 20524 12638 20580
rect 14802 20524 14812 20580
rect 14868 20524 21644 20580
rect 21700 20524 21710 20580
rect 22838 20524 22876 20580
rect 22932 20524 22942 20580
rect 24892 20524 27468 20580
rect 27524 20524 27534 20580
rect 27682 20524 27692 20580
rect 27748 20524 29036 20580
rect 29092 20524 29102 20580
rect 30034 20524 30044 20580
rect 30100 20524 30380 20580
rect 30436 20524 31948 20580
rect 32004 20524 32014 20580
rect 32498 20524 32508 20580
rect 32564 20524 33628 20580
rect 33684 20524 36204 20580
rect 36260 20524 36270 20580
rect 36754 20524 36764 20580
rect 36820 20524 37436 20580
rect 37492 20524 38444 20580
rect 38500 20524 39956 20580
rect 40338 20524 40348 20580
rect 40404 20524 40796 20580
rect 40852 20524 40862 20580
rect 41020 20524 43932 20580
rect 43988 20524 43998 20580
rect 48598 20524 48636 20580
rect 48692 20524 48702 20580
rect 48850 20524 48860 20580
rect 48916 20524 49980 20580
rect 50036 20524 50046 20580
rect 50372 20524 52052 20580
rect 52210 20524 52220 20580
rect 52276 20524 53004 20580
rect 53060 20524 54572 20580
rect 54628 20524 54638 20580
rect 56354 20524 56364 20580
rect 56420 20524 57932 20580
rect 57988 20524 57998 20580
rect 3378 20412 3388 20468
rect 3444 20412 3612 20468
rect 3668 20412 3678 20468
rect 9090 20412 9100 20468
rect 9156 20412 11564 20468
rect 11620 20412 16716 20468
rect 16772 20412 18284 20468
rect 18340 20412 18508 20468
rect 18564 20412 18574 20468
rect 20710 20412 20748 20468
rect 20804 20412 20814 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 24892 20356 24948 20524
rect 50372 20468 50428 20524
rect 26002 20412 26012 20468
rect 26068 20412 26796 20468
rect 26852 20412 28140 20468
rect 28196 20412 28206 20468
rect 33170 20412 33180 20468
rect 33236 20412 33246 20468
rect 35298 20412 35308 20468
rect 35364 20412 35532 20468
rect 35588 20412 35756 20468
rect 35812 20412 35822 20468
rect 36866 20412 36876 20468
rect 36932 20412 41468 20468
rect 41524 20412 41534 20468
rect 42466 20412 42476 20468
rect 42532 20412 43036 20468
rect 43092 20412 43102 20468
rect 44268 20412 45612 20468
rect 45668 20412 45678 20468
rect 47618 20412 47628 20468
rect 47684 20412 48580 20468
rect 48738 20412 48748 20468
rect 48804 20412 49084 20468
rect 49140 20412 50428 20468
rect 51996 20468 52052 20524
rect 51996 20412 59052 20468
rect 59108 20412 59118 20468
rect 33180 20356 33236 20412
rect 44268 20356 44324 20412
rect 48524 20356 48580 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 3042 20300 3052 20356
rect 3108 20300 4172 20356
rect 4228 20300 4956 20356
rect 5012 20300 11676 20356
rect 11732 20300 11742 20356
rect 12226 20300 12236 20356
rect 12292 20300 12404 20356
rect 12786 20300 12796 20356
rect 12852 20300 18060 20356
rect 18116 20300 18126 20356
rect 20514 20300 20524 20356
rect 20580 20300 21756 20356
rect 21812 20300 21822 20356
rect 23874 20300 23884 20356
rect 23940 20300 24892 20356
rect 24948 20300 24958 20356
rect 25862 20300 25900 20356
rect 25956 20300 25966 20356
rect 33180 20300 33628 20356
rect 33684 20300 34860 20356
rect 34916 20300 34926 20356
rect 35186 20300 35196 20356
rect 35252 20300 35756 20356
rect 35812 20300 35822 20356
rect 37090 20300 37100 20356
rect 37156 20300 40348 20356
rect 40404 20300 40414 20356
rect 40674 20300 40684 20356
rect 40740 20300 44324 20356
rect 44594 20300 44604 20356
rect 44660 20300 46620 20356
rect 46676 20300 48300 20356
rect 48356 20300 48366 20356
rect 48524 20300 50316 20356
rect 50372 20300 50382 20356
rect 52322 20300 52332 20356
rect 52388 20300 54628 20356
rect 12348 20244 12404 20300
rect 2146 20188 2156 20244
rect 2212 20188 5404 20244
rect 5460 20188 6412 20244
rect 6468 20188 6478 20244
rect 7298 20188 7308 20244
rect 7364 20188 7980 20244
rect 8036 20188 8046 20244
rect 12348 20188 14700 20244
rect 14756 20188 14766 20244
rect 18162 20188 18172 20244
rect 18228 20188 19404 20244
rect 19460 20188 22316 20244
rect 22372 20188 22382 20244
rect 24406 20188 24444 20244
rect 24500 20188 24510 20244
rect 25778 20188 25788 20244
rect 25844 20188 26012 20244
rect 26068 20188 26078 20244
rect 28354 20188 28364 20244
rect 28420 20188 29092 20244
rect 31826 20188 31836 20244
rect 31892 20188 35364 20244
rect 39106 20188 39116 20244
rect 39172 20188 40124 20244
rect 40180 20188 40190 20244
rect 40786 20188 40796 20244
rect 40852 20188 41804 20244
rect 41860 20188 41870 20244
rect 42802 20188 42812 20244
rect 42868 20188 43484 20244
rect 43540 20188 45836 20244
rect 45892 20188 46284 20244
rect 46340 20188 46350 20244
rect 46722 20188 46732 20244
rect 46788 20188 46798 20244
rect 48626 20188 48636 20244
rect 48692 20188 51212 20244
rect 51268 20188 51278 20244
rect 51846 20188 51884 20244
rect 51940 20188 51950 20244
rect 53554 20188 53564 20244
rect 53620 20188 54124 20244
rect 54180 20188 54190 20244
rect 54338 20188 54348 20244
rect 54404 20188 54414 20244
rect 29036 20132 29092 20188
rect 35308 20132 35364 20188
rect 46732 20132 46788 20188
rect 54348 20132 54404 20188
rect 1922 20076 1932 20132
rect 1988 20076 2604 20132
rect 2660 20076 2670 20132
rect 4722 20076 4732 20132
rect 4788 20076 4956 20132
rect 5012 20076 7196 20132
rect 7252 20076 7262 20132
rect 15698 20076 15708 20132
rect 15764 20076 21868 20132
rect 21924 20076 21934 20132
rect 22642 20076 22652 20132
rect 22708 20076 23772 20132
rect 23828 20076 24668 20132
rect 24724 20076 26964 20132
rect 27122 20076 27132 20132
rect 27188 20076 27692 20132
rect 27748 20076 27758 20132
rect 29026 20076 29036 20132
rect 29092 20076 29102 20132
rect 29782 20076 29820 20132
rect 29876 20076 29886 20132
rect 35308 20076 43596 20132
rect 43652 20076 43662 20132
rect 43820 20076 44940 20132
rect 44996 20076 45006 20132
rect 46732 20076 47404 20132
rect 47460 20076 47470 20132
rect 49074 20076 49084 20132
rect 49140 20076 49420 20132
rect 49476 20076 49486 20132
rect 49746 20076 49756 20132
rect 49812 20076 51772 20132
rect 51828 20076 51838 20132
rect 53666 20076 53676 20132
rect 53732 20076 54404 20132
rect 54572 20132 54628 20300
rect 59200 20244 59800 20272
rect 56018 20188 56028 20244
rect 56084 20188 59800 20244
rect 59200 20160 59800 20188
rect 54572 20076 56476 20132
rect 56532 20076 56542 20132
rect 56690 20076 56700 20132
rect 56756 20076 57484 20132
rect 57540 20076 58044 20132
rect 58100 20076 58716 20132
rect 58772 20076 58782 20132
rect 26908 20020 26964 20076
rect 43820 20020 43876 20076
rect 3378 19964 3388 20020
rect 3444 19964 4508 20020
rect 4564 19964 4574 20020
rect 4946 19964 4956 20020
rect 5012 19964 7308 20020
rect 7364 19964 7374 20020
rect 8082 19964 8092 20020
rect 8148 19964 10444 20020
rect 10500 19964 10510 20020
rect 12674 19964 12684 20020
rect 12740 19964 14028 20020
rect 14084 19964 14094 20020
rect 19030 19964 19068 20020
rect 19124 19964 19134 20020
rect 19282 19964 19292 20020
rect 19348 19964 24332 20020
rect 24388 19964 24398 20020
rect 25554 19964 25564 20020
rect 25620 19964 26236 20020
rect 26292 19964 26302 20020
rect 26908 19964 28140 20020
rect 28196 19964 29708 20020
rect 29764 19964 31724 20020
rect 31780 19964 31790 20020
rect 34514 19964 34524 20020
rect 34580 19964 37548 20020
rect 37604 19964 37614 20020
rect 41010 19964 41020 20020
rect 41076 19964 42588 20020
rect 42644 19964 42654 20020
rect 42812 19964 43876 20020
rect 44230 19964 44268 20020
rect 44324 19964 48300 20020
rect 48356 19964 48366 20020
rect 48850 19964 48860 20020
rect 48916 19964 50204 20020
rect 50260 19964 50316 20020
rect 50372 19964 50382 20020
rect 50754 19964 50764 20020
rect 50820 19964 51660 20020
rect 51716 19964 51726 20020
rect 51874 19964 51884 20020
rect 51940 19964 52388 20020
rect 54338 19964 54348 20020
rect 54404 19964 55804 20020
rect 55860 19964 55870 20020
rect 42812 19908 42868 19964
rect 52332 19908 52388 19964
rect 5702 19852 5740 19908
rect 5796 19852 5806 19908
rect 6626 19852 6636 19908
rect 6692 19852 10892 19908
rect 10948 19852 13580 19908
rect 13636 19852 13646 19908
rect 13794 19852 13804 19908
rect 13860 19852 13916 19908
rect 13972 19852 13982 19908
rect 14690 19852 14700 19908
rect 14756 19852 15932 19908
rect 15988 19852 15998 19908
rect 16146 19852 16156 19908
rect 16212 19852 16716 19908
rect 16772 19852 16782 19908
rect 17938 19852 17948 19908
rect 18004 19852 21084 19908
rect 21140 19852 21980 19908
rect 22036 19852 24332 19908
rect 24388 19852 24398 19908
rect 28242 19852 28252 19908
rect 28308 19852 30156 19908
rect 30212 19852 31276 19908
rect 31332 19852 31342 19908
rect 36082 19852 36092 19908
rect 36148 19852 36876 19908
rect 36932 19852 36942 19908
rect 37958 19852 37996 19908
rect 38052 19852 38062 19908
rect 40226 19852 40236 19908
rect 40292 19852 40572 19908
rect 40628 19852 40638 19908
rect 42018 19852 42028 19908
rect 42084 19852 42868 19908
rect 46498 19852 46508 19908
rect 46564 19852 47180 19908
rect 47236 19852 52108 19908
rect 52164 19852 52174 19908
rect 52332 19852 53116 19908
rect 53172 19852 54460 19908
rect 54516 19852 54526 19908
rect 55234 19852 55244 19908
rect 55300 19852 55468 19908
rect 55524 19852 55534 19908
rect 2594 19740 2604 19796
rect 2660 19740 12460 19796
rect 12516 19740 14252 19796
rect 14308 19740 14318 19796
rect 15810 19740 15820 19796
rect 15876 19740 16604 19796
rect 16660 19740 16670 19796
rect 17154 19740 17164 19796
rect 17220 19740 22764 19796
rect 22820 19740 23548 19796
rect 23604 19740 23614 19796
rect 24546 19740 24556 19796
rect 24612 19740 25452 19796
rect 25508 19740 25518 19796
rect 32946 19740 32956 19796
rect 33012 19740 33852 19796
rect 33908 19740 34748 19796
rect 34804 19740 38668 19796
rect 43362 19740 43372 19796
rect 43428 19740 43484 19796
rect 43540 19740 43550 19796
rect 44034 19740 44044 19796
rect 44100 19740 44604 19796
rect 44660 19740 44670 19796
rect 49494 19740 49532 19796
rect 49588 19740 49598 19796
rect 50642 19740 50652 19796
rect 50708 19740 51548 19796
rect 51604 19740 51996 19796
rect 52052 19740 52062 19796
rect 38612 19684 38668 19740
rect 6066 19628 6076 19684
rect 6132 19628 10332 19684
rect 10388 19628 11116 19684
rect 11172 19628 11182 19684
rect 11330 19628 11340 19684
rect 11396 19628 19740 19684
rect 19796 19628 20860 19684
rect 20916 19628 20926 19684
rect 21858 19628 21868 19684
rect 21924 19628 23548 19684
rect 23604 19628 23614 19684
rect 23762 19628 23772 19684
rect 23828 19628 26460 19684
rect 26516 19628 31724 19684
rect 31780 19628 31790 19684
rect 38612 19628 42700 19684
rect 42756 19628 42924 19684
rect 42980 19628 44380 19684
rect 44436 19628 44446 19684
rect 45154 19628 45164 19684
rect 45220 19628 46172 19684
rect 46228 19628 51548 19684
rect 51604 19628 51614 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 45164 19572 45220 19628
rect 7532 19516 8988 19572
rect 9044 19516 9054 19572
rect 10098 19516 10108 19572
rect 10164 19516 10780 19572
rect 10836 19516 10846 19572
rect 13458 19516 13468 19572
rect 13524 19516 13916 19572
rect 13972 19516 13982 19572
rect 15362 19516 15372 19572
rect 15428 19516 15820 19572
rect 15876 19516 15886 19572
rect 19394 19516 19404 19572
rect 19460 19516 22428 19572
rect 22484 19516 22988 19572
rect 23044 19516 23054 19572
rect 24322 19516 24332 19572
rect 24388 19516 24556 19572
rect 24612 19516 27580 19572
rect 27636 19516 27646 19572
rect 40002 19516 40012 19572
rect 40068 19516 42812 19572
rect 42868 19516 44044 19572
rect 44100 19516 44110 19572
rect 44258 19516 44268 19572
rect 44324 19516 45220 19572
rect 47506 19516 47516 19572
rect 47572 19516 54908 19572
rect 54964 19516 54974 19572
rect 7532 19460 7588 19516
rect 3714 19404 3724 19460
rect 3780 19404 7588 19460
rect 7746 19404 7756 19460
rect 7812 19404 13356 19460
rect 13412 19404 13422 19460
rect 13570 19404 13580 19460
rect 13636 19404 14700 19460
rect 14756 19404 14766 19460
rect 15474 19404 15484 19460
rect 15540 19404 15932 19460
rect 15988 19404 15998 19460
rect 18498 19404 18508 19460
rect 18564 19404 21308 19460
rect 21364 19404 30044 19460
rect 30100 19404 30110 19460
rect 36418 19404 36428 19460
rect 36484 19404 38668 19460
rect 38724 19404 38734 19460
rect 41682 19404 41692 19460
rect 41748 19404 45612 19460
rect 45668 19404 45678 19460
rect 46162 19404 46172 19460
rect 46228 19404 47404 19460
rect 47460 19404 47852 19460
rect 47908 19404 47918 19460
rect 48290 19404 48300 19460
rect 48356 19404 49252 19460
rect 49634 19404 49644 19460
rect 49700 19404 53116 19460
rect 53172 19404 53182 19460
rect 53442 19404 53452 19460
rect 53508 19404 54012 19460
rect 54068 19404 54078 19460
rect 49196 19348 49252 19404
rect 2930 19292 2940 19348
rect 2996 19292 8092 19348
rect 8148 19292 8158 19348
rect 10294 19292 10332 19348
rect 10388 19292 10398 19348
rect 12450 19292 12460 19348
rect 12516 19292 13132 19348
rect 13188 19292 13916 19348
rect 13972 19292 19404 19348
rect 19460 19292 19470 19348
rect 19590 19292 19628 19348
rect 19684 19292 19694 19348
rect 23538 19292 23548 19348
rect 23604 19292 24780 19348
rect 24836 19292 26460 19348
rect 26516 19292 26572 19348
rect 26628 19292 26638 19348
rect 37202 19292 37212 19348
rect 37268 19292 37884 19348
rect 37940 19292 41468 19348
rect 41524 19292 41534 19348
rect 43586 19292 43596 19348
rect 43652 19292 44156 19348
rect 44212 19292 45388 19348
rect 45444 19292 45454 19348
rect 45910 19292 45948 19348
rect 46004 19292 46014 19348
rect 46610 19292 46620 19348
rect 46676 19292 46956 19348
rect 47012 19292 47022 19348
rect 48934 19292 48972 19348
rect 49028 19292 49038 19348
rect 49196 19292 54012 19348
rect 54068 19292 54078 19348
rect 55122 19292 55132 19348
rect 55188 19292 56812 19348
rect 56868 19292 56878 19348
rect 2370 19180 2380 19236
rect 2436 19180 3612 19236
rect 3668 19180 3678 19236
rect 3938 19180 3948 19236
rect 4004 19180 6524 19236
rect 6580 19180 6590 19236
rect 8418 19180 8428 19236
rect 8484 19180 8652 19236
rect 8708 19180 8718 19236
rect 8978 19180 8988 19236
rect 9044 19180 10444 19236
rect 10500 19180 10892 19236
rect 10948 19180 12684 19236
rect 12740 19180 12750 19236
rect 12898 19180 12908 19236
rect 12964 19180 13692 19236
rect 13748 19180 13804 19236
rect 13860 19180 13870 19236
rect 14914 19180 14924 19236
rect 14980 19180 15260 19236
rect 15316 19180 17612 19236
rect 17668 19180 17678 19236
rect 19404 19124 19460 19292
rect 45388 19236 45444 19292
rect 23314 19180 23324 19236
rect 23380 19180 24332 19236
rect 24388 19180 26348 19236
rect 26404 19180 26414 19236
rect 32946 19180 32956 19236
rect 33012 19180 34748 19236
rect 34804 19180 40012 19236
rect 40068 19180 40078 19236
rect 42802 19180 42812 19236
rect 42868 19180 43820 19236
rect 43876 19180 43886 19236
rect 44930 19180 44940 19236
rect 44996 19180 45164 19236
rect 45220 19180 45230 19236
rect 45388 19180 47404 19236
rect 47460 19180 47470 19236
rect 48738 19180 48748 19236
rect 48804 19180 49868 19236
rect 49924 19180 49934 19236
rect 50530 19180 50540 19236
rect 50596 19180 50988 19236
rect 51044 19180 51054 19236
rect 51426 19180 51436 19236
rect 51492 19180 53228 19236
rect 53284 19180 53452 19236
rect 53508 19180 53788 19236
rect 53844 19180 53854 19236
rect 56578 19180 56588 19236
rect 56644 19180 57316 19236
rect 57260 19124 57316 19180
rect 3266 19068 3276 19124
rect 3332 19068 4060 19124
rect 4116 19068 4956 19124
rect 5012 19068 10220 19124
rect 10276 19068 14140 19124
rect 14196 19068 15148 19124
rect 15204 19068 15260 19124
rect 15316 19068 16044 19124
rect 16100 19068 16110 19124
rect 19404 19068 19628 19124
rect 19684 19068 19694 19124
rect 27682 19068 27692 19124
rect 27748 19068 29932 19124
rect 29988 19068 30268 19124
rect 30324 19068 30334 19124
rect 34850 19068 34860 19124
rect 34916 19068 35868 19124
rect 35924 19068 35934 19124
rect 37874 19068 37884 19124
rect 37940 19068 39228 19124
rect 39284 19068 39294 19124
rect 39442 19068 39452 19124
rect 39508 19068 39676 19124
rect 39732 19068 40348 19124
rect 40404 19068 40414 19124
rect 41906 19068 41916 19124
rect 41972 19068 42924 19124
rect 42980 19068 45836 19124
rect 45892 19068 46620 19124
rect 46676 19068 46686 19124
rect 47618 19068 47628 19124
rect 47684 19068 47852 19124
rect 47908 19068 49532 19124
rect 49588 19068 49598 19124
rect 50194 19068 50204 19124
rect 50260 19068 50652 19124
rect 50708 19068 50718 19124
rect 51538 19068 51548 19124
rect 51604 19068 52220 19124
rect 52276 19068 52286 19124
rect 55794 19068 55804 19124
rect 55860 19068 56924 19124
rect 56980 19068 56990 19124
rect 57222 19068 57260 19124
rect 57316 19068 57326 19124
rect 3714 18956 3724 19012
rect 3780 18956 4620 19012
rect 4676 18956 5964 19012
rect 6020 18956 6030 19012
rect 8082 18956 8092 19012
rect 8148 18956 10780 19012
rect 10836 18956 10846 19012
rect 11778 18956 11788 19012
rect 11844 18956 13972 19012
rect 14242 18956 14252 19012
rect 14308 18956 16604 19012
rect 16660 18956 16670 19012
rect 17154 18956 17164 19012
rect 17220 18956 17948 19012
rect 18004 18956 18014 19012
rect 18162 18956 18172 19012
rect 18228 18956 19852 19012
rect 19908 18956 19918 19012
rect 21746 18956 21756 19012
rect 21812 18956 22876 19012
rect 22932 18956 23100 19012
rect 23156 18956 23166 19012
rect 24182 18956 24220 19012
rect 24276 18956 24286 19012
rect 26422 18956 26460 19012
rect 26516 18956 26526 19012
rect 26786 18956 26796 19012
rect 26852 18956 27132 19012
rect 27188 18956 27198 19012
rect 32498 18956 32508 19012
rect 32564 18956 35084 19012
rect 35140 18956 36092 19012
rect 36148 18956 36428 19012
rect 36484 18956 36494 19012
rect 37090 18956 37100 19012
rect 37156 18956 37772 19012
rect 37828 18956 37838 19012
rect 39106 18956 39116 19012
rect 39172 18956 39900 19012
rect 39956 18956 42532 19012
rect 43138 18956 43148 19012
rect 43204 18956 44716 19012
rect 44772 18956 46172 19012
rect 46228 18956 46238 19012
rect 46946 18956 46956 19012
rect 47012 18956 51996 19012
rect 52052 18956 52062 19012
rect 54674 18956 54684 19012
rect 54740 18956 55132 19012
rect 55188 18956 55198 19012
rect 55430 18956 55468 19012
rect 55524 18956 55534 19012
rect 56242 18956 56252 19012
rect 56308 18956 56476 19012
rect 56532 18956 59164 19012
rect 59220 18956 59230 19012
rect 3602 18844 3612 18900
rect 3668 18844 12460 18900
rect 12516 18844 12526 18900
rect 13916 18788 13972 18956
rect 16034 18844 16044 18900
rect 16100 18844 18172 18900
rect 18228 18844 18238 18900
rect 18498 18844 18508 18900
rect 18564 18844 18620 18900
rect 18676 18844 18686 18900
rect 30258 18844 30268 18900
rect 30324 18844 31276 18900
rect 31332 18844 31342 18900
rect 39666 18844 39676 18900
rect 39732 18844 40236 18900
rect 40292 18844 40302 18900
rect 40674 18844 40684 18900
rect 40740 18844 40796 18900
rect 40852 18844 40862 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 42476 18788 42532 18956
rect 46386 18844 46396 18900
rect 46452 18844 47516 18900
rect 47572 18844 50204 18900
rect 50260 18844 50270 18900
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 51324 18788 51380 18956
rect 52434 18844 52444 18900
rect 52500 18844 58828 18900
rect 58884 18844 58894 18900
rect 2818 18732 2828 18788
rect 2884 18732 8988 18788
rect 9044 18732 9996 18788
rect 10052 18732 10220 18788
rect 10276 18732 10286 18788
rect 11666 18732 11676 18788
rect 11732 18732 12124 18788
rect 12180 18732 12190 18788
rect 12310 18732 12348 18788
rect 12404 18732 12414 18788
rect 13906 18732 13916 18788
rect 13972 18732 18172 18788
rect 18228 18732 18238 18788
rect 23986 18732 23996 18788
rect 24052 18732 24892 18788
rect 24948 18732 24958 18788
rect 25890 18732 25900 18788
rect 25956 18732 27020 18788
rect 27076 18732 27086 18788
rect 29698 18732 29708 18788
rect 29764 18732 30156 18788
rect 30212 18732 30604 18788
rect 30660 18732 30670 18788
rect 31826 18732 31836 18788
rect 31892 18732 32508 18788
rect 32564 18732 32574 18788
rect 36642 18732 36652 18788
rect 36708 18732 37100 18788
rect 37156 18732 37548 18788
rect 37604 18732 37614 18788
rect 42466 18732 42476 18788
rect 42532 18732 45892 18788
rect 48626 18732 48636 18788
rect 48692 18732 49308 18788
rect 49364 18732 49374 18788
rect 49746 18732 49756 18788
rect 49812 18732 50316 18788
rect 50372 18732 50382 18788
rect 51314 18732 51324 18788
rect 51380 18732 51390 18788
rect 52098 18732 52108 18788
rect 52164 18732 52780 18788
rect 52836 18732 52892 18788
rect 52948 18732 52958 18788
rect 54450 18732 54460 18788
rect 54516 18732 54908 18788
rect 54964 18732 54974 18788
rect 1922 18620 1932 18676
rect 1988 18620 8428 18676
rect 8484 18620 8494 18676
rect 9090 18620 9100 18676
rect 9156 18620 11788 18676
rect 11844 18620 12460 18676
rect 12516 18620 13020 18676
rect 13076 18620 13086 18676
rect 15670 18620 15708 18676
rect 15764 18620 15774 18676
rect 15922 18620 15932 18676
rect 15988 18620 17500 18676
rect 17556 18620 17566 18676
rect 17938 18620 17948 18676
rect 18004 18620 18284 18676
rect 18340 18620 21980 18676
rect 22036 18620 22046 18676
rect 23314 18620 23324 18676
rect 23380 18620 23436 18676
rect 23492 18620 23502 18676
rect 26198 18620 26236 18676
rect 26292 18620 26302 18676
rect 28354 18620 28364 18676
rect 28420 18620 31276 18676
rect 31332 18620 31342 18676
rect 31490 18620 31500 18676
rect 31556 18620 32620 18676
rect 32676 18620 32686 18676
rect 36194 18620 36204 18676
rect 36260 18620 38780 18676
rect 38836 18620 41580 18676
rect 41636 18620 41646 18676
rect 43474 18620 43484 18676
rect 43540 18620 43596 18676
rect 43652 18620 43662 18676
rect 28924 18564 28980 18620
rect 5292 18508 5516 18564
rect 5572 18508 5582 18564
rect 6178 18508 6188 18564
rect 6244 18508 6636 18564
rect 6692 18508 6702 18564
rect 7858 18508 7868 18564
rect 7924 18508 8764 18564
rect 8820 18508 8830 18564
rect 10546 18508 10556 18564
rect 10612 18508 11564 18564
rect 11620 18508 11630 18564
rect 12114 18508 12124 18564
rect 12180 18508 15372 18564
rect 15428 18508 15438 18564
rect 15586 18508 15596 18564
rect 15652 18508 15820 18564
rect 15876 18508 15886 18564
rect 16594 18508 16604 18564
rect 16660 18508 20412 18564
rect 20468 18508 20478 18564
rect 20636 18508 24220 18564
rect 24276 18508 24286 18564
rect 28914 18508 28924 18564
rect 28980 18508 28990 18564
rect 31154 18508 31164 18564
rect 31220 18508 32172 18564
rect 32228 18508 32238 18564
rect 35970 18508 35980 18564
rect 36036 18508 37324 18564
rect 37380 18508 37390 18564
rect 37538 18508 37548 18564
rect 37604 18508 38668 18564
rect 39078 18508 39116 18564
rect 39172 18508 39182 18564
rect 40562 18508 40572 18564
rect 40628 18508 42588 18564
rect 42644 18508 42654 18564
rect 44258 18508 44268 18564
rect 44324 18508 45668 18564
rect 5292 18452 5348 18508
rect 20636 18452 20692 18508
rect 38612 18452 38668 18508
rect 45612 18452 45668 18508
rect 45836 18452 45892 18732
rect 46050 18620 46060 18676
rect 46116 18620 46956 18676
rect 47012 18620 54796 18676
rect 54852 18620 54862 18676
rect 56438 18620 56476 18676
rect 56532 18620 56542 18676
rect 57026 18620 57036 18676
rect 57092 18620 57820 18676
rect 57876 18620 57886 18676
rect 47394 18508 47404 18564
rect 47460 18508 50428 18564
rect 50866 18508 50876 18564
rect 50932 18508 51324 18564
rect 51380 18508 51390 18564
rect 51874 18508 51884 18564
rect 51940 18508 52444 18564
rect 52500 18508 53676 18564
rect 53732 18508 54012 18564
rect 54068 18508 54078 18564
rect 54898 18508 54908 18564
rect 54964 18508 55804 18564
rect 55860 18508 55870 18564
rect 56690 18508 56700 18564
rect 56756 18508 57708 18564
rect 57764 18508 57774 18564
rect 50372 18452 50428 18508
rect 3490 18396 3500 18452
rect 3556 18396 3724 18452
rect 3780 18396 3790 18452
rect 3938 18396 3948 18452
rect 4004 18396 4620 18452
rect 4676 18396 4686 18452
rect 4844 18396 5348 18452
rect 5404 18396 7532 18452
rect 7588 18396 8540 18452
rect 8596 18396 8606 18452
rect 9090 18396 9100 18452
rect 9156 18396 11340 18452
rect 11396 18396 11406 18452
rect 12674 18396 12684 18452
rect 12740 18396 16716 18452
rect 16772 18396 16782 18452
rect 16930 18396 16940 18452
rect 16996 18396 17164 18452
rect 17220 18396 17230 18452
rect 18274 18396 18284 18452
rect 18340 18396 18956 18452
rect 19012 18396 19022 18452
rect 19170 18396 19180 18452
rect 19236 18396 19404 18452
rect 19460 18396 19470 18452
rect 19618 18396 19628 18452
rect 19684 18396 20692 18452
rect 21970 18396 21980 18452
rect 22036 18396 23772 18452
rect 23828 18396 23838 18452
rect 28354 18396 28364 18452
rect 28420 18396 28700 18452
rect 28756 18396 29596 18452
rect 29652 18396 29662 18452
rect 34290 18396 34300 18452
rect 34356 18396 35532 18452
rect 35588 18396 35598 18452
rect 38612 18396 40684 18452
rect 40740 18396 40750 18452
rect 42242 18396 42252 18452
rect 42308 18396 43036 18452
rect 43092 18396 43102 18452
rect 45602 18396 45612 18452
rect 45668 18396 45678 18452
rect 45836 18396 47180 18452
rect 47236 18396 48300 18452
rect 48356 18396 48366 18452
rect 49494 18396 49532 18452
rect 49588 18396 49598 18452
rect 50372 18396 52108 18452
rect 52164 18396 52174 18452
rect 53218 18396 53228 18452
rect 53284 18396 54236 18452
rect 54292 18396 54302 18452
rect 54674 18396 54684 18452
rect 54740 18396 55916 18452
rect 55972 18396 55982 18452
rect 4844 18340 4900 18396
rect 3042 18284 3052 18340
rect 3108 18284 4284 18340
rect 4340 18284 4900 18340
rect 5404 18228 5460 18396
rect 8642 18284 8652 18340
rect 8708 18284 9772 18340
rect 9828 18284 9838 18340
rect 9996 18284 11452 18340
rect 11508 18284 12460 18340
rect 12516 18284 12526 18340
rect 13346 18284 13356 18340
rect 13412 18284 19292 18340
rect 19348 18284 19358 18340
rect 20076 18284 21084 18340
rect 21140 18284 21150 18340
rect 21830 18284 21868 18340
rect 21924 18284 21934 18340
rect 22978 18284 22988 18340
rect 23044 18284 23436 18340
rect 23492 18284 23502 18340
rect 25638 18284 25676 18340
rect 25732 18284 28028 18340
rect 28084 18284 28094 18340
rect 34402 18284 34412 18340
rect 34468 18284 36876 18340
rect 36932 18284 37996 18340
rect 38052 18284 38062 18340
rect 40898 18284 40908 18340
rect 40964 18284 43036 18340
rect 43092 18284 47628 18340
rect 47684 18284 47694 18340
rect 49410 18284 49420 18340
rect 49476 18284 49980 18340
rect 50036 18284 50046 18340
rect 50754 18284 50764 18340
rect 50820 18284 51100 18340
rect 51156 18284 51166 18340
rect 51762 18284 51772 18340
rect 51828 18284 53340 18340
rect 53396 18284 53788 18340
rect 53844 18284 53854 18340
rect 9996 18228 10052 18284
rect 20076 18228 20132 18284
rect 1810 18172 1820 18228
rect 1876 18172 5460 18228
rect 5516 18172 10052 18228
rect 10770 18172 10780 18228
rect 10836 18172 13244 18228
rect 13300 18172 13310 18228
rect 13458 18172 13468 18228
rect 13524 18172 13580 18228
rect 13636 18172 13646 18228
rect 14690 18172 14700 18228
rect 14756 18172 15708 18228
rect 15764 18172 15774 18228
rect 17042 18172 17052 18228
rect 17108 18172 20132 18228
rect 20738 18172 20748 18228
rect 20804 18172 21532 18228
rect 21588 18172 22092 18228
rect 22148 18172 22158 18228
rect 23538 18172 23548 18228
rect 23604 18172 24444 18228
rect 24500 18172 24510 18228
rect 32722 18172 32732 18228
rect 32788 18172 33740 18228
rect 33796 18172 33806 18228
rect 34290 18172 34300 18228
rect 34356 18172 34748 18228
rect 34804 18172 36876 18228
rect 36932 18172 36942 18228
rect 37090 18172 37100 18228
rect 37156 18172 37194 18228
rect 37650 18172 37660 18228
rect 37716 18172 38108 18228
rect 38164 18172 38174 18228
rect 41906 18172 41916 18228
rect 41972 18172 42252 18228
rect 42308 18172 42318 18228
rect 43250 18172 43260 18228
rect 43316 18172 44156 18228
rect 44212 18172 44222 18228
rect 47954 18172 47964 18228
rect 48020 18172 48412 18228
rect 48468 18172 48478 18228
rect 48626 18172 48636 18228
rect 48692 18172 52220 18228
rect 52276 18172 53564 18228
rect 53620 18172 53630 18228
rect 57474 18172 57484 18228
rect 57540 18172 58716 18228
rect 58772 18172 58782 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 5516 18004 5572 18172
rect 48412 18116 48468 18172
rect 7186 18060 7196 18116
rect 7252 18060 7532 18116
rect 7588 18060 8204 18116
rect 8260 18060 8270 18116
rect 9202 18060 9212 18116
rect 9268 18060 16828 18116
rect 16884 18060 18060 18116
rect 18116 18060 18126 18116
rect 18834 18060 18844 18116
rect 18900 18060 19068 18116
rect 19124 18060 19134 18116
rect 21858 18060 21868 18116
rect 21924 18060 28364 18116
rect 28420 18060 28430 18116
rect 36978 18060 36988 18116
rect 37044 18060 41804 18116
rect 41860 18060 44604 18116
rect 44660 18060 44940 18116
rect 44996 18060 45006 18116
rect 48412 18060 55580 18116
rect 55636 18060 55646 18116
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 5058 17948 5068 18004
rect 5124 17948 5516 18004
rect 5572 17948 5582 18004
rect 6626 17948 6636 18004
rect 6692 17948 9044 18004
rect 9538 17948 9548 18004
rect 9604 17948 11452 18004
rect 11508 17948 11518 18004
rect 11666 17948 11676 18004
rect 11732 17948 11770 18004
rect 13346 17948 13356 18004
rect 13412 17948 15372 18004
rect 15428 17948 15438 18004
rect 19170 17948 19180 18004
rect 19236 17948 25340 18004
rect 25396 17948 26012 18004
rect 26068 17948 26078 18004
rect 38612 17948 43820 18004
rect 43876 17948 44156 18004
rect 44212 17948 44222 18004
rect 44370 17948 44380 18004
rect 44436 17948 45164 18004
rect 45220 17948 45230 18004
rect 46162 17948 46172 18004
rect 46228 17948 49196 18004
rect 49252 17948 49262 18004
rect 50082 17948 50092 18004
rect 50148 17948 51884 18004
rect 51940 17948 51950 18004
rect 52098 17948 52108 18004
rect 52164 17948 52444 18004
rect 52500 17948 52510 18004
rect 52658 17948 52668 18004
rect 52724 17948 56252 18004
rect 56308 17948 56318 18004
rect 2258 17836 2268 17892
rect 2324 17836 8652 17892
rect 8708 17836 8718 17892
rect 1586 17724 1596 17780
rect 1652 17724 3052 17780
rect 3108 17724 3118 17780
rect 4050 17724 4060 17780
rect 4116 17724 8204 17780
rect 8260 17724 8270 17780
rect 8988 17668 9044 17948
rect 38612 17892 38668 17948
rect 9762 17836 9772 17892
rect 9828 17836 14924 17892
rect 14980 17836 14990 17892
rect 15698 17836 15708 17892
rect 15764 17836 16380 17892
rect 16436 17836 16446 17892
rect 17042 17836 17052 17892
rect 17108 17836 17164 17892
rect 17220 17836 17230 17892
rect 18834 17836 18844 17892
rect 18900 17836 19516 17892
rect 19572 17836 19740 17892
rect 19796 17836 19806 17892
rect 22754 17836 22764 17892
rect 22820 17836 23324 17892
rect 23380 17836 23390 17892
rect 23874 17836 23884 17892
rect 23940 17836 27244 17892
rect 27300 17836 28476 17892
rect 28532 17836 28542 17892
rect 34178 17836 34188 17892
rect 34244 17836 34636 17892
rect 34692 17836 38668 17892
rect 40310 17836 40348 17892
rect 40404 17836 40414 17892
rect 44034 17836 44044 17892
rect 44100 17836 45500 17892
rect 45556 17836 53564 17892
rect 53620 17836 53630 17892
rect 54114 17836 54124 17892
rect 54180 17836 54796 17892
rect 54852 17836 54862 17892
rect 9314 17724 9324 17780
rect 9380 17724 9660 17780
rect 9716 17724 9726 17780
rect 12450 17724 12460 17780
rect 12516 17724 13468 17780
rect 13524 17724 13916 17780
rect 13972 17724 13982 17780
rect 14140 17724 15428 17780
rect 16258 17724 16268 17780
rect 16324 17724 20412 17780
rect 20468 17724 21756 17780
rect 21812 17724 22652 17780
rect 22708 17724 22718 17780
rect 23426 17724 23436 17780
rect 23492 17724 23660 17780
rect 23716 17724 23726 17780
rect 28242 17724 28252 17780
rect 28308 17724 28588 17780
rect 28644 17724 29484 17780
rect 29540 17724 29550 17780
rect 33058 17724 33068 17780
rect 33124 17724 33404 17780
rect 33460 17724 33470 17780
rect 33730 17724 33740 17780
rect 33796 17724 33964 17780
rect 34020 17724 34030 17780
rect 36418 17724 36428 17780
rect 36484 17724 36876 17780
rect 36932 17724 36942 17780
rect 37398 17724 37436 17780
rect 37492 17724 37502 17780
rect 40786 17724 40796 17780
rect 40852 17724 41804 17780
rect 41860 17724 43596 17780
rect 43652 17724 43662 17780
rect 47142 17724 47180 17780
rect 47236 17724 47246 17780
rect 47730 17724 47740 17780
rect 47796 17724 48748 17780
rect 48804 17724 48814 17780
rect 49634 17724 49644 17780
rect 49700 17724 52108 17780
rect 52164 17724 52174 17780
rect 52322 17724 52332 17780
rect 52388 17724 52426 17780
rect 52994 17724 53004 17780
rect 53060 17724 53228 17780
rect 53284 17724 53452 17780
rect 53508 17724 53518 17780
rect 4134 17612 4172 17668
rect 4228 17612 4238 17668
rect 5058 17612 5068 17668
rect 5124 17612 6972 17668
rect 7028 17612 7038 17668
rect 7634 17612 7644 17668
rect 7700 17612 8316 17668
rect 8372 17612 8382 17668
rect 8988 17612 12908 17668
rect 12964 17612 12974 17668
rect 13458 17612 13468 17668
rect 13524 17612 13804 17668
rect 13860 17612 13870 17668
rect 14140 17556 14196 17724
rect 14354 17612 14364 17668
rect 14420 17612 15148 17668
rect 15204 17612 15214 17668
rect 5618 17500 5628 17556
rect 5684 17500 7084 17556
rect 7140 17500 7150 17556
rect 7858 17500 7868 17556
rect 7924 17500 8092 17556
rect 8148 17500 8540 17556
rect 8596 17500 8606 17556
rect 9650 17500 9660 17556
rect 9716 17500 14196 17556
rect 15372 17556 15428 17724
rect 17714 17612 17724 17668
rect 17780 17612 19628 17668
rect 19684 17612 19694 17668
rect 23314 17612 23324 17668
rect 23380 17612 25116 17668
rect 25172 17612 25182 17668
rect 26338 17612 26348 17668
rect 26404 17612 26684 17668
rect 26740 17612 26750 17668
rect 27346 17612 27356 17668
rect 27412 17612 29260 17668
rect 29316 17612 29820 17668
rect 29876 17612 29886 17668
rect 41458 17612 41468 17668
rect 41524 17612 41916 17668
rect 41972 17612 41982 17668
rect 43362 17612 43372 17668
rect 43428 17612 44716 17668
rect 44772 17612 45836 17668
rect 45892 17612 46844 17668
rect 46900 17612 46910 17668
rect 48290 17612 48300 17668
rect 48356 17612 49644 17668
rect 49700 17612 49710 17668
rect 49858 17612 49868 17668
rect 49924 17612 50316 17668
rect 50372 17612 57372 17668
rect 57428 17612 57438 17668
rect 15372 17500 18396 17556
rect 18452 17500 19180 17556
rect 19236 17500 19246 17556
rect 21410 17500 21420 17556
rect 21476 17500 23212 17556
rect 23268 17500 23278 17556
rect 24994 17500 25004 17556
rect 25060 17500 25788 17556
rect 25844 17500 26236 17556
rect 26292 17500 26302 17556
rect 32050 17500 32060 17556
rect 32116 17500 33852 17556
rect 33908 17500 33918 17556
rect 34962 17500 34972 17556
rect 35028 17500 37436 17556
rect 37492 17500 37502 17556
rect 41010 17500 41020 17556
rect 41076 17500 42140 17556
rect 42196 17500 42206 17556
rect 43372 17444 43428 17612
rect 44034 17500 44044 17556
rect 44100 17500 46172 17556
rect 46228 17500 46844 17556
rect 46900 17500 46910 17556
rect 48402 17500 48412 17556
rect 48468 17500 49980 17556
rect 50036 17500 54684 17556
rect 54740 17500 54750 17556
rect 55682 17500 55692 17556
rect 55748 17500 56476 17556
rect 56532 17500 56542 17556
rect 4610 17388 4620 17444
rect 4676 17388 4844 17444
rect 4900 17388 5964 17444
rect 6020 17388 6030 17444
rect 6402 17388 6412 17444
rect 6468 17388 10164 17444
rect 10322 17388 10332 17444
rect 10388 17388 11004 17444
rect 11060 17388 11070 17444
rect 13794 17388 13804 17444
rect 13860 17388 20860 17444
rect 20916 17388 22540 17444
rect 22596 17388 22606 17444
rect 23286 17388 23324 17444
rect 23380 17388 23390 17444
rect 25106 17388 25116 17444
rect 25172 17388 27916 17444
rect 27972 17388 27982 17444
rect 28914 17388 28924 17444
rect 28980 17388 29484 17444
rect 29540 17388 30492 17444
rect 30548 17388 30558 17444
rect 32722 17388 32732 17444
rect 32788 17388 33180 17444
rect 33236 17388 33246 17444
rect 35410 17388 35420 17444
rect 35476 17388 35644 17444
rect 35700 17388 35710 17444
rect 38322 17388 38332 17444
rect 38388 17388 43428 17444
rect 44192 17388 44268 17444
rect 44324 17388 44940 17444
rect 44996 17388 45006 17444
rect 45266 17388 45276 17444
rect 45332 17388 45500 17444
rect 45556 17388 45566 17444
rect 47954 17388 47964 17444
rect 48020 17388 48030 17444
rect 49298 17388 49308 17444
rect 49364 17388 50428 17444
rect 50484 17388 50876 17444
rect 50932 17388 50942 17444
rect 54562 17388 54572 17444
rect 54628 17388 54638 17444
rect 54870 17388 54908 17444
rect 54964 17388 54974 17444
rect 55570 17388 55580 17444
rect 55636 17388 56252 17444
rect 56308 17388 56318 17444
rect 57250 17388 57260 17444
rect 57316 17388 57708 17444
rect 57764 17388 57774 17444
rect 10108 17332 10164 17388
rect 47964 17332 48020 17388
rect 54572 17332 54628 17388
rect 3332 17276 9884 17332
rect 9940 17276 9950 17332
rect 10108 17276 14532 17332
rect 17378 17276 17388 17332
rect 17444 17276 18956 17332
rect 19012 17276 19022 17332
rect 20626 17276 20636 17332
rect 20692 17276 21756 17332
rect 21812 17276 21822 17332
rect 27010 17276 27020 17332
rect 27076 17276 28252 17332
rect 28308 17276 28318 17332
rect 31042 17276 31052 17332
rect 31108 17276 31612 17332
rect 31668 17276 31678 17332
rect 32162 17276 32172 17332
rect 32228 17276 33068 17332
rect 33124 17276 33134 17332
rect 36082 17276 36092 17332
rect 36148 17276 41580 17332
rect 41636 17276 41646 17332
rect 43810 17276 43820 17332
rect 43876 17276 46396 17332
rect 46452 17276 48020 17332
rect 49074 17276 49084 17332
rect 49140 17276 50204 17332
rect 50260 17276 50270 17332
rect 53890 17276 53900 17332
rect 53956 17276 54628 17332
rect 3332 17220 3388 17276
rect 9884 17220 9940 17276
rect 3042 17164 3052 17220
rect 3108 17164 3388 17220
rect 3490 17164 3500 17220
rect 3556 17164 4284 17220
rect 4340 17164 4956 17220
rect 5012 17164 5022 17220
rect 5180 17164 6636 17220
rect 6692 17164 6702 17220
rect 7298 17164 7308 17220
rect 7364 17164 8316 17220
rect 8372 17164 8382 17220
rect 9884 17164 12964 17220
rect 5180 16996 5236 17164
rect 6402 17052 6412 17108
rect 6468 17052 7532 17108
rect 7588 17052 7598 17108
rect 8316 17052 10108 17108
rect 10164 17052 10332 17108
rect 10388 17052 10892 17108
rect 10948 17052 10958 17108
rect 11862 17052 11900 17108
rect 11956 17052 11966 17108
rect 12236 17052 12684 17108
rect 12740 17052 12750 17108
rect 8316 16996 8372 17052
rect 12236 16996 12292 17052
rect 12908 16996 12964 17164
rect 14476 17108 14532 17276
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 36876 17220 36932 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 21298 17164 21308 17220
rect 21364 17164 21644 17220
rect 21700 17164 21710 17220
rect 24668 17164 30380 17220
rect 30436 17164 31724 17220
rect 31780 17164 32284 17220
rect 32340 17164 32350 17220
rect 36866 17164 36876 17220
rect 36932 17164 36942 17220
rect 43362 17164 43372 17220
rect 43428 17164 47068 17220
rect 47124 17164 47740 17220
rect 47796 17164 47806 17220
rect 54562 17164 54572 17220
rect 54628 17164 55356 17220
rect 55412 17164 55422 17220
rect 24668 17108 24724 17164
rect 14466 17052 14476 17108
rect 14532 17052 14812 17108
rect 14868 17052 14878 17108
rect 16930 17052 16940 17108
rect 16996 17052 17500 17108
rect 17556 17052 18172 17108
rect 18228 17052 18844 17108
rect 18900 17052 18910 17108
rect 19282 17052 19292 17108
rect 19348 17052 24724 17108
rect 25554 17052 25564 17108
rect 25620 17052 26348 17108
rect 26404 17052 26414 17108
rect 31266 17052 31276 17108
rect 31332 17052 32172 17108
rect 32228 17052 32238 17108
rect 33954 17052 33964 17108
rect 34020 17052 35532 17108
rect 35588 17052 35868 17108
rect 35924 17052 35980 17108
rect 36036 17052 36046 17108
rect 36978 17052 36988 17108
rect 37044 17052 37548 17108
rect 37604 17052 37614 17108
rect 40338 17052 40348 17108
rect 40404 17052 41804 17108
rect 41860 17052 41916 17108
rect 41972 17052 41982 17108
rect 43026 17052 43036 17108
rect 43092 17052 47964 17108
rect 48020 17052 48030 17108
rect 49074 17052 49084 17108
rect 49140 17052 49980 17108
rect 50036 17052 51772 17108
rect 51828 17052 51838 17108
rect 53526 17052 53564 17108
rect 53620 17052 53630 17108
rect 54422 17052 54460 17108
rect 54516 17052 54526 17108
rect 3266 16940 3276 16996
rect 3332 16940 5236 16996
rect 5394 16940 5404 16996
rect 5460 16940 5740 16996
rect 5796 16940 5806 16996
rect 6850 16940 6860 16996
rect 6916 16940 7308 16996
rect 7364 16940 7374 16996
rect 8306 16940 8316 16996
rect 8372 16940 8382 16996
rect 10994 16940 11004 16996
rect 11060 16940 12236 16996
rect 12292 16940 12302 16996
rect 12908 16940 15484 16996
rect 15540 16940 17724 16996
rect 17780 16940 18060 16996
rect 18116 16940 18126 16996
rect 19404 16940 22652 16996
rect 22708 16940 22718 16996
rect 26562 16940 26572 16996
rect 26628 16940 27020 16996
rect 27076 16940 28028 16996
rect 28084 16940 28094 16996
rect 31938 16940 31948 16996
rect 32004 16940 32732 16996
rect 32788 16940 33796 16996
rect 34402 16940 34412 16996
rect 34468 16940 35196 16996
rect 35252 16940 36428 16996
rect 36484 16940 36494 16996
rect 39974 16940 40012 16996
rect 40068 16940 40078 16996
rect 40226 16940 40236 16996
rect 40292 16940 41692 16996
rect 41748 16940 41758 16996
rect 43586 16940 43596 16996
rect 43652 16940 44156 16996
rect 44212 16940 44222 16996
rect 44706 16940 44716 16996
rect 44772 16940 45052 16996
rect 45108 16940 45118 16996
rect 45378 16940 45388 16996
rect 45444 16940 45836 16996
rect 45892 16940 46732 16996
rect 46788 16940 49644 16996
rect 49700 16940 49710 16996
rect 50306 16940 50316 16996
rect 50372 16940 51548 16996
rect 51604 16940 51614 16996
rect 52994 16940 53004 16996
rect 53060 16940 57484 16996
rect 57540 16940 57550 16996
rect 200 16884 800 16912
rect 200 16828 2044 16884
rect 2100 16828 2110 16884
rect 4386 16828 4396 16884
rect 4452 16828 5180 16884
rect 5236 16828 6412 16884
rect 6468 16828 6478 16884
rect 7186 16828 7196 16884
rect 7252 16828 11732 16884
rect 13206 16828 13244 16884
rect 13300 16828 13310 16884
rect 16146 16828 16156 16884
rect 16212 16828 17948 16884
rect 18004 16828 18014 16884
rect 18806 16828 18844 16884
rect 18900 16828 18910 16884
rect 200 16800 800 16828
rect 11676 16772 11732 16828
rect 19404 16772 19460 16940
rect 33740 16884 33796 16940
rect 19590 16828 19628 16884
rect 19684 16828 19694 16884
rect 19954 16828 19964 16884
rect 20020 16828 20972 16884
rect 21028 16828 21038 16884
rect 21420 16828 23660 16884
rect 23716 16828 23726 16884
rect 25218 16828 25228 16884
rect 25284 16828 28812 16884
rect 28868 16828 29148 16884
rect 29204 16828 29214 16884
rect 32050 16828 32060 16884
rect 32116 16828 32508 16884
rect 32564 16828 33516 16884
rect 33572 16828 33582 16884
rect 33740 16828 35644 16884
rect 35700 16828 35710 16884
rect 37986 16828 37996 16884
rect 38052 16828 40124 16884
rect 40180 16828 40190 16884
rect 40338 16828 40348 16884
rect 40404 16828 40572 16884
rect 40628 16828 40638 16884
rect 41010 16828 41020 16884
rect 41076 16828 41132 16884
rect 41188 16828 41198 16884
rect 41570 16828 41580 16884
rect 41636 16828 46172 16884
rect 46228 16828 46238 16884
rect 47170 16828 47180 16884
rect 47236 16828 48188 16884
rect 48244 16828 50540 16884
rect 50596 16828 50606 16884
rect 53554 16828 53564 16884
rect 53620 16828 54012 16884
rect 54068 16828 55916 16884
rect 55972 16828 55982 16884
rect 21420 16772 21476 16828
rect 2482 16716 2492 16772
rect 2548 16716 4060 16772
rect 4116 16716 4126 16772
rect 5814 16716 5852 16772
rect 5908 16716 5918 16772
rect 7410 16716 7420 16772
rect 7476 16716 9772 16772
rect 9828 16716 9838 16772
rect 11676 16716 14924 16772
rect 14980 16716 14990 16772
rect 16034 16716 16044 16772
rect 16100 16716 16268 16772
rect 16324 16716 16334 16772
rect 18274 16716 18284 16772
rect 18340 16716 19460 16772
rect 21410 16716 21420 16772
rect 21476 16716 21486 16772
rect 23212 16716 24780 16772
rect 24836 16716 24846 16772
rect 23212 16660 23268 16716
rect 33740 16660 33796 16828
rect 50540 16772 50596 16828
rect 40562 16716 40572 16772
rect 40628 16716 40638 16772
rect 41122 16716 41132 16772
rect 41188 16716 41468 16772
rect 41524 16716 41534 16772
rect 42466 16716 42476 16772
rect 42532 16716 45500 16772
rect 45556 16716 48076 16772
rect 48132 16716 48142 16772
rect 50540 16716 53340 16772
rect 53396 16716 53676 16772
rect 53732 16716 53742 16772
rect 58258 16716 58268 16772
rect 58324 16716 58492 16772
rect 58548 16716 58558 16772
rect 3574 16604 3612 16660
rect 3668 16604 3678 16660
rect 7410 16604 7420 16660
rect 7476 16604 7756 16660
rect 7812 16604 7822 16660
rect 8194 16604 8204 16660
rect 8260 16604 12348 16660
rect 12404 16604 12414 16660
rect 12898 16604 12908 16660
rect 12964 16604 15372 16660
rect 15428 16604 16156 16660
rect 16212 16604 16222 16660
rect 16482 16604 16492 16660
rect 16548 16604 19852 16660
rect 19908 16604 19918 16660
rect 20962 16604 20972 16660
rect 21028 16604 23268 16660
rect 23398 16604 23436 16660
rect 23492 16604 23502 16660
rect 26534 16604 26572 16660
rect 26628 16604 26638 16660
rect 33506 16604 33516 16660
rect 33572 16604 33796 16660
rect 40572 16660 40628 16716
rect 47180 16660 47236 16716
rect 40572 16604 43372 16660
rect 43428 16604 43820 16660
rect 43876 16604 43886 16660
rect 44594 16604 44604 16660
rect 44660 16604 45836 16660
rect 45892 16604 45902 16660
rect 47170 16604 47180 16660
rect 47236 16604 47246 16660
rect 47618 16604 47628 16660
rect 47684 16604 55020 16660
rect 55076 16604 55086 16660
rect 4834 16492 4844 16548
rect 4900 16492 6860 16548
rect 6916 16492 7308 16548
rect 7364 16492 7374 16548
rect 7522 16492 7532 16548
rect 7588 16492 8764 16548
rect 8820 16492 15148 16548
rect 19282 16492 19292 16548
rect 19348 16492 20188 16548
rect 20244 16492 20254 16548
rect 21074 16492 21084 16548
rect 21140 16492 21868 16548
rect 21924 16492 21934 16548
rect 23986 16492 23996 16548
rect 24052 16492 24556 16548
rect 24612 16492 24780 16548
rect 24836 16492 24846 16548
rect 24994 16492 25004 16548
rect 25060 16492 28924 16548
rect 28980 16492 28990 16548
rect 38406 16492 38444 16548
rect 38500 16492 38510 16548
rect 40562 16492 40572 16548
rect 40628 16492 42700 16548
rect 42756 16492 51884 16548
rect 51940 16492 51950 16548
rect 52658 16492 52668 16548
rect 52724 16492 54124 16548
rect 54180 16492 54190 16548
rect 58482 16492 58492 16548
rect 58548 16492 58828 16548
rect 58884 16492 58894 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 15092 16436 15148 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 8418 16380 8428 16436
rect 8484 16380 9324 16436
rect 9380 16380 12460 16436
rect 12516 16380 12526 16436
rect 15092 16380 16268 16436
rect 16324 16380 16334 16436
rect 23202 16380 23212 16436
rect 23268 16380 24276 16436
rect 25442 16380 25452 16436
rect 25508 16380 27916 16436
rect 27972 16380 28812 16436
rect 28868 16380 28878 16436
rect 36642 16380 36652 16436
rect 36708 16380 43484 16436
rect 43540 16380 43550 16436
rect 47842 16380 47852 16436
rect 47908 16380 48748 16436
rect 48804 16380 49532 16436
rect 49588 16380 49598 16436
rect 51314 16380 51324 16436
rect 51380 16380 53788 16436
rect 53844 16380 53854 16436
rect 24220 16324 24276 16380
rect 2594 16268 2604 16324
rect 2660 16268 9660 16324
rect 9716 16268 9726 16324
rect 10332 16268 11788 16324
rect 11844 16268 15148 16324
rect 15810 16268 15820 16324
rect 15876 16268 16044 16324
rect 16100 16268 23548 16324
rect 23604 16268 23614 16324
rect 24210 16268 24220 16324
rect 24276 16268 30828 16324
rect 30884 16268 30894 16324
rect 37986 16268 37996 16324
rect 38052 16268 39116 16324
rect 39172 16268 39340 16324
rect 39396 16268 39406 16324
rect 39666 16268 39676 16324
rect 39732 16268 40460 16324
rect 40516 16268 40908 16324
rect 40964 16268 40974 16324
rect 46610 16268 46620 16324
rect 46676 16268 51436 16324
rect 51492 16268 53228 16324
rect 53284 16268 53294 16324
rect 57334 16268 57372 16324
rect 57428 16268 57438 16324
rect 1250 16156 1260 16212
rect 1316 16156 4620 16212
rect 4676 16156 4686 16212
rect 4844 16156 7084 16212
rect 7140 16156 7150 16212
rect 8418 16156 8428 16212
rect 8484 16156 9100 16212
rect 9156 16156 9166 16212
rect 4134 16044 4172 16100
rect 4228 16044 4238 16100
rect 4844 15988 4900 16156
rect 10332 16100 10388 16268
rect 15092 16212 15148 16268
rect 12898 16156 12908 16212
rect 12964 16156 13356 16212
rect 13412 16156 13422 16212
rect 15092 16156 16156 16212
rect 16212 16156 17052 16212
rect 17108 16156 17118 16212
rect 18274 16156 18284 16212
rect 18340 16156 21084 16212
rect 21140 16156 21150 16212
rect 21980 16156 23660 16212
rect 23716 16156 23726 16212
rect 34514 16156 34524 16212
rect 34580 16156 35308 16212
rect 35364 16156 36540 16212
rect 36596 16156 36606 16212
rect 37874 16156 37884 16212
rect 37940 16156 38500 16212
rect 39218 16156 39228 16212
rect 39284 16156 39564 16212
rect 39620 16156 39630 16212
rect 42354 16156 42364 16212
rect 42420 16156 44492 16212
rect 44548 16156 44558 16212
rect 45378 16156 45388 16212
rect 45444 16156 46508 16212
rect 46564 16156 46574 16212
rect 46834 16156 46844 16212
rect 46900 16156 48300 16212
rect 48356 16156 48366 16212
rect 49298 16156 49308 16212
rect 49364 16156 52220 16212
rect 52276 16156 52286 16212
rect 52882 16156 52892 16212
rect 52948 16156 53564 16212
rect 53620 16156 53630 16212
rect 54674 16156 54684 16212
rect 54740 16156 58268 16212
rect 58324 16156 58334 16212
rect 21980 16100 22036 16156
rect 5058 16044 5068 16100
rect 5124 16044 10388 16100
rect 10546 16044 10556 16100
rect 10612 16044 11340 16100
rect 11396 16044 11406 16100
rect 12002 16044 12012 16100
rect 12068 16044 13020 16100
rect 13076 16044 13086 16100
rect 18722 16044 18732 16100
rect 18788 16044 19068 16100
rect 19124 16044 19134 16100
rect 20514 16044 20524 16100
rect 20580 16044 22036 16100
rect 23314 16044 23324 16100
rect 23380 16044 23548 16100
rect 23604 16044 23614 16100
rect 24518 16044 24556 16100
rect 24612 16044 24622 16100
rect 24770 16044 24780 16100
rect 24836 16044 25116 16100
rect 25172 16044 25182 16100
rect 26450 16044 26460 16100
rect 26516 16044 26572 16100
rect 26628 16044 26638 16100
rect 29894 16044 29932 16100
rect 29988 16044 30380 16100
rect 30436 16044 30828 16100
rect 30884 16044 30894 16100
rect 34626 16044 34636 16100
rect 34692 16044 35084 16100
rect 35140 16044 35150 16100
rect 35746 16044 35756 16100
rect 35812 16044 35980 16100
rect 36036 16044 36988 16100
rect 37044 16044 38108 16100
rect 38164 16044 38174 16100
rect 4274 15932 4284 15988
rect 4340 15932 4900 15988
rect 5730 15932 5740 15988
rect 5796 15932 6636 15988
rect 6692 15932 6702 15988
rect 7410 15932 7420 15988
rect 7476 15932 7980 15988
rect 8036 15932 10668 15988
rect 10724 15932 10734 15988
rect 16370 15932 16380 15988
rect 16436 15932 17836 15988
rect 17892 15932 17902 15988
rect 18386 15932 18396 15988
rect 18452 15932 21756 15988
rect 21812 15932 21822 15988
rect 22082 15932 22092 15988
rect 22148 15932 22988 15988
rect 23044 15932 23054 15988
rect 23314 15932 23324 15988
rect 23380 15932 25228 15988
rect 25284 15932 25294 15988
rect 26002 15932 26012 15988
rect 26068 15932 26908 15988
rect 26964 15932 26974 15988
rect 32946 15932 32956 15988
rect 33012 15932 34076 15988
rect 34132 15932 34860 15988
rect 34916 15932 36316 15988
rect 36372 15932 36382 15988
rect 36642 15932 36652 15988
rect 36708 15932 37660 15988
rect 37716 15932 37884 15988
rect 37940 15932 37950 15988
rect 21756 15876 21812 15932
rect 36316 15876 36372 15932
rect 38444 15876 38500 16156
rect 43586 16044 43596 16100
rect 43652 16044 43932 16100
rect 43988 16044 47628 16100
rect 47684 16044 47694 16100
rect 49568 16044 49644 16100
rect 49700 16044 51212 16100
rect 51268 16044 51278 16100
rect 54114 16044 54124 16100
rect 54180 16044 55356 16100
rect 55412 16044 55422 16100
rect 41010 15932 41020 15988
rect 41076 15932 42028 15988
rect 42084 15932 42094 15988
rect 44146 15932 44156 15988
rect 44212 15932 46620 15988
rect 46676 15932 46686 15988
rect 50754 15932 50764 15988
rect 50820 15932 53676 15988
rect 53732 15932 54460 15988
rect 54516 15932 54526 15988
rect 3602 15820 3612 15876
rect 3668 15820 7532 15876
rect 7588 15820 7598 15876
rect 8978 15820 8988 15876
rect 9044 15820 13132 15876
rect 13188 15820 13804 15876
rect 13860 15820 17948 15876
rect 18004 15820 18014 15876
rect 19394 15820 19404 15876
rect 19460 15820 19516 15876
rect 19572 15820 19582 15876
rect 21756 15820 24780 15876
rect 24836 15820 24846 15876
rect 30818 15820 30828 15876
rect 30884 15820 31724 15876
rect 31780 15820 31790 15876
rect 36316 15820 37548 15876
rect 37604 15820 37614 15876
rect 38434 15820 38444 15876
rect 38500 15820 38510 15876
rect 39824 15820 39900 15876
rect 39956 15820 41132 15876
rect 41188 15820 41198 15876
rect 45826 15820 45836 15876
rect 45892 15820 48972 15876
rect 49028 15820 49038 15876
rect 50418 15820 50428 15876
rect 50484 15820 51212 15876
rect 51268 15820 51278 15876
rect 54898 15820 54908 15876
rect 54964 15820 56252 15876
rect 56308 15820 56924 15876
rect 56980 15820 57484 15876
rect 57540 15820 57932 15876
rect 57988 15820 57998 15876
rect 2706 15708 2716 15764
rect 2772 15708 8092 15764
rect 8148 15708 8876 15764
rect 8932 15708 8942 15764
rect 9090 15708 9100 15764
rect 9156 15708 12124 15764
rect 12180 15708 12190 15764
rect 14242 15708 14252 15764
rect 14308 15708 16380 15764
rect 16436 15708 17836 15764
rect 17892 15708 17902 15764
rect 18274 15708 18284 15764
rect 18340 15708 19628 15764
rect 19684 15708 19694 15764
rect 23314 15708 23324 15764
rect 23380 15708 24220 15764
rect 24276 15708 24286 15764
rect 26608 15708 26684 15764
rect 26740 15708 29484 15764
rect 29540 15708 29550 15764
rect 37062 15708 37100 15764
rect 37156 15708 37166 15764
rect 38658 15708 38668 15764
rect 38724 15708 38762 15764
rect 49746 15708 49756 15764
rect 49812 15708 50316 15764
rect 50372 15708 50382 15764
rect 51314 15708 51324 15764
rect 51380 15708 51884 15764
rect 51940 15708 51996 15764
rect 52052 15708 52062 15764
rect 52210 15708 52220 15764
rect 52276 15708 52780 15764
rect 52836 15708 52846 15764
rect 53666 15708 53676 15764
rect 53732 15708 57820 15764
rect 57876 15708 57886 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 2594 15596 2604 15652
rect 2660 15596 10220 15652
rect 10276 15596 10556 15652
rect 10612 15596 10622 15652
rect 12562 15596 12572 15652
rect 12628 15596 13356 15652
rect 13412 15596 13422 15652
rect 13794 15596 13804 15652
rect 13860 15596 16044 15652
rect 16100 15596 16110 15652
rect 16706 15596 16716 15652
rect 16772 15596 17052 15652
rect 17108 15596 18732 15652
rect 18788 15596 18798 15652
rect 19170 15596 19180 15652
rect 19236 15596 19246 15652
rect 20514 15596 20524 15652
rect 20580 15596 22316 15652
rect 22372 15596 22382 15652
rect 28242 15596 28252 15652
rect 28308 15596 29596 15652
rect 29652 15596 29932 15652
rect 29988 15596 29998 15652
rect 34962 15596 34972 15652
rect 35028 15596 35644 15652
rect 35700 15596 35710 15652
rect 38332 15596 42364 15652
rect 42420 15596 43260 15652
rect 43316 15596 43326 15652
rect 46050 15596 46060 15652
rect 46116 15596 46126 15652
rect 46274 15596 46284 15652
rect 46340 15596 46396 15652
rect 46452 15596 46462 15652
rect 47730 15596 47740 15652
rect 47796 15596 49308 15652
rect 49364 15596 49374 15652
rect 51660 15596 53452 15652
rect 53508 15596 55468 15652
rect 55524 15596 55534 15652
rect 19180 15540 19236 15596
rect 38332 15540 38388 15596
rect 46060 15540 46116 15596
rect 51660 15540 51716 15596
rect 3938 15484 3948 15540
rect 4004 15484 4844 15540
rect 4900 15484 4910 15540
rect 5282 15484 5292 15540
rect 5348 15484 5404 15540
rect 5460 15484 6412 15540
rect 6468 15484 6478 15540
rect 7634 15484 7644 15540
rect 7700 15484 7710 15540
rect 8642 15484 8652 15540
rect 8708 15484 14700 15540
rect 14756 15484 14766 15540
rect 15138 15484 15148 15540
rect 15204 15484 16324 15540
rect 16482 15484 16492 15540
rect 16548 15484 17500 15540
rect 17556 15484 17566 15540
rect 18134 15484 18172 15540
rect 18228 15484 18620 15540
rect 18676 15484 18686 15540
rect 19180 15484 19796 15540
rect 20514 15484 20524 15540
rect 20580 15484 20590 15540
rect 21410 15484 21420 15540
rect 21476 15484 21644 15540
rect 21700 15484 21710 15540
rect 22418 15484 22428 15540
rect 22484 15484 22988 15540
rect 23044 15484 23054 15540
rect 23538 15484 23548 15540
rect 23604 15484 24556 15540
rect 24612 15484 24780 15540
rect 24836 15484 24846 15540
rect 29250 15484 29260 15540
rect 29316 15484 30604 15540
rect 30660 15484 30670 15540
rect 31686 15484 31724 15540
rect 31780 15484 32508 15540
rect 32564 15484 33740 15540
rect 33796 15484 34300 15540
rect 34356 15484 34366 15540
rect 37090 15484 37100 15540
rect 37156 15484 37772 15540
rect 37828 15484 37838 15540
rect 38098 15484 38108 15540
rect 38164 15484 38332 15540
rect 38388 15484 38398 15540
rect 38546 15484 38556 15540
rect 38612 15484 39228 15540
rect 39284 15484 39294 15540
rect 39526 15484 39564 15540
rect 39620 15484 39630 15540
rect 40450 15484 40460 15540
rect 40516 15484 40684 15540
rect 40740 15484 40750 15540
rect 44342 15484 44380 15540
rect 44436 15484 44446 15540
rect 46060 15484 46508 15540
rect 46564 15484 51716 15540
rect 51846 15484 51884 15540
rect 51940 15484 51950 15540
rect 54002 15484 54012 15540
rect 54068 15484 55580 15540
rect 55636 15484 55646 15540
rect 56550 15484 56588 15540
rect 56644 15484 56654 15540
rect 7644 15428 7700 15484
rect 16268 15428 16324 15484
rect 1922 15372 1932 15428
rect 1988 15372 3388 15428
rect 4722 15372 4732 15428
rect 4788 15372 5180 15428
rect 5236 15372 5246 15428
rect 6850 15372 6860 15428
rect 6916 15372 6972 15428
rect 7028 15372 7038 15428
rect 7186 15372 7196 15428
rect 7252 15372 9660 15428
rect 9716 15372 9726 15428
rect 9874 15372 9884 15428
rect 9940 15372 10780 15428
rect 10836 15372 10846 15428
rect 12898 15372 12908 15428
rect 12964 15372 13580 15428
rect 13636 15372 16044 15428
rect 16100 15372 16110 15428
rect 16268 15372 18844 15428
rect 18900 15372 19516 15428
rect 19572 15372 19582 15428
rect 3332 15316 3388 15372
rect 19740 15316 19796 15484
rect 20524 15428 20580 15484
rect 46060 15428 46116 15484
rect 20178 15372 20188 15428
rect 20244 15372 20300 15428
rect 20356 15372 23884 15428
rect 23940 15372 23950 15428
rect 24668 15372 25452 15428
rect 25508 15372 25518 15428
rect 42242 15372 42252 15428
rect 42308 15372 43708 15428
rect 43764 15372 46116 15428
rect 46946 15372 46956 15428
rect 47012 15372 47740 15428
rect 47796 15372 48188 15428
rect 48244 15372 48254 15428
rect 49298 15372 49308 15428
rect 49364 15372 50428 15428
rect 50484 15372 50494 15428
rect 52210 15372 52220 15428
rect 52276 15372 53004 15428
rect 53060 15372 53070 15428
rect 54674 15372 54684 15428
rect 54740 15372 55468 15428
rect 55524 15372 55534 15428
rect 24668 15316 24724 15372
rect 2706 15260 2716 15316
rect 2772 15260 3052 15316
rect 3108 15260 3118 15316
rect 3332 15260 7924 15316
rect 8082 15260 8092 15316
rect 8148 15260 11676 15316
rect 11732 15260 11742 15316
rect 16258 15260 16268 15316
rect 16324 15260 18396 15316
rect 18452 15260 18462 15316
rect 19740 15260 21084 15316
rect 21140 15260 21150 15316
rect 21858 15260 21868 15316
rect 21924 15260 24724 15316
rect 24882 15260 24892 15316
rect 24948 15260 25900 15316
rect 25956 15260 26572 15316
rect 26628 15260 26638 15316
rect 27234 15260 27244 15316
rect 27300 15260 27804 15316
rect 27860 15260 28588 15316
rect 28644 15260 28654 15316
rect 28802 15260 28812 15316
rect 28868 15260 29820 15316
rect 29876 15260 30380 15316
rect 30436 15260 30446 15316
rect 30818 15260 30828 15316
rect 30884 15260 32284 15316
rect 32340 15260 32350 15316
rect 32946 15260 32956 15316
rect 33012 15260 33516 15316
rect 33572 15260 33582 15316
rect 36530 15260 36540 15316
rect 36596 15260 37212 15316
rect 37268 15260 37996 15316
rect 38052 15260 38062 15316
rect 40450 15260 40460 15316
rect 40516 15260 40684 15316
rect 40740 15260 40750 15316
rect 41234 15260 41244 15316
rect 41300 15260 42028 15316
rect 42084 15260 42094 15316
rect 42914 15260 42924 15316
rect 42980 15260 43708 15316
rect 43764 15260 43774 15316
rect 46806 15260 46844 15316
rect 46900 15260 46910 15316
rect 48514 15260 48524 15316
rect 48580 15260 52668 15316
rect 52724 15260 52734 15316
rect 7868 15204 7924 15260
rect 28812 15204 28868 15260
rect 54684 15204 54740 15372
rect 55906 15260 55916 15316
rect 55972 15260 56364 15316
rect 56420 15260 57260 15316
rect 57316 15260 57326 15316
rect 57670 15260 57708 15316
rect 57764 15260 57774 15316
rect 1250 15148 1260 15204
rect 1316 15148 1708 15204
rect 1764 15148 1774 15204
rect 4134 15148 4172 15204
rect 4228 15148 4238 15204
rect 6850 15148 6860 15204
rect 6916 15148 7644 15204
rect 7700 15148 7710 15204
rect 7868 15148 8988 15204
rect 9044 15148 9054 15204
rect 12002 15148 12012 15204
rect 12068 15148 13020 15204
rect 13076 15148 13086 15204
rect 15026 15148 15036 15204
rect 15092 15148 22204 15204
rect 22260 15148 22270 15204
rect 23314 15148 23324 15204
rect 23380 15148 23436 15204
rect 23492 15148 23502 15204
rect 23650 15148 23660 15204
rect 23716 15148 23772 15204
rect 23828 15148 23838 15204
rect 27458 15148 27468 15204
rect 27524 15148 28868 15204
rect 30146 15148 30156 15204
rect 30212 15148 30716 15204
rect 30772 15148 31276 15204
rect 31332 15148 31342 15204
rect 40796 15148 42028 15204
rect 42084 15148 42094 15204
rect 43026 15148 43036 15204
rect 43092 15148 43932 15204
rect 43988 15148 43998 15204
rect 44156 15148 47740 15204
rect 47796 15148 47806 15204
rect 48514 15148 48524 15204
rect 48580 15148 48748 15204
rect 48804 15148 49756 15204
rect 49812 15148 49822 15204
rect 50866 15148 50876 15204
rect 50932 15148 50988 15204
rect 51044 15148 51054 15204
rect 52434 15148 52444 15204
rect 52500 15148 54740 15204
rect 40796 15092 40852 15148
rect 44156 15092 44212 15148
rect 1922 15036 1932 15092
rect 1988 15036 3388 15092
rect 3826 15036 3836 15092
rect 3892 15036 6748 15092
rect 6804 15036 6814 15092
rect 7410 15036 7420 15092
rect 7476 15036 11900 15092
rect 11956 15036 11966 15092
rect 12114 15036 12124 15092
rect 12180 15036 13804 15092
rect 13860 15036 13870 15092
rect 15922 15036 15932 15092
rect 15988 15036 19068 15092
rect 19124 15036 19134 15092
rect 29362 15036 29372 15092
rect 29428 15036 30044 15092
rect 30100 15036 30110 15092
rect 35074 15036 35084 15092
rect 35140 15036 36092 15092
rect 36148 15036 36158 15092
rect 40786 15036 40796 15092
rect 40852 15036 40862 15092
rect 43474 15036 43484 15092
rect 43540 15036 44212 15092
rect 44818 15036 44828 15092
rect 44884 15036 45276 15092
rect 45332 15036 45342 15092
rect 46274 15036 46284 15092
rect 46340 15036 46956 15092
rect 47012 15036 47022 15092
rect 50306 15036 50316 15092
rect 50372 15036 51100 15092
rect 51156 15036 51166 15092
rect 52322 15036 52332 15092
rect 52388 15036 54236 15092
rect 54292 15036 55692 15092
rect 55748 15036 55758 15092
rect 1698 14924 1708 14980
rect 1764 14924 2044 14980
rect 2100 14924 2110 14980
rect 3332 14756 3388 15036
rect 6748 14980 6804 15036
rect 4134 14924 4172 14980
rect 4228 14924 4238 14980
rect 4946 14924 4956 14980
rect 5012 14924 6524 14980
rect 6580 14924 6590 14980
rect 6748 14924 14252 14980
rect 14308 14924 14318 14980
rect 18498 14924 18508 14980
rect 18564 14924 19292 14980
rect 19348 14924 21084 14980
rect 21140 14924 21150 14980
rect 37062 14924 37100 14980
rect 37156 14924 37166 14980
rect 39554 14924 39564 14980
rect 39620 14924 48524 14980
rect 48580 14924 48590 14980
rect 54674 14924 54684 14980
rect 54740 14924 57708 14980
rect 57764 14924 57774 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 5730 14812 5740 14868
rect 5796 14812 8540 14868
rect 8596 14812 8606 14868
rect 9324 14812 11004 14868
rect 11060 14812 11676 14868
rect 11732 14812 11742 14868
rect 13682 14812 13692 14868
rect 13748 14812 15260 14868
rect 15316 14812 15326 14868
rect 17052 14812 21420 14868
rect 21476 14812 21486 14868
rect 21970 14812 21980 14868
rect 22036 14812 31164 14868
rect 31220 14812 31230 14868
rect 38658 14812 38668 14868
rect 38724 14812 43316 14868
rect 43474 14812 43484 14868
rect 43540 14812 43932 14868
rect 43988 14812 44380 14868
rect 44436 14812 47404 14868
rect 47460 14812 47470 14868
rect 57026 14812 57036 14868
rect 57092 14812 58828 14868
rect 58884 14812 59276 14868
rect 59332 14812 59342 14868
rect 9324 14756 9380 14812
rect 3332 14700 9380 14756
rect 9538 14700 9548 14756
rect 9604 14700 9660 14756
rect 9716 14700 9726 14756
rect 12114 14700 12124 14756
rect 12180 14700 12684 14756
rect 12740 14700 14028 14756
rect 14084 14700 14094 14756
rect 17052 14644 17108 14812
rect 43260 14756 43316 14812
rect 19842 14700 19852 14756
rect 19908 14700 21644 14756
rect 21700 14700 21710 14756
rect 36754 14700 36764 14756
rect 36820 14700 38892 14756
rect 38948 14700 38958 14756
rect 43260 14700 48412 14756
rect 48468 14700 48748 14756
rect 48804 14700 48814 14756
rect 2930 14588 2940 14644
rect 2996 14588 3612 14644
rect 3668 14588 3678 14644
rect 4284 14588 7420 14644
rect 7476 14588 7486 14644
rect 7606 14588 7644 14644
rect 7700 14588 7710 14644
rect 8642 14588 8652 14644
rect 8708 14588 13916 14644
rect 13972 14588 13982 14644
rect 16380 14588 17108 14644
rect 18050 14588 18060 14644
rect 18116 14588 18620 14644
rect 18676 14588 18686 14644
rect 19058 14588 19068 14644
rect 19124 14588 21532 14644
rect 21588 14588 21598 14644
rect 23062 14588 23100 14644
rect 23156 14588 23166 14644
rect 27010 14588 27020 14644
rect 27076 14588 29708 14644
rect 29764 14588 30268 14644
rect 30324 14588 30334 14644
rect 37314 14588 37324 14644
rect 37380 14588 38444 14644
rect 38500 14588 38510 14644
rect 39106 14588 39116 14644
rect 39172 14588 39788 14644
rect 39844 14588 41748 14644
rect 47842 14588 47852 14644
rect 47908 14588 48188 14644
rect 48244 14588 48254 14644
rect 49858 14588 49868 14644
rect 49924 14588 50316 14644
rect 50372 14588 50382 14644
rect 53330 14588 53340 14644
rect 53396 14588 57148 14644
rect 57204 14588 57214 14644
rect 4284 14532 4340 14588
rect 16380 14532 16436 14588
rect 18060 14532 18116 14588
rect 2818 14476 2828 14532
rect 2884 14476 2894 14532
rect 3602 14476 3612 14532
rect 3668 14476 4340 14532
rect 4498 14476 4508 14532
rect 4564 14476 6188 14532
rect 6244 14476 6254 14532
rect 6850 14476 6860 14532
rect 6916 14476 6972 14532
rect 7028 14476 7038 14532
rect 7186 14476 7196 14532
rect 7252 14476 8652 14532
rect 8708 14476 8718 14532
rect 8866 14476 8876 14532
rect 8932 14476 10444 14532
rect 10500 14476 10510 14532
rect 10658 14476 10668 14532
rect 10724 14476 11788 14532
rect 11844 14476 16436 14532
rect 16594 14476 16604 14532
rect 16660 14476 18116 14532
rect 19292 14476 19740 14532
rect 19796 14476 19806 14532
rect 19954 14476 19964 14532
rect 20020 14476 20524 14532
rect 20580 14476 20590 14532
rect 29474 14476 29484 14532
rect 29540 14476 30044 14532
rect 30100 14476 30828 14532
rect 30884 14476 30894 14532
rect 36306 14476 36316 14532
rect 36372 14476 38668 14532
rect 38724 14476 38734 14532
rect 39442 14476 39452 14532
rect 39508 14476 40460 14532
rect 40516 14476 40526 14532
rect 2828 14420 2884 14476
rect 19292 14420 19348 14476
rect 41692 14420 41748 14588
rect 46162 14476 46172 14532
rect 46228 14476 48972 14532
rect 49028 14476 49038 14532
rect 50978 14476 50988 14532
rect 51044 14476 51054 14532
rect 53666 14476 53676 14532
rect 53732 14476 53788 14532
rect 53844 14476 53854 14532
rect 54898 14476 54908 14532
rect 54964 14476 56140 14532
rect 56196 14476 57596 14532
rect 57652 14476 57662 14532
rect 2828 14364 5572 14420
rect 5730 14364 5740 14420
rect 5796 14364 6412 14420
rect 6468 14364 7532 14420
rect 7588 14364 7598 14420
rect 8530 14364 8540 14420
rect 8596 14364 9772 14420
rect 9828 14364 9838 14420
rect 10770 14364 10780 14420
rect 10836 14364 12012 14420
rect 12068 14364 12078 14420
rect 14914 14364 14924 14420
rect 14980 14364 16044 14420
rect 16100 14364 16110 14420
rect 18274 14364 18284 14420
rect 18340 14364 19348 14420
rect 19404 14364 20300 14420
rect 20356 14364 20366 14420
rect 22418 14364 22428 14420
rect 22484 14364 25564 14420
rect 25620 14364 25630 14420
rect 36530 14364 36540 14420
rect 36596 14364 37884 14420
rect 37940 14364 39004 14420
rect 39060 14364 41132 14420
rect 41188 14364 41198 14420
rect 41654 14364 41692 14420
rect 41748 14364 41758 14420
rect 42018 14364 42028 14420
rect 42084 14364 42924 14420
rect 42980 14364 43708 14420
rect 43764 14364 43774 14420
rect 45602 14364 45612 14420
rect 45668 14364 47684 14420
rect 48626 14364 48636 14420
rect 48692 14364 49588 14420
rect 5516 14308 5572 14364
rect 19404 14308 19460 14364
rect 47628 14308 47684 14364
rect 49532 14308 49588 14364
rect 50988 14308 51044 14476
rect 55682 14364 55692 14420
rect 55748 14364 56700 14420
rect 56756 14364 56766 14420
rect 3332 14252 3612 14308
rect 3668 14252 3678 14308
rect 3826 14252 3836 14308
rect 3892 14252 4060 14308
rect 4116 14252 4956 14308
rect 5012 14252 5022 14308
rect 5516 14252 7980 14308
rect 8036 14252 10332 14308
rect 10388 14252 11564 14308
rect 11620 14252 11630 14308
rect 12786 14252 12796 14308
rect 12852 14252 15932 14308
rect 15988 14252 15998 14308
rect 17938 14252 17948 14308
rect 18004 14252 18508 14308
rect 18564 14252 18956 14308
rect 19012 14252 19022 14308
rect 19170 14252 19180 14308
rect 19236 14252 19460 14308
rect 20066 14252 20076 14308
rect 20132 14252 20636 14308
rect 20692 14252 21532 14308
rect 21588 14252 22092 14308
rect 22148 14252 23212 14308
rect 23268 14252 23278 14308
rect 23426 14252 23436 14308
rect 23492 14252 24332 14308
rect 24388 14252 24398 14308
rect 27906 14252 27916 14308
rect 27972 14252 28476 14308
rect 28532 14252 28542 14308
rect 30594 14252 30604 14308
rect 30660 14252 33516 14308
rect 33572 14252 33582 14308
rect 34290 14252 34300 14308
rect 34356 14252 44044 14308
rect 44100 14252 44110 14308
rect 44482 14252 44492 14308
rect 44548 14252 47068 14308
rect 47124 14252 47134 14308
rect 47618 14252 47628 14308
rect 47684 14252 48188 14308
rect 48244 14252 48636 14308
rect 48692 14252 48702 14308
rect 49494 14252 49532 14308
rect 49588 14252 49598 14308
rect 50642 14252 50652 14308
rect 50708 14252 53340 14308
rect 53396 14252 53406 14308
rect 55990 14252 56028 14308
rect 56084 14252 58380 14308
rect 58436 14252 58446 14308
rect 3332 14196 3388 14252
rect 59200 14196 59800 14224
rect 2482 14140 2492 14196
rect 2548 14140 3388 14196
rect 3490 14140 3500 14196
rect 3556 14140 11116 14196
rect 11172 14140 14476 14196
rect 14532 14140 14542 14196
rect 15092 14140 19068 14196
rect 19124 14140 19628 14196
rect 19684 14140 19694 14196
rect 23286 14140 23324 14196
rect 23380 14140 23390 14196
rect 38994 14140 39004 14196
rect 39060 14140 39340 14196
rect 39396 14140 40124 14196
rect 40180 14140 40190 14196
rect 42690 14140 42700 14196
rect 42756 14140 43820 14196
rect 43876 14140 45276 14196
rect 45332 14140 45836 14196
rect 45892 14140 45902 14196
rect 46610 14140 46620 14196
rect 46676 14140 46732 14196
rect 46788 14140 46798 14196
rect 49410 14140 49420 14196
rect 49476 14140 49644 14196
rect 49700 14140 49710 14196
rect 52098 14140 52108 14196
rect 52164 14140 53564 14196
rect 53620 14140 53630 14196
rect 55346 14140 55356 14196
rect 55412 14140 59800 14196
rect 15092 14084 15148 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 39004 14084 39060 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 59200 14112 59800 14140
rect 2930 14028 2940 14084
rect 2996 14028 5292 14084
rect 5348 14028 5358 14084
rect 6822 14028 6860 14084
rect 6916 14028 6926 14084
rect 7410 14028 7420 14084
rect 7476 14028 10332 14084
rect 10388 14028 12572 14084
rect 12628 14028 12638 14084
rect 13234 14028 13244 14084
rect 13300 14028 13692 14084
rect 13748 14028 13758 14084
rect 13906 14028 13916 14084
rect 13972 14028 15148 14084
rect 15586 14028 15596 14084
rect 15652 14028 18340 14084
rect 19058 14028 19068 14084
rect 19124 14028 19516 14084
rect 19572 14028 19582 14084
rect 22978 14028 22988 14084
rect 23044 14028 23436 14084
rect 23492 14028 23502 14084
rect 24322 14028 24332 14084
rect 24388 14028 30492 14084
rect 30548 14028 31724 14084
rect 31780 14028 31790 14084
rect 32732 14028 39060 14084
rect 18284 13972 18340 14028
rect 32732 13972 32788 14028
rect 2706 13916 2716 13972
rect 2772 13916 3500 13972
rect 3556 13916 3566 13972
rect 4498 13916 4508 13972
rect 4564 13916 5068 13972
rect 5124 13916 5134 13972
rect 5282 13916 5292 13972
rect 5348 13916 5740 13972
rect 5796 13916 7756 13972
rect 7812 13916 7822 13972
rect 8082 13916 8092 13972
rect 8148 13916 13468 13972
rect 13524 13916 13534 13972
rect 14690 13916 14700 13972
rect 14756 13916 15148 13972
rect 15204 13916 15214 13972
rect 15698 13916 15708 13972
rect 15764 13916 15932 13972
rect 15988 13916 15998 13972
rect 16342 13916 16380 13972
rect 16436 13916 16446 13972
rect 16818 13916 16828 13972
rect 16884 13916 17612 13972
rect 17668 13916 17678 13972
rect 18284 13916 19740 13972
rect 19796 13916 19806 13972
rect 23650 13916 23660 13972
rect 23716 13916 24220 13972
rect 24276 13916 24780 13972
rect 24836 13916 24846 13972
rect 30930 13916 30940 13972
rect 30996 13916 32788 13972
rect 33394 13916 33404 13972
rect 33460 13916 33628 13972
rect 33684 13916 34412 13972
rect 34468 13916 34478 13972
rect 36978 13916 36988 13972
rect 37044 13916 37660 13972
rect 37716 13916 37726 13972
rect 42242 13916 42252 13972
rect 42308 13916 43484 13972
rect 43540 13916 43550 13972
rect 44146 13916 44156 13972
rect 44212 13916 44268 13972
rect 44324 13916 44334 13972
rect 45238 13916 45276 13972
rect 45332 13916 45342 13972
rect 46386 13916 46396 13972
rect 46452 13916 46508 13972
rect 46564 13916 46574 13972
rect 51090 13916 51100 13972
rect 51156 13916 51772 13972
rect 51828 13916 56364 13972
rect 56420 13916 56430 13972
rect 46396 13860 46452 13916
rect 5058 13804 5068 13860
rect 5124 13804 6188 13860
rect 6244 13804 6254 13860
rect 6514 13804 6524 13860
rect 6580 13804 7644 13860
rect 7700 13804 8652 13860
rect 8708 13804 8718 13860
rect 8866 13804 8876 13860
rect 8932 13804 9772 13860
rect 9828 13804 9838 13860
rect 10108 13804 16436 13860
rect 18722 13804 18732 13860
rect 18788 13804 19180 13860
rect 19236 13804 19246 13860
rect 44482 13804 44492 13860
rect 44548 13804 46452 13860
rect 49074 13804 49084 13860
rect 49140 13804 49644 13860
rect 49700 13804 52108 13860
rect 52164 13804 52174 13860
rect 53190 13804 53228 13860
rect 53284 13804 56140 13860
rect 56196 13804 56206 13860
rect 10108 13748 10164 13804
rect 16380 13748 16436 13804
rect 4162 13692 4172 13748
rect 4228 13692 5180 13748
rect 5236 13692 5246 13748
rect 6626 13692 6636 13748
rect 6692 13692 7756 13748
rect 7812 13692 7822 13748
rect 8194 13692 8204 13748
rect 8260 13692 10164 13748
rect 10556 13692 14252 13748
rect 14308 13692 14318 13748
rect 14466 13692 14476 13748
rect 14532 13692 15148 13748
rect 15204 13692 15214 13748
rect 15474 13692 15484 13748
rect 15540 13692 15708 13748
rect 15764 13692 15774 13748
rect 16380 13692 22428 13748
rect 22484 13692 22494 13748
rect 26338 13692 26348 13748
rect 26404 13692 30380 13748
rect 30436 13692 30446 13748
rect 35298 13692 35308 13748
rect 35364 13692 36540 13748
rect 36596 13692 36606 13748
rect 44034 13692 44044 13748
rect 44100 13692 52108 13748
rect 52164 13692 52174 13748
rect 52322 13692 52332 13748
rect 52388 13692 53116 13748
rect 53172 13692 53182 13748
rect 54450 13692 54460 13748
rect 54516 13692 55020 13748
rect 55076 13692 55692 13748
rect 55748 13692 55758 13748
rect 2370 13580 2380 13636
rect 2436 13580 9212 13636
rect 9268 13580 9278 13636
rect 2818 13468 2828 13524
rect 2884 13468 4844 13524
rect 4900 13468 4956 13524
rect 5012 13468 5022 13524
rect 5282 13468 5292 13524
rect 5348 13468 5964 13524
rect 6020 13468 6030 13524
rect 8204 13468 8316 13524
rect 8372 13468 8382 13524
rect 8754 13468 8764 13524
rect 8820 13468 10332 13524
rect 10388 13468 10398 13524
rect 8204 13412 8260 13468
rect 4844 13356 8260 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 4844 13188 4900 13356
rect 10556 13300 10612 13692
rect 11218 13580 11228 13636
rect 11284 13580 12012 13636
rect 12068 13580 13468 13636
rect 13524 13580 13534 13636
rect 14578 13580 14588 13636
rect 14644 13580 15260 13636
rect 15316 13580 15326 13636
rect 15586 13580 15596 13636
rect 15652 13580 17052 13636
rect 17108 13580 17118 13636
rect 17714 13580 17724 13636
rect 17780 13580 18284 13636
rect 18340 13580 18350 13636
rect 18722 13580 18732 13636
rect 18788 13580 19180 13636
rect 19236 13580 19246 13636
rect 21186 13580 21196 13636
rect 21252 13580 23436 13636
rect 23492 13580 23502 13636
rect 27346 13580 27356 13636
rect 27412 13580 27804 13636
rect 27860 13580 29932 13636
rect 29988 13580 31388 13636
rect 31444 13580 31454 13636
rect 37202 13580 37212 13636
rect 37268 13580 37772 13636
rect 37828 13580 37838 13636
rect 38770 13580 38780 13636
rect 38836 13580 41356 13636
rect 41412 13580 41422 13636
rect 41570 13580 41580 13636
rect 41636 13580 41916 13636
rect 41972 13580 42700 13636
rect 42756 13580 42766 13636
rect 47058 13580 47068 13636
rect 47124 13580 47162 13636
rect 49858 13580 49868 13636
rect 49924 13580 51660 13636
rect 51716 13580 51726 13636
rect 51986 13580 51996 13636
rect 52052 13580 53900 13636
rect 53956 13580 53966 13636
rect 54226 13580 54236 13636
rect 54292 13580 54908 13636
rect 54964 13580 54974 13636
rect 11554 13468 11564 13524
rect 11620 13468 17388 13524
rect 17444 13468 17454 13524
rect 17948 13468 28252 13524
rect 28308 13468 28318 13524
rect 31938 13468 31948 13524
rect 32004 13468 33852 13524
rect 33908 13468 33918 13524
rect 38658 13468 38668 13524
rect 38724 13468 39788 13524
rect 39844 13468 40180 13524
rect 40338 13468 40348 13524
rect 40404 13468 43540 13524
rect 43810 13468 43820 13524
rect 43876 13468 44604 13524
rect 44660 13468 44670 13524
rect 46946 13468 46956 13524
rect 17948 13412 18004 13468
rect 40124 13412 40180 13468
rect 43484 13412 43540 13468
rect 47012 13412 47068 13524
rect 48178 13468 48188 13524
rect 48244 13468 50204 13524
rect 50260 13468 50270 13524
rect 51090 13468 51100 13524
rect 51156 13468 53900 13524
rect 53956 13468 53966 13524
rect 55570 13468 55580 13524
rect 55636 13468 59500 13524
rect 59556 13468 59566 13524
rect 12114 13356 12124 13412
rect 12180 13356 13580 13412
rect 13636 13356 17948 13412
rect 18004 13356 18014 13412
rect 20290 13356 20300 13412
rect 20356 13356 20748 13412
rect 20804 13356 22540 13412
rect 22596 13356 22606 13412
rect 38546 13356 38556 13412
rect 38612 13356 39116 13412
rect 39172 13356 39676 13412
rect 39732 13356 39742 13412
rect 40124 13356 40572 13412
rect 40628 13356 40908 13412
rect 40964 13356 40974 13412
rect 43474 13356 43484 13412
rect 43540 13356 43550 13412
rect 44482 13356 44492 13412
rect 44548 13356 44716 13412
rect 44772 13356 44782 13412
rect 47012 13356 47852 13412
rect 47908 13356 47918 13412
rect 50194 13356 50204 13412
rect 50260 13356 50428 13412
rect 50484 13356 50494 13412
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 5618 13244 5628 13300
rect 5684 13244 7868 13300
rect 7924 13244 10612 13300
rect 12338 13244 12348 13300
rect 12404 13244 21532 13300
rect 21588 13244 21868 13300
rect 21924 13244 21934 13300
rect 22418 13244 22428 13300
rect 22484 13244 22876 13300
rect 22932 13244 23436 13300
rect 23492 13244 23502 13300
rect 25218 13244 25228 13300
rect 25284 13244 26348 13300
rect 26404 13244 27020 13300
rect 27076 13244 27086 13300
rect 41682 13244 41692 13300
rect 41748 13244 48860 13300
rect 48916 13244 48926 13300
rect 51090 13244 51100 13300
rect 51156 13244 55580 13300
rect 55636 13244 55646 13300
rect 1922 13132 1932 13188
rect 1988 13132 3500 13188
rect 3556 13132 3566 13188
rect 4610 13132 4620 13188
rect 4676 13132 4900 13188
rect 5394 13132 5404 13188
rect 5460 13132 5852 13188
rect 5908 13132 5918 13188
rect 13346 13132 13356 13188
rect 13412 13132 15036 13188
rect 15092 13132 15102 13188
rect 15250 13132 15260 13188
rect 15316 13132 16828 13188
rect 16884 13132 18732 13188
rect 18788 13132 18798 13188
rect 18946 13132 18956 13188
rect 19012 13132 19628 13188
rect 19684 13132 22988 13188
rect 23044 13132 23054 13188
rect 36754 13132 36764 13188
rect 36820 13132 37324 13188
rect 37380 13132 42028 13188
rect 42084 13132 42140 13188
rect 42196 13132 42206 13188
rect 42364 13132 55916 13188
rect 55972 13132 56364 13188
rect 56420 13132 56430 13188
rect 42364 13076 42420 13132
rect 1474 13020 1484 13076
rect 1540 13020 6636 13076
rect 6692 13020 6702 13076
rect 7718 13020 7756 13076
rect 7812 13020 7822 13076
rect 8082 13020 8092 13076
rect 8148 13020 9940 13076
rect 10098 13020 10108 13076
rect 10164 13020 16380 13076
rect 16436 13020 16446 13076
rect 17826 13020 17836 13076
rect 17892 13020 20188 13076
rect 20244 13020 21308 13076
rect 21364 13020 21644 13076
rect 21700 13020 21710 13076
rect 29810 13020 29820 13076
rect 29876 13020 30492 13076
rect 30548 13020 30828 13076
rect 30884 13020 30894 13076
rect 34626 13020 34636 13076
rect 34692 13020 35196 13076
rect 35252 13020 35262 13076
rect 39666 13020 39676 13076
rect 39732 13020 42420 13076
rect 43026 13020 43036 13076
rect 43092 13020 46060 13076
rect 46116 13020 47292 13076
rect 47348 13020 47358 13076
rect 48962 13020 48972 13076
rect 49028 13020 49700 13076
rect 51986 13020 51996 13076
rect 52052 13020 55804 13076
rect 55860 13020 55870 13076
rect 57810 13020 57820 13076
rect 57876 13020 59052 13076
rect 59108 13020 59118 13076
rect 9884 12964 9940 13020
rect 49644 12964 49700 13020
rect 1362 12908 1372 12964
rect 1428 12908 2044 12964
rect 2100 12908 2380 12964
rect 2436 12908 2446 12964
rect 3266 12908 3276 12964
rect 3332 12908 4620 12964
rect 4676 12908 4686 12964
rect 4946 12908 4956 12964
rect 5012 12908 6188 12964
rect 6244 12908 6254 12964
rect 7158 12908 7196 12964
rect 7252 12908 7262 12964
rect 9090 12908 9100 12964
rect 9156 12908 9660 12964
rect 9716 12908 9726 12964
rect 9884 12908 12964 12964
rect 16034 12908 16044 12964
rect 16100 12908 20300 12964
rect 20356 12908 20366 12964
rect 20514 12908 20524 12964
rect 20580 12908 21980 12964
rect 22036 12908 22046 12964
rect 25330 12908 25340 12964
rect 25396 12908 31276 12964
rect 31332 12908 31342 12964
rect 32834 12908 32844 12964
rect 32900 12908 33628 12964
rect 33684 12908 33694 12964
rect 39106 12908 39116 12964
rect 39172 12908 40236 12964
rect 40292 12908 40302 12964
rect 40562 12908 40572 12964
rect 40628 12908 41020 12964
rect 41076 12908 41086 12964
rect 46386 12908 46396 12964
rect 46452 12908 47628 12964
rect 47684 12908 47964 12964
rect 48020 12908 48636 12964
rect 48692 12908 48702 12964
rect 49644 12908 51100 12964
rect 51156 12908 51166 12964
rect 51762 12908 51772 12964
rect 51828 12908 52668 12964
rect 52724 12908 52734 12964
rect 12908 12852 12964 12908
rect 3602 12796 3612 12852
rect 3668 12796 4284 12852
rect 4340 12796 5852 12852
rect 5908 12796 5918 12852
rect 6178 12796 6188 12852
rect 6244 12796 12684 12852
rect 12740 12796 12750 12852
rect 12898 12796 12908 12852
rect 12964 12796 15036 12852
rect 15092 12796 19404 12852
rect 19460 12796 19470 12852
rect 20738 12796 20748 12852
rect 20804 12796 24220 12852
rect 24276 12796 24286 12852
rect 26572 12740 26628 12908
rect 28466 12796 28476 12852
rect 28532 12796 29820 12852
rect 29876 12796 29886 12852
rect 33282 12796 33292 12852
rect 33348 12796 33740 12852
rect 33796 12796 34524 12852
rect 34580 12796 34590 12852
rect 39414 12796 39452 12852
rect 39508 12796 39518 12852
rect 40898 12796 40908 12852
rect 40964 12796 41132 12852
rect 41188 12796 41804 12852
rect 41860 12796 41870 12852
rect 48738 12796 48748 12852
rect 48804 12796 49196 12852
rect 49252 12796 49262 12852
rect 49606 12796 49644 12852
rect 49700 12796 51436 12852
rect 51492 12796 51502 12852
rect 52322 12796 52332 12852
rect 52388 12796 54684 12852
rect 54740 12796 54750 12852
rect 57026 12796 57036 12852
rect 57092 12796 57932 12852
rect 57988 12796 58380 12852
rect 58436 12796 58446 12852
rect 8082 12684 8092 12740
rect 8148 12684 9324 12740
rect 9380 12684 10108 12740
rect 10164 12684 10174 12740
rect 13794 12684 13804 12740
rect 13860 12684 15820 12740
rect 15876 12684 15886 12740
rect 16146 12684 16156 12740
rect 16212 12684 16268 12740
rect 16324 12684 16334 12740
rect 18722 12684 18732 12740
rect 18788 12684 19180 12740
rect 19236 12684 19246 12740
rect 19618 12684 19628 12740
rect 19684 12684 19740 12740
rect 19796 12684 19806 12740
rect 21382 12684 21420 12740
rect 21476 12684 21486 12740
rect 23090 12684 23100 12740
rect 23156 12684 23324 12740
rect 23380 12684 23390 12740
rect 26562 12684 26572 12740
rect 26628 12684 26638 12740
rect 36866 12684 36876 12740
rect 36932 12684 40124 12740
rect 40180 12684 41580 12740
rect 41636 12684 41646 12740
rect 44818 12684 44828 12740
rect 44884 12684 46172 12740
rect 46228 12684 52108 12740
rect 52164 12684 54124 12740
rect 54180 12684 54190 12740
rect 5058 12572 5068 12628
rect 5124 12572 11676 12628
rect 11732 12572 12572 12628
rect 12628 12572 13020 12628
rect 13076 12572 13916 12628
rect 13972 12572 13982 12628
rect 14242 12572 14252 12628
rect 14308 12572 14924 12628
rect 14980 12572 14990 12628
rect 16258 12572 16268 12628
rect 16324 12572 17388 12628
rect 17444 12572 17454 12628
rect 18498 12572 18508 12628
rect 18564 12572 18620 12628
rect 18676 12572 19236 12628
rect 26674 12572 26684 12628
rect 26740 12572 29708 12628
rect 29764 12572 29932 12628
rect 29988 12572 29998 12628
rect 38658 12572 38668 12628
rect 38724 12572 49532 12628
rect 49588 12572 49598 12628
rect 49746 12572 49756 12628
rect 49812 12572 49850 12628
rect 52322 12572 52332 12628
rect 52388 12572 52556 12628
rect 52612 12572 54348 12628
rect 54404 12572 54414 12628
rect 3714 12460 3724 12516
rect 3780 12460 3948 12516
rect 4004 12460 4014 12516
rect 4386 12460 4396 12516
rect 4452 12460 5628 12516
rect 5684 12460 5694 12516
rect 7298 12460 7308 12516
rect 7364 12460 12796 12516
rect 12852 12460 12862 12516
rect 16034 12460 16044 12516
rect 16100 12460 18060 12516
rect 18116 12460 18956 12516
rect 19012 12460 19022 12516
rect 3938 12348 3948 12404
rect 4004 12348 4956 12404
rect 5012 12348 5068 12404
rect 5124 12348 10220 12404
rect 10276 12348 10668 12404
rect 10724 12348 10734 12404
rect 11554 12348 11564 12404
rect 11620 12348 12236 12404
rect 12292 12348 13132 12404
rect 13188 12348 13198 12404
rect 15138 12348 15148 12404
rect 15204 12348 15242 12404
rect 15698 12348 15708 12404
rect 15764 12348 16828 12404
rect 16884 12348 16894 12404
rect 19180 12292 19236 12572
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 19394 12460 19404 12516
rect 19460 12460 19516 12516
rect 19572 12460 19582 12516
rect 43586 12460 43596 12516
rect 43652 12460 43932 12516
rect 43988 12460 43998 12516
rect 46134 12460 46172 12516
rect 46228 12460 46238 12516
rect 46498 12460 46508 12516
rect 46564 12460 46956 12516
rect 47012 12460 47022 12516
rect 48738 12460 48748 12516
rect 48804 12460 49644 12516
rect 49700 12460 50316 12516
rect 50372 12460 50382 12516
rect 19394 12348 19404 12404
rect 19460 12348 19852 12404
rect 19908 12348 19918 12404
rect 33964 12348 35644 12404
rect 35700 12348 36092 12404
rect 36148 12348 36158 12404
rect 40562 12348 40572 12404
rect 40628 12348 41468 12404
rect 41524 12348 41534 12404
rect 43698 12348 43708 12404
rect 43764 12348 44268 12404
rect 44324 12348 44334 12404
rect 45378 12348 45388 12404
rect 45444 12348 45454 12404
rect 45714 12348 45724 12404
rect 45780 12348 47740 12404
rect 47796 12348 47806 12404
rect 48738 12348 48748 12404
rect 48804 12348 50876 12404
rect 50932 12348 50942 12404
rect 55122 12348 55132 12404
rect 55188 12348 56588 12404
rect 56644 12348 56654 12404
rect 57362 12348 57372 12404
rect 57428 12348 58492 12404
rect 58548 12348 58558 12404
rect 33964 12292 34020 12348
rect 45388 12292 45444 12348
rect 5282 12236 5292 12292
rect 5348 12236 10556 12292
rect 10612 12236 11116 12292
rect 11172 12236 11182 12292
rect 12786 12236 12796 12292
rect 12852 12236 13468 12292
rect 13524 12236 16772 12292
rect 19170 12236 19180 12292
rect 19236 12236 21868 12292
rect 21924 12236 21934 12292
rect 22194 12236 22204 12292
rect 22260 12236 22876 12292
rect 22932 12236 22942 12292
rect 27458 12236 27468 12292
rect 27524 12236 28476 12292
rect 28532 12236 31164 12292
rect 31220 12236 31230 12292
rect 32834 12236 32844 12292
rect 32900 12236 33964 12292
rect 34020 12236 34030 12292
rect 34850 12236 34860 12292
rect 34916 12236 36316 12292
rect 36372 12236 36382 12292
rect 41010 12236 41020 12292
rect 41076 12236 42364 12292
rect 42420 12236 42700 12292
rect 42756 12236 46620 12292
rect 46676 12236 46686 12292
rect 47842 12236 47852 12292
rect 47908 12236 49868 12292
rect 49924 12236 50316 12292
rect 50372 12236 50382 12292
rect 16716 12180 16772 12236
rect 5954 12124 5964 12180
rect 6020 12124 6412 12180
rect 6468 12124 6972 12180
rect 7028 12124 7038 12180
rect 7634 12124 7644 12180
rect 7700 12124 8428 12180
rect 8484 12124 8494 12180
rect 9874 12124 9884 12180
rect 9940 12124 11228 12180
rect 11284 12124 11294 12180
rect 15026 12124 15036 12180
rect 15092 12124 16044 12180
rect 16100 12124 16110 12180
rect 16706 12124 16716 12180
rect 16772 12124 18172 12180
rect 18228 12124 18238 12180
rect 19058 12124 19068 12180
rect 19124 12124 22092 12180
rect 22148 12124 22158 12180
rect 24182 12124 24220 12180
rect 24276 12124 24286 12180
rect 28914 12124 28924 12180
rect 28980 12124 30716 12180
rect 30772 12124 30782 12180
rect 44594 12124 44604 12180
rect 44660 12124 45388 12180
rect 45444 12124 45454 12180
rect 51212 12124 54908 12180
rect 54964 12124 54974 12180
rect 51212 12068 51268 12124
rect 7298 12012 7308 12068
rect 7364 12012 8092 12068
rect 8148 12012 8158 12068
rect 10098 12012 10108 12068
rect 10164 12012 11004 12068
rect 11060 12012 11070 12068
rect 17042 12012 17052 12068
rect 17108 12012 26684 12068
rect 26740 12012 26750 12068
rect 41458 12012 41468 12068
rect 41524 12012 46172 12068
rect 46228 12012 47740 12068
rect 47796 12012 47806 12068
rect 51202 12012 51212 12068
rect 51268 12012 51278 12068
rect 53330 12012 53340 12068
rect 53396 12012 54348 12068
rect 54404 12012 55692 12068
rect 55748 12012 55758 12068
rect 15586 11900 15596 11956
rect 15652 11900 21980 11956
rect 22036 11900 22046 11956
rect 43698 11900 43708 11956
rect 43764 11900 47180 11956
rect 47236 11900 47246 11956
rect 49410 11900 49420 11956
rect 49476 11900 50540 11956
rect 50596 11900 54236 11956
rect 54292 11900 54302 11956
rect 8978 11788 8988 11844
rect 9044 11788 10444 11844
rect 10500 11788 11004 11844
rect 11060 11788 11844 11844
rect 12450 11788 12460 11844
rect 12516 11788 12908 11844
rect 12964 11788 16380 11844
rect 16436 11788 16446 11844
rect 19618 11788 19628 11844
rect 19684 11788 19852 11844
rect 19908 11788 19918 11844
rect 29474 11788 29484 11844
rect 29540 11788 29596 11844
rect 29652 11788 30268 11844
rect 30324 11788 32004 11844
rect 36866 11788 36876 11844
rect 36932 11788 38780 11844
rect 38836 11788 39116 11844
rect 39172 11788 39182 11844
rect 39442 11788 39452 11844
rect 39508 11788 40124 11844
rect 40180 11788 40190 11844
rect 49522 11788 49532 11844
rect 49588 11788 50764 11844
rect 50820 11788 50830 11844
rect 55010 11788 55020 11844
rect 55076 11788 57148 11844
rect 57204 11788 57214 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 11788 11732 11844 11788
rect 8306 11676 8316 11732
rect 8372 11676 9324 11732
rect 9380 11676 9390 11732
rect 11788 11676 15148 11732
rect 15250 11676 15260 11732
rect 15316 11676 16604 11732
rect 16660 11676 16670 11732
rect 16818 11676 16828 11732
rect 16884 11676 21196 11732
rect 21252 11676 21262 11732
rect 22082 11676 22092 11732
rect 22148 11676 23660 11732
rect 23716 11676 24108 11732
rect 24164 11676 24174 11732
rect 15092 11620 15148 11676
rect 31948 11620 32004 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 47058 11676 47068 11732
rect 47124 11676 48076 11732
rect 48132 11676 48636 11732
rect 48692 11676 48702 11732
rect 50082 11676 50092 11732
rect 50148 11676 50158 11732
rect 50306 11676 50316 11732
rect 50372 11676 50540 11732
rect 50596 11676 50606 11732
rect 51650 11676 51660 11732
rect 51716 11676 53340 11732
rect 53396 11676 53406 11732
rect 53564 11676 56924 11732
rect 56980 11676 56990 11732
rect 50092 11620 50148 11676
rect 53564 11620 53620 11676
rect 5058 11564 5068 11620
rect 5124 11564 8204 11620
rect 8260 11564 8270 11620
rect 8866 11564 8876 11620
rect 8932 11564 10948 11620
rect 11778 11564 11788 11620
rect 11844 11564 12012 11620
rect 12068 11564 14924 11620
rect 14980 11564 14990 11620
rect 15092 11564 19012 11620
rect 20962 11564 20972 11620
rect 21028 11564 26124 11620
rect 26180 11564 26190 11620
rect 31948 11564 41804 11620
rect 41860 11564 41870 11620
rect 48066 11564 48076 11620
rect 48132 11564 49868 11620
rect 49924 11564 49934 11620
rect 50092 11564 50652 11620
rect 50708 11564 50718 11620
rect 52032 11564 52108 11620
rect 52164 11564 53620 11620
rect 54898 11564 54908 11620
rect 54964 11564 55356 11620
rect 55412 11564 55422 11620
rect 200 11508 800 11536
rect 10892 11508 10948 11564
rect 18956 11508 19012 11564
rect 200 11452 1932 11508
rect 1988 11452 1998 11508
rect 3154 11452 3164 11508
rect 3220 11452 3388 11508
rect 3444 11452 3454 11508
rect 7970 11452 7980 11508
rect 8036 11452 10668 11508
rect 10724 11452 10734 11508
rect 10892 11452 11116 11508
rect 11172 11452 16940 11508
rect 16996 11452 17006 11508
rect 18946 11452 18956 11508
rect 19012 11452 22764 11508
rect 22820 11452 28028 11508
rect 28084 11452 28094 11508
rect 34402 11452 34412 11508
rect 34468 11452 35756 11508
rect 35812 11452 35822 11508
rect 37762 11452 37772 11508
rect 37828 11452 38892 11508
rect 38948 11452 38958 11508
rect 41682 11452 41692 11508
rect 41748 11452 42252 11508
rect 42308 11452 42318 11508
rect 42998 11452 43036 11508
rect 43092 11452 43102 11508
rect 44370 11452 44380 11508
rect 44436 11452 47628 11508
rect 47684 11452 47694 11508
rect 49410 11452 49420 11508
rect 49476 11452 50988 11508
rect 51044 11452 51054 11508
rect 53554 11452 53564 11508
rect 53620 11452 56252 11508
rect 56308 11452 56318 11508
rect 57362 11452 57372 11508
rect 57428 11452 57596 11508
rect 57652 11452 58940 11508
rect 58996 11452 59006 11508
rect 200 11424 800 11452
rect 2258 11340 2268 11396
rect 2324 11340 4060 11396
rect 4116 11340 4126 11396
rect 4274 11340 4284 11396
rect 4340 11340 4956 11396
rect 5012 11340 5022 11396
rect 6626 11340 6636 11396
rect 6692 11340 7420 11396
rect 7476 11340 7486 11396
rect 10434 11340 10444 11396
rect 10500 11340 13804 11396
rect 13860 11340 13870 11396
rect 14914 11340 14924 11396
rect 14980 11340 16604 11396
rect 16660 11340 16670 11396
rect 16818 11340 16828 11396
rect 16884 11340 18396 11396
rect 18452 11340 19628 11396
rect 19684 11340 19694 11396
rect 20738 11340 20748 11396
rect 20804 11340 21532 11396
rect 21588 11340 23212 11396
rect 23268 11340 23278 11396
rect 24658 11340 24668 11396
rect 24724 11340 25788 11396
rect 25844 11340 25854 11396
rect 26898 11340 26908 11396
rect 26964 11340 29036 11396
rect 29092 11340 29102 11396
rect 33058 11340 33068 11396
rect 33124 11340 37996 11396
rect 38052 11340 38668 11396
rect 38724 11340 38734 11396
rect 50372 11340 51324 11396
rect 51380 11340 51390 11396
rect 54786 11340 54796 11396
rect 54852 11340 56700 11396
rect 56756 11340 57484 11396
rect 57540 11340 57550 11396
rect 1810 11228 1820 11284
rect 1876 11228 8316 11284
rect 8372 11228 8382 11284
rect 10098 11228 10108 11284
rect 10164 11228 12348 11284
rect 12404 11228 12414 11284
rect 14130 11228 14140 11284
rect 14196 11228 14476 11284
rect 14532 11228 19180 11284
rect 19236 11228 25228 11284
rect 25284 11228 25294 11284
rect 27234 11228 27244 11284
rect 27300 11228 29596 11284
rect 29652 11228 29662 11284
rect 48850 11228 48860 11284
rect 48916 11228 50316 11284
rect 50372 11228 50428 11340
rect 53330 11228 53340 11284
rect 53396 11228 57372 11284
rect 57428 11228 57438 11284
rect 4386 11116 4396 11172
rect 4452 11116 6188 11172
rect 6244 11116 6254 11172
rect 14354 11116 14364 11172
rect 14420 11116 14812 11172
rect 14868 11116 14878 11172
rect 15474 11116 15484 11172
rect 15540 11116 22092 11172
rect 22148 11116 22158 11172
rect 22642 11116 22652 11172
rect 22708 11116 23772 11172
rect 23828 11116 23838 11172
rect 25554 11116 25564 11172
rect 25620 11116 26124 11172
rect 26180 11116 28252 11172
rect 28308 11116 28318 11172
rect 34066 11116 34076 11172
rect 34132 11116 34636 11172
rect 34692 11116 35308 11172
rect 35364 11116 40908 11172
rect 40964 11116 40974 11172
rect 41794 11116 41804 11172
rect 41860 11116 42588 11172
rect 42644 11116 42654 11172
rect 44482 11116 44492 11172
rect 44548 11116 50204 11172
rect 50260 11116 50270 11172
rect 50642 11116 50652 11172
rect 50708 11116 51044 11172
rect 54786 11116 54796 11172
rect 54852 11116 54908 11172
rect 54964 11116 54974 11172
rect 23772 11060 23828 11116
rect 3602 11004 3612 11060
rect 3668 11004 4620 11060
rect 4676 11004 8092 11060
rect 8148 11004 8876 11060
rect 8932 11004 17724 11060
rect 17780 11004 17790 11060
rect 22754 11004 22764 11060
rect 22820 11004 23100 11060
rect 23156 11004 23166 11060
rect 23772 11004 30828 11060
rect 30884 11004 30894 11060
rect 36194 11004 36204 11060
rect 36260 11004 45388 11060
rect 45444 11004 45454 11060
rect 46498 11004 46508 11060
rect 46564 11004 47740 11060
rect 47796 11004 47806 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 45388 10948 45444 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 50988 10948 51044 11116
rect 51650 11004 51660 11060
rect 51716 11004 56476 11060
rect 56532 11004 56542 11060
rect 11554 10892 11564 10948
rect 11620 10892 16940 10948
rect 16996 10892 19684 10948
rect 23202 10892 23212 10948
rect 23268 10892 27020 10948
rect 27076 10892 27086 10948
rect 42578 10892 42588 10948
rect 42644 10892 43596 10948
rect 43652 10892 43662 10948
rect 45388 10892 47628 10948
rect 47684 10892 47694 10948
rect 50978 10892 50988 10948
rect 51044 10892 51054 10948
rect 19628 10836 19684 10892
rect 1250 10780 1260 10836
rect 1316 10780 4284 10836
rect 4340 10780 4350 10836
rect 6738 10780 6748 10836
rect 6804 10780 7420 10836
rect 7476 10780 7486 10836
rect 14690 10780 14700 10836
rect 14756 10780 17948 10836
rect 18004 10780 18014 10836
rect 19628 10780 22204 10836
rect 22260 10780 25564 10836
rect 25620 10780 25630 10836
rect 25778 10780 25788 10836
rect 25844 10780 27244 10836
rect 27300 10780 27310 10836
rect 28578 10780 28588 10836
rect 28644 10780 29820 10836
rect 29876 10780 29886 10836
rect 35746 10780 35756 10836
rect 35812 10780 51772 10836
rect 51828 10780 51996 10836
rect 52052 10780 52062 10836
rect 52658 10780 52668 10836
rect 52724 10780 53564 10836
rect 53620 10780 53630 10836
rect 55346 10780 55356 10836
rect 55412 10780 58716 10836
rect 58772 10780 58782 10836
rect 2080 10668 2156 10724
rect 2212 10668 2380 10724
rect 2436 10668 2446 10724
rect 3154 10668 3164 10724
rect 3220 10668 4508 10724
rect 4564 10668 6300 10724
rect 6356 10668 7868 10724
rect 7924 10668 7934 10724
rect 8306 10668 8316 10724
rect 8372 10668 10780 10724
rect 10836 10668 20412 10724
rect 20468 10668 20860 10724
rect 20916 10668 20926 10724
rect 24098 10668 24108 10724
rect 24164 10668 30156 10724
rect 30212 10668 30222 10724
rect 50194 10668 50204 10724
rect 50260 10668 52108 10724
rect 52164 10668 52174 10724
rect 4946 10556 4956 10612
rect 5012 10556 5180 10612
rect 5236 10556 5246 10612
rect 6402 10556 6412 10612
rect 6468 10556 7084 10612
rect 7140 10556 7150 10612
rect 7634 10556 7644 10612
rect 7700 10556 7756 10612
rect 7812 10556 8204 10612
rect 8260 10556 8270 10612
rect 11218 10556 11228 10612
rect 11284 10556 13356 10612
rect 13412 10556 14588 10612
rect 14644 10556 14654 10612
rect 14802 10556 14812 10612
rect 14868 10556 15596 10612
rect 15652 10556 16044 10612
rect 16100 10556 16110 10612
rect 17042 10556 17052 10612
rect 17108 10556 18284 10612
rect 18340 10556 18350 10612
rect 19170 10556 19180 10612
rect 19236 10556 20300 10612
rect 20356 10556 20636 10612
rect 20692 10556 22092 10612
rect 22148 10556 22158 10612
rect 23874 10556 23884 10612
rect 23940 10556 25676 10612
rect 25732 10556 25742 10612
rect 28064 10556 28140 10612
rect 28196 10556 28700 10612
rect 28756 10556 28766 10612
rect 31490 10556 31500 10612
rect 31556 10556 45388 10612
rect 45444 10556 45454 10612
rect 49970 10556 49980 10612
rect 50036 10556 51212 10612
rect 51268 10556 56588 10612
rect 56644 10556 56654 10612
rect 3154 10444 3164 10500
rect 3220 10444 6748 10500
rect 6804 10444 6814 10500
rect 17714 10444 17724 10500
rect 17780 10444 20188 10500
rect 20244 10444 20254 10500
rect 21298 10444 21308 10500
rect 21364 10444 24780 10500
rect 24836 10444 24846 10500
rect 28466 10444 28476 10500
rect 28532 10444 29260 10500
rect 29316 10444 29932 10500
rect 29988 10444 29998 10500
rect 37986 10444 37996 10500
rect 38052 10444 38220 10500
rect 38276 10444 38286 10500
rect 39442 10444 39452 10500
rect 39508 10444 39788 10500
rect 39844 10444 43036 10500
rect 43092 10444 43102 10500
rect 48524 10444 54908 10500
rect 54964 10444 54974 10500
rect 56438 10444 56476 10500
rect 56532 10444 56542 10500
rect 57362 10444 57372 10500
rect 57428 10444 57438 10500
rect 48524 10388 48580 10444
rect 3266 10332 3276 10388
rect 3332 10332 4732 10388
rect 4788 10332 10108 10388
rect 10164 10332 10174 10388
rect 19842 10332 19852 10388
rect 19908 10332 20300 10388
rect 20356 10332 20366 10388
rect 23538 10332 23548 10388
rect 23604 10332 24332 10388
rect 24388 10332 24398 10388
rect 30706 10332 30716 10388
rect 30772 10332 48524 10388
rect 48580 10332 48590 10388
rect 5506 10220 5516 10276
rect 5572 10220 6412 10276
rect 6468 10220 6478 10276
rect 13840 10220 13916 10276
rect 13972 10220 15316 10276
rect 16034 10220 16044 10276
rect 16100 10220 24668 10276
rect 24724 10220 24734 10276
rect 51212 10220 53004 10276
rect 53060 10220 53070 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 15260 10164 15316 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 51212 10164 51268 10220
rect 57372 10164 57428 10444
rect 4844 10108 5404 10164
rect 5460 10108 5470 10164
rect 14028 10108 15148 10164
rect 15260 10108 19068 10164
rect 19124 10108 19134 10164
rect 48626 10108 48636 10164
rect 48692 10108 50876 10164
rect 50932 10108 51268 10164
rect 51426 10108 51436 10164
rect 51492 10108 51548 10164
rect 51604 10108 51614 10164
rect 57260 10108 57428 10164
rect 4844 9940 4900 10108
rect 14028 10052 14084 10108
rect 15092 10052 15148 10108
rect 57260 10052 57316 10108
rect 9762 9996 9772 10052
rect 9828 9996 10556 10052
rect 10612 9996 12684 10052
rect 12740 9996 14084 10052
rect 14242 9996 14252 10052
rect 14308 9996 14924 10052
rect 14980 9996 14990 10052
rect 15092 9996 16492 10052
rect 16548 9996 16558 10052
rect 22754 9996 22764 10052
rect 22820 9996 23324 10052
rect 23380 9996 24220 10052
rect 24276 9996 24286 10052
rect 26114 9996 26124 10052
rect 26180 9996 27132 10052
rect 27188 9996 27198 10052
rect 41234 9996 41244 10052
rect 41300 9996 41916 10052
rect 41972 9996 43596 10052
rect 43652 9996 43662 10052
rect 45042 9996 45052 10052
rect 45108 9996 45500 10052
rect 45556 9996 45566 10052
rect 48850 9996 48860 10052
rect 48916 9996 49084 10052
rect 49140 9996 49150 10052
rect 49522 9996 49532 10052
rect 49588 9996 51324 10052
rect 51380 9996 51390 10052
rect 53778 9996 53788 10052
rect 53844 9996 56924 10052
rect 56980 9996 56990 10052
rect 57250 9996 57260 10052
rect 57316 9996 57326 10052
rect 2370 9884 2380 9940
rect 2436 9884 3500 9940
rect 3556 9884 4060 9940
rect 4116 9884 4900 9940
rect 6514 9884 6524 9940
rect 6580 9884 8092 9940
rect 8148 9884 8158 9940
rect 11890 9884 11900 9940
rect 11956 9884 12796 9940
rect 12852 9884 14140 9940
rect 14196 9884 14206 9940
rect 15894 9884 15932 9940
rect 15988 9884 15998 9940
rect 19954 9884 19964 9940
rect 20020 9884 20748 9940
rect 20804 9884 20814 9940
rect 23090 9884 23100 9940
rect 23156 9884 27356 9940
rect 27412 9884 28364 9940
rect 28420 9884 29484 9940
rect 29540 9884 29550 9940
rect 43474 9884 43484 9940
rect 43540 9884 45612 9940
rect 45668 9884 45678 9940
rect 47954 9884 47964 9940
rect 48020 9884 48300 9940
rect 48356 9884 49420 9940
rect 49476 9884 49486 9940
rect 51874 9884 51884 9940
rect 51940 9884 52444 9940
rect 52500 9884 52510 9940
rect 55570 9884 55580 9940
rect 55636 9884 56252 9940
rect 56308 9884 56318 9940
rect 58034 9884 58044 9940
rect 58100 9884 59164 9940
rect 59220 9884 59230 9940
rect 4946 9772 4956 9828
rect 5012 9772 6188 9828
rect 6244 9772 7308 9828
rect 7364 9772 7374 9828
rect 9650 9772 9660 9828
rect 9716 9772 11228 9828
rect 11284 9772 11294 9828
rect 14018 9772 14028 9828
rect 14084 9772 14364 9828
rect 14420 9772 14700 9828
rect 14756 9772 14924 9828
rect 14980 9772 14990 9828
rect 15250 9772 15260 9828
rect 15316 9772 16044 9828
rect 16100 9772 18956 9828
rect 19012 9772 21756 9828
rect 21812 9772 22540 9828
rect 22596 9772 22606 9828
rect 23762 9772 23772 9828
rect 23828 9772 25900 9828
rect 25956 9772 26348 9828
rect 26404 9772 27020 9828
rect 27076 9772 27086 9828
rect 36082 9772 36092 9828
rect 36148 9772 38668 9828
rect 38724 9772 38734 9828
rect 43474 9772 43484 9828
rect 43540 9772 54684 9828
rect 54740 9772 54750 9828
rect 3938 9660 3948 9716
rect 4004 9660 4620 9716
rect 4676 9660 4686 9716
rect 5394 9660 5404 9716
rect 5460 9660 16268 9716
rect 16324 9660 16334 9716
rect 36642 9660 36652 9716
rect 36708 9660 45948 9716
rect 46004 9660 46014 9716
rect 48066 9660 48076 9716
rect 48132 9660 52332 9716
rect 52388 9660 52892 9716
rect 52948 9660 52958 9716
rect 3714 9548 3724 9604
rect 3780 9548 10668 9604
rect 10724 9548 10734 9604
rect 16146 9548 16156 9604
rect 16212 9548 19964 9604
rect 20020 9548 20030 9604
rect 40338 9548 40348 9604
rect 40404 9548 41020 9604
rect 41076 9548 42140 9604
rect 42196 9548 42206 9604
rect 44034 9548 44044 9604
rect 44100 9548 44716 9604
rect 44772 9548 45276 9604
rect 45332 9548 45342 9604
rect 47170 9548 47180 9604
rect 47236 9548 52108 9604
rect 52164 9548 52174 9604
rect 2706 9436 2716 9492
rect 2772 9436 3164 9492
rect 3220 9436 6300 9492
rect 6356 9436 6636 9492
rect 6692 9436 14812 9492
rect 14868 9436 15148 9492
rect 15810 9436 15820 9492
rect 15876 9436 16268 9492
rect 16324 9436 16334 9492
rect 19618 9436 19628 9492
rect 19684 9436 19694 9492
rect 21308 9436 22316 9492
rect 22372 9436 23100 9492
rect 23156 9436 23166 9492
rect 28690 9436 28700 9492
rect 28756 9436 41132 9492
rect 41188 9436 41198 9492
rect 51874 9436 51884 9492
rect 51940 9436 52556 9492
rect 52612 9436 54684 9492
rect 54740 9436 54750 9492
rect 15092 9380 15148 9436
rect 19628 9380 19684 9436
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 3714 9324 3724 9380
rect 3780 9324 7196 9380
rect 7252 9324 9548 9380
rect 9604 9324 9614 9380
rect 11676 9324 14812 9380
rect 14868 9324 14878 9380
rect 15092 9324 15932 9380
rect 15988 9324 15998 9380
rect 16594 9324 16604 9380
rect 16660 9324 19684 9380
rect 11676 9268 11732 9324
rect 19628 9268 19684 9324
rect 8194 9212 8204 9268
rect 8260 9212 10220 9268
rect 10276 9212 10286 9268
rect 11638 9212 11676 9268
rect 11732 9212 11742 9268
rect 13654 9212 13692 9268
rect 13748 9212 13758 9268
rect 13916 9212 15148 9268
rect 15204 9212 15214 9268
rect 16118 9212 16156 9268
rect 16212 9212 16222 9268
rect 17042 9212 17052 9268
rect 17108 9212 18620 9268
rect 18676 9212 18686 9268
rect 19628 9212 19964 9268
rect 20020 9212 20030 9268
rect 13916 9156 13972 9212
rect 1922 9100 1932 9156
rect 1988 9100 3948 9156
rect 4004 9100 6524 9156
rect 6580 9100 7700 9156
rect 9762 9100 9772 9156
rect 9828 9100 13972 9156
rect 14914 9100 14924 9156
rect 14980 9100 15820 9156
rect 15876 9100 15886 9156
rect 7644 9044 7700 9100
rect 14924 9044 14980 9100
rect 21308 9044 21364 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 21522 9324 21532 9380
rect 21588 9324 23996 9380
rect 24052 9324 24062 9380
rect 33954 9324 33964 9380
rect 34020 9324 41804 9380
rect 41860 9324 41870 9380
rect 55458 9324 55468 9380
rect 55524 9324 56700 9380
rect 56756 9324 56766 9380
rect 21858 9212 21868 9268
rect 21924 9212 22540 9268
rect 22596 9212 22606 9268
rect 24210 9212 24220 9268
rect 24276 9212 28364 9268
rect 28420 9212 28430 9268
rect 48262 9212 48300 9268
rect 48356 9212 51100 9268
rect 51156 9212 51166 9268
rect 51874 9212 51884 9268
rect 51940 9212 52556 9268
rect 52612 9212 52622 9268
rect 53666 9212 53676 9268
rect 53732 9212 54012 9268
rect 54068 9212 54078 9268
rect 54338 9212 54348 9268
rect 54404 9212 55916 9268
rect 55972 9212 56140 9268
rect 56196 9212 56206 9268
rect 22978 9100 22988 9156
rect 23044 9100 23212 9156
rect 23268 9100 24556 9156
rect 24612 9100 24622 9156
rect 40450 9100 40460 9156
rect 40516 9100 42588 9156
rect 42644 9100 45276 9156
rect 45332 9100 45342 9156
rect 2818 8988 2828 9044
rect 2884 8988 3948 9044
rect 4004 8988 5068 9044
rect 5124 8988 5134 9044
rect 6402 8988 6412 9044
rect 6468 8988 7420 9044
rect 7476 8988 7486 9044
rect 7644 8988 12236 9044
rect 12292 8988 12302 9044
rect 12562 8988 12572 9044
rect 12628 8988 13916 9044
rect 13972 8988 14980 9044
rect 15250 8988 15260 9044
rect 15316 8988 21364 9044
rect 24882 8988 24892 9044
rect 24948 8988 25788 9044
rect 25844 8988 25854 9044
rect 26002 8988 26012 9044
rect 26068 8988 26460 9044
rect 26516 8988 26908 9044
rect 26964 8988 27468 9044
rect 27524 8988 27534 9044
rect 34962 8988 34972 9044
rect 35028 8988 37772 9044
rect 37828 8988 37838 9044
rect 41346 8988 41356 9044
rect 41412 8988 44828 9044
rect 44884 8988 44894 9044
rect 51062 8988 51100 9044
rect 51156 8988 51166 9044
rect 5590 8876 5628 8932
rect 5684 8876 5694 8932
rect 7746 8876 7756 8932
rect 7812 8876 8540 8932
rect 8596 8876 8876 8932
rect 8932 8876 8942 8932
rect 14774 8876 14812 8932
rect 14868 8876 14878 8932
rect 18610 8876 18620 8932
rect 18676 8876 19180 8932
rect 19236 8876 19628 8932
rect 19684 8876 19694 8932
rect 20738 8876 20748 8932
rect 20804 8876 22428 8932
rect 22484 8876 22494 8932
rect 36866 8876 36876 8932
rect 36932 8876 37436 8932
rect 37492 8876 37502 8932
rect 50306 8876 50316 8932
rect 50372 8876 50428 8932
rect 50484 8876 51548 8932
rect 51604 8876 51614 8932
rect 5506 8764 5516 8820
rect 5572 8764 9100 8820
rect 9156 8764 9436 8820
rect 9492 8764 9502 8820
rect 19030 8764 19068 8820
rect 19124 8764 19134 8820
rect 45602 8764 45612 8820
rect 45668 8764 46396 8820
rect 46452 8764 53788 8820
rect 53844 8764 53854 8820
rect 56914 8764 56924 8820
rect 56980 8764 57260 8820
rect 57316 8764 57326 8820
rect 44706 8652 44716 8708
rect 44772 8652 52332 8708
rect 52388 8652 53228 8708
rect 53284 8652 53294 8708
rect 56130 8652 56140 8708
rect 56196 8652 57484 8708
rect 57540 8652 57550 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 16146 8540 16156 8596
rect 16212 8540 16492 8596
rect 16548 8540 18956 8596
rect 19012 8540 19740 8596
rect 19796 8540 19806 8596
rect 20402 8540 20412 8596
rect 20468 8540 21980 8596
rect 22036 8540 22988 8596
rect 23044 8540 23054 8596
rect 38612 8540 39116 8596
rect 39172 8540 57708 8596
rect 57764 8540 57774 8596
rect 4498 8428 4508 8484
rect 4564 8428 4956 8484
rect 5012 8428 5022 8484
rect 12226 8428 12236 8484
rect 12292 8428 16828 8484
rect 16884 8428 17388 8484
rect 17444 8428 17454 8484
rect 17602 8428 17612 8484
rect 17668 8428 17948 8484
rect 18004 8428 18508 8484
rect 18564 8428 19516 8484
rect 19572 8428 22764 8484
rect 22820 8428 22830 8484
rect 38612 8372 38668 8540
rect 40898 8428 40908 8484
rect 40964 8428 41356 8484
rect 41412 8428 41422 8484
rect 50866 8428 50876 8484
rect 50932 8428 51212 8484
rect 51268 8428 52220 8484
rect 52276 8428 52286 8484
rect 8978 8316 8988 8372
rect 9044 8316 9884 8372
rect 9940 8316 10332 8372
rect 10388 8316 10398 8372
rect 11666 8316 11676 8372
rect 11732 8316 13580 8372
rect 13636 8316 13860 8372
rect 15810 8316 15820 8372
rect 15876 8316 16044 8372
rect 16100 8316 16110 8372
rect 19282 8316 19292 8372
rect 19348 8316 19740 8372
rect 19796 8316 19806 8372
rect 19954 8316 19964 8372
rect 20020 8316 20300 8372
rect 20356 8316 20366 8372
rect 20850 8316 20860 8372
rect 20916 8316 22092 8372
rect 22148 8316 25452 8372
rect 25508 8316 25518 8372
rect 32722 8316 32732 8372
rect 32788 8316 38668 8372
rect 43250 8316 43260 8372
rect 43316 8316 43820 8372
rect 43876 8316 44156 8372
rect 44212 8316 44222 8372
rect 44818 8316 44828 8372
rect 44884 8316 52892 8372
rect 52948 8316 53340 8372
rect 53396 8316 53406 8372
rect 54674 8316 54684 8372
rect 54740 8316 55132 8372
rect 55188 8316 56252 8372
rect 56308 8316 56588 8372
rect 56644 8316 56654 8372
rect 7522 8204 7532 8260
rect 7588 8204 8428 8260
rect 8484 8204 8764 8260
rect 8820 8204 8830 8260
rect 9986 8204 9996 8260
rect 10052 8204 10780 8260
rect 10836 8204 12348 8260
rect 12404 8204 12414 8260
rect 8978 8092 8988 8148
rect 9044 8092 11788 8148
rect 11844 8092 13580 8148
rect 13636 8092 13646 8148
rect 2482 7980 2492 8036
rect 2548 7980 3612 8036
rect 3668 7980 3678 8036
rect 6412 7980 8204 8036
rect 8260 7980 8270 8036
rect 6412 7924 6468 7980
rect 13804 7924 13860 8316
rect 17826 8204 17836 8260
rect 17892 8204 21532 8260
rect 21588 8204 21598 8260
rect 29362 8204 29372 8260
rect 29428 8204 38332 8260
rect 38388 8204 38398 8260
rect 39554 8204 39564 8260
rect 39620 8204 45948 8260
rect 46004 8204 46014 8260
rect 49942 8204 49980 8260
rect 50036 8204 50046 8260
rect 51202 8204 51212 8260
rect 51268 8204 51436 8260
rect 51492 8204 53452 8260
rect 53508 8204 54236 8260
rect 54292 8204 54302 8260
rect 49980 8148 50036 8204
rect 59200 8148 59800 8176
rect 19628 8092 22036 8148
rect 22194 8092 22204 8148
rect 22260 8092 23100 8148
rect 23156 8092 23166 8148
rect 25554 8092 25564 8148
rect 25620 8092 26124 8148
rect 26180 8092 26190 8148
rect 33394 8092 33404 8148
rect 33460 8092 41804 8148
rect 41860 8092 41870 8148
rect 42690 8092 42700 8148
rect 42756 8092 50036 8148
rect 51650 8092 51660 8148
rect 51716 8092 52108 8148
rect 52164 8092 52174 8148
rect 55346 8092 55356 8148
rect 55412 8092 59800 8148
rect 14018 7980 14028 8036
rect 14084 7980 15820 8036
rect 15876 7980 15886 8036
rect 2370 7868 2380 7924
rect 2436 7868 6468 7924
rect 7410 7868 7420 7924
rect 7476 7868 11676 7924
rect 11732 7868 11742 7924
rect 13794 7868 13804 7924
rect 13860 7868 13870 7924
rect 19628 7812 19684 8092
rect 21980 8036 22036 8092
rect 59200 8064 59800 8092
rect 21980 7980 22540 8036
rect 22596 7980 25340 8036
rect 25396 7980 25406 8036
rect 26674 7980 26684 8036
rect 26740 7980 27244 8036
rect 27300 7980 27310 8036
rect 29596 7980 38668 8036
rect 43922 7980 43932 8036
rect 43988 7980 49420 8036
rect 49476 7980 49486 8036
rect 50372 7980 51044 8036
rect 52770 7980 52780 8036
rect 52836 7980 53116 8036
rect 53172 7980 54236 8036
rect 54292 7980 54796 8036
rect 54852 7980 54862 8036
rect 57586 7980 57596 8036
rect 57652 7980 58828 8036
rect 58884 7980 58894 8036
rect 29596 7924 29652 7980
rect 26114 7868 26124 7924
rect 26180 7868 26908 7924
rect 26964 7868 27692 7924
rect 27748 7868 29652 7924
rect 38612 7924 38668 7980
rect 38612 7868 45164 7924
rect 45220 7868 45230 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50372 7812 50428 7980
rect 50988 7924 51044 7980
rect 50988 7868 59612 7924
rect 59668 7868 59678 7924
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 6066 7756 6076 7812
rect 6132 7756 7980 7812
rect 8036 7756 8316 7812
rect 8372 7756 8382 7812
rect 8530 7756 8540 7812
rect 8596 7756 10220 7812
rect 10276 7756 19684 7812
rect 37202 7756 37212 7812
rect 37268 7756 39564 7812
rect 39620 7756 39630 7812
rect 41906 7756 41916 7812
rect 41972 7756 50428 7812
rect 53106 7756 53116 7812
rect 53172 7756 53788 7812
rect 53844 7756 53854 7812
rect 2930 7644 2940 7700
rect 2996 7644 3388 7700
rect 3444 7644 3454 7700
rect 6738 7644 6748 7700
rect 6804 7644 7308 7700
rect 7364 7644 7374 7700
rect 7746 7644 7756 7700
rect 7812 7644 11788 7700
rect 11844 7644 12012 7700
rect 12068 7644 12078 7700
rect 12450 7644 12460 7700
rect 12516 7644 14252 7700
rect 14308 7644 14318 7700
rect 17826 7644 17836 7700
rect 17892 7644 18620 7700
rect 18676 7644 18686 7700
rect 19506 7644 19516 7700
rect 19572 7644 19852 7700
rect 19908 7644 19918 7700
rect 20290 7644 20300 7700
rect 20356 7644 21084 7700
rect 21140 7644 21150 7700
rect 23874 7644 23884 7700
rect 23940 7644 24444 7700
rect 24500 7644 24510 7700
rect 33618 7644 33628 7700
rect 33684 7644 37996 7700
rect 38052 7644 38668 7700
rect 38724 7644 38734 7700
rect 46498 7644 46508 7700
rect 46564 7644 47292 7700
rect 47348 7644 47358 7700
rect 47954 7644 47964 7700
rect 48020 7644 49532 7700
rect 49588 7644 49598 7700
rect 50306 7644 50316 7700
rect 50372 7644 51772 7700
rect 51828 7644 52108 7700
rect 52164 7644 52174 7700
rect 53554 7644 53564 7700
rect 53620 7644 56588 7700
rect 56644 7644 57484 7700
rect 57540 7644 57550 7700
rect 7756 7588 7812 7644
rect 14252 7588 14308 7644
rect 2034 7532 2044 7588
rect 2100 7532 3164 7588
rect 3220 7532 4620 7588
rect 4676 7532 4686 7588
rect 5394 7532 5404 7588
rect 5460 7532 6636 7588
rect 6692 7532 7812 7588
rect 10882 7532 10892 7588
rect 10948 7532 12124 7588
rect 12180 7532 12684 7588
rect 12740 7532 12750 7588
rect 14252 7532 22876 7588
rect 22932 7532 22942 7588
rect 46946 7532 46956 7588
rect 47012 7532 50092 7588
rect 50148 7532 55244 7588
rect 55300 7532 55310 7588
rect 5506 7420 5516 7476
rect 5572 7420 6748 7476
rect 6804 7420 7084 7476
rect 7140 7420 7150 7476
rect 14578 7420 14588 7476
rect 14644 7420 15036 7476
rect 15092 7420 15102 7476
rect 16370 7420 16380 7476
rect 16436 7420 17500 7476
rect 17556 7420 17566 7476
rect 18162 7420 18172 7476
rect 18228 7420 19292 7476
rect 19348 7420 21868 7476
rect 21924 7420 22204 7476
rect 22260 7420 22270 7476
rect 24882 7420 24892 7476
rect 24948 7420 25452 7476
rect 25508 7420 25518 7476
rect 25666 7420 25676 7476
rect 25732 7420 26460 7476
rect 26516 7420 26526 7476
rect 46610 7420 46620 7476
rect 46676 7420 50876 7476
rect 50932 7420 50942 7476
rect 3826 7308 3836 7364
rect 3892 7308 8652 7364
rect 8708 7308 9660 7364
rect 9716 7308 9726 7364
rect 13682 7308 13692 7364
rect 13748 7308 18844 7364
rect 18900 7308 22764 7364
rect 22820 7308 23548 7364
rect 23604 7308 23614 7364
rect 38322 7308 38332 7364
rect 38388 7308 38780 7364
rect 38836 7308 38846 7364
rect 40002 7308 40012 7364
rect 40068 7308 42588 7364
rect 42644 7308 42654 7364
rect 49858 7308 49868 7364
rect 49924 7308 50764 7364
rect 50820 7308 50830 7364
rect 56690 7308 56700 7364
rect 56756 7308 57820 7364
rect 57876 7308 57886 7364
rect 40012 7252 40068 7308
rect 4162 7196 4172 7252
rect 4228 7196 4396 7252
rect 4452 7196 10556 7252
rect 10612 7196 10622 7252
rect 12338 7196 12348 7252
rect 12404 7196 16380 7252
rect 16436 7196 16446 7252
rect 20178 7196 20188 7252
rect 20244 7196 20860 7252
rect 20916 7196 23436 7252
rect 23492 7196 23772 7252
rect 23828 7196 23838 7252
rect 26908 7196 40068 7252
rect 49410 7196 49420 7252
rect 49476 7196 55692 7252
rect 55748 7196 55758 7252
rect 26908 7140 26964 7196
rect 10210 7084 10220 7140
rect 10276 7084 11564 7140
rect 11620 7084 18732 7140
rect 18788 7084 18798 7140
rect 19618 7084 19628 7140
rect 19684 7084 22316 7140
rect 22372 7084 22382 7140
rect 26898 7084 26908 7140
rect 26964 7084 26974 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 15810 6972 15820 7028
rect 15876 6972 23884 7028
rect 23940 6972 23950 7028
rect 18732 6916 18788 6972
rect 1922 6860 1932 6916
rect 1988 6860 2268 6916
rect 2324 6860 3836 6916
rect 3892 6860 6076 6916
rect 6132 6860 6142 6916
rect 9202 6860 9212 6916
rect 9268 6860 15036 6916
rect 15092 6860 18396 6916
rect 18452 6860 18462 6916
rect 18722 6860 18732 6916
rect 18788 6860 18798 6916
rect 23538 6860 23548 6916
rect 23604 6860 25228 6916
rect 25284 6860 25788 6916
rect 25844 6860 25854 6916
rect 43362 6860 43372 6916
rect 43428 6860 48188 6916
rect 48244 6860 48254 6916
rect 58034 6860 58044 6916
rect 58100 6860 58110 6916
rect 58044 6804 58100 6860
rect 5170 6748 5180 6804
rect 5236 6748 5740 6804
rect 5796 6748 5806 6804
rect 7634 6748 7644 6804
rect 7700 6748 7710 6804
rect 10658 6748 10668 6804
rect 10724 6748 11004 6804
rect 11060 6748 11340 6804
rect 11396 6748 11406 6804
rect 11788 6748 12236 6804
rect 12292 6748 16716 6804
rect 16772 6748 16782 6804
rect 17238 6748 17276 6804
rect 17332 6748 17342 6804
rect 22306 6748 22316 6804
rect 22372 6748 22876 6804
rect 22932 6748 22942 6804
rect 24322 6748 24332 6804
rect 24388 6748 28028 6804
rect 28084 6748 28094 6804
rect 29362 6748 29372 6804
rect 29428 6748 43708 6804
rect 43764 6748 43774 6804
rect 50866 6748 50876 6804
rect 50932 6748 52556 6804
rect 52612 6748 52622 6804
rect 54450 6748 54460 6804
rect 54516 6748 55580 6804
rect 55636 6748 58100 6804
rect 7644 6692 7700 6748
rect 11788 6692 11844 6748
rect 1138 6636 1148 6692
rect 1204 6636 2604 6692
rect 2660 6636 3164 6692
rect 3220 6636 3230 6692
rect 7074 6636 7084 6692
rect 7140 6636 7700 6692
rect 10322 6636 10332 6692
rect 10388 6636 11844 6692
rect 12114 6636 12124 6692
rect 12180 6636 13020 6692
rect 13076 6636 13580 6692
rect 13636 6636 13646 6692
rect 15698 6636 15708 6692
rect 15764 6636 16380 6692
rect 16436 6636 16446 6692
rect 16930 6636 16940 6692
rect 16996 6636 19516 6692
rect 19572 6636 22092 6692
rect 22148 6636 22540 6692
rect 22596 6636 23772 6692
rect 23828 6636 23838 6692
rect 37762 6636 37772 6692
rect 37828 6636 38220 6692
rect 38276 6636 38286 6692
rect 38434 6636 38444 6692
rect 38500 6636 45948 6692
rect 46004 6636 47068 6692
rect 47124 6636 47134 6692
rect 49074 6636 49084 6692
rect 49140 6636 50428 6692
rect 51202 6636 51212 6692
rect 51268 6636 51884 6692
rect 51940 6636 53564 6692
rect 53620 6636 53630 6692
rect 54114 6636 54124 6692
rect 54180 6636 54908 6692
rect 54964 6636 55804 6692
rect 55860 6636 55870 6692
rect 56690 6636 56700 6692
rect 56756 6636 57372 6692
rect 57428 6636 57438 6692
rect 4498 6524 4508 6580
rect 4564 6524 5516 6580
rect 5572 6524 8092 6580
rect 8148 6524 8158 6580
rect 9762 6524 9772 6580
rect 9828 6524 13692 6580
rect 13748 6524 14028 6580
rect 14084 6524 14094 6580
rect 14242 6524 14252 6580
rect 14308 6524 15148 6580
rect 15204 6524 15214 6580
rect 18050 6524 18060 6580
rect 18116 6524 18956 6580
rect 19012 6524 20076 6580
rect 20132 6524 20142 6580
rect 22726 6524 22764 6580
rect 22820 6524 22830 6580
rect 23426 6524 23436 6580
rect 23492 6524 23884 6580
rect 23940 6524 23950 6580
rect 24546 6524 24556 6580
rect 24612 6524 26124 6580
rect 26180 6524 26190 6580
rect 44482 6524 44492 6580
rect 44548 6524 47740 6580
rect 47796 6524 47806 6580
rect 48514 6524 48524 6580
rect 48580 6524 49420 6580
rect 49476 6524 49868 6580
rect 49924 6524 49934 6580
rect 23884 6468 23940 6524
rect 50372 6468 50428 6636
rect 52994 6524 53004 6580
rect 53060 6524 54236 6580
rect 54292 6524 54460 6580
rect 54516 6524 55356 6580
rect 55412 6524 55422 6580
rect 4946 6412 4956 6468
rect 5012 6412 8988 6468
rect 9044 6412 10332 6468
rect 10388 6412 10398 6468
rect 10658 6412 10668 6468
rect 10724 6412 11452 6468
rect 11508 6412 16604 6468
rect 16660 6412 20300 6468
rect 20356 6412 20366 6468
rect 23884 6412 26572 6468
rect 26628 6412 26638 6468
rect 40562 6412 40572 6468
rect 40628 6412 41356 6468
rect 41412 6412 44604 6468
rect 44660 6412 44670 6468
rect 50372 6412 52108 6468
rect 52164 6412 55020 6468
rect 55076 6412 57596 6468
rect 57652 6412 57820 6468
rect 57876 6412 57886 6468
rect 10668 6356 10724 6412
rect 3714 6300 3724 6356
rect 3780 6300 6524 6356
rect 6580 6300 10108 6356
rect 10164 6300 10724 6356
rect 12898 6300 12908 6356
rect 12964 6300 13244 6356
rect 13300 6300 13310 6356
rect 18050 6300 18060 6356
rect 18116 6300 18284 6356
rect 18340 6300 18350 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 2706 6188 2716 6244
rect 2772 6188 5628 6244
rect 5684 6188 5740 6244
rect 5796 6188 5806 6244
rect 8082 6188 8092 6244
rect 8148 6188 10780 6244
rect 10836 6188 10846 6244
rect 14018 6188 14028 6244
rect 14084 6188 14924 6244
rect 14980 6188 15708 6244
rect 15764 6188 15774 6244
rect 3910 6076 3948 6132
rect 4004 6076 4014 6132
rect 4498 6076 4508 6132
rect 4564 6076 5292 6132
rect 5348 6076 10220 6132
rect 10276 6076 10286 6132
rect 15138 6076 15148 6132
rect 15204 6076 15484 6132
rect 15540 6076 15550 6132
rect 15810 6076 15820 6132
rect 15876 6076 19628 6132
rect 19684 6076 19694 6132
rect 20626 6076 20636 6132
rect 20692 6076 21420 6132
rect 21476 6076 21486 6132
rect 30370 6076 30380 6132
rect 30436 6076 36316 6132
rect 36372 6076 37772 6132
rect 37828 6076 37838 6132
rect 47618 6076 47628 6132
rect 47684 6076 48524 6132
rect 48580 6076 48972 6132
rect 49028 6076 49038 6132
rect 49858 6076 49868 6132
rect 49924 6076 54684 6132
rect 54740 6076 54750 6132
rect 56018 6076 56028 6132
rect 56084 6076 56476 6132
rect 56532 6076 56542 6132
rect 6402 5964 6412 6020
rect 6468 5964 6636 6020
rect 6692 5964 13132 6020
rect 13188 5964 21756 6020
rect 21812 5964 22540 6020
rect 22596 5964 28476 6020
rect 28532 5964 28542 6020
rect 35074 5964 35084 6020
rect 35140 5964 49980 6020
rect 50036 5964 50046 6020
rect 13234 5852 13244 5908
rect 13300 5852 17836 5908
rect 17892 5852 17902 5908
rect 40786 5852 40796 5908
rect 40852 5852 41468 5908
rect 41524 5852 41534 5908
rect 3490 5740 3500 5796
rect 3556 5740 7084 5796
rect 7140 5740 7150 5796
rect 7634 5740 7644 5796
rect 7700 5740 7868 5796
rect 7924 5740 8428 5796
rect 8484 5740 9660 5796
rect 9716 5740 9726 5796
rect 18274 5740 18284 5796
rect 18340 5740 19068 5796
rect 19124 5740 21644 5796
rect 21700 5740 21710 5796
rect 33506 5740 33516 5796
rect 33572 5740 41356 5796
rect 41412 5740 42028 5796
rect 42084 5740 42094 5796
rect 48178 5740 48188 5796
rect 48244 5740 55916 5796
rect 55972 5740 55982 5796
rect 8194 5628 8204 5684
rect 8260 5628 15820 5684
rect 15876 5628 15886 5684
rect 40226 5628 40236 5684
rect 40292 5628 49084 5684
rect 49140 5628 57148 5684
rect 57204 5628 58380 5684
rect 58436 5628 58446 5684
rect 9986 5516 9996 5572
rect 10052 5516 12460 5572
rect 12516 5516 12908 5572
rect 12964 5516 12974 5572
rect 14242 5516 14252 5572
rect 14308 5516 19628 5572
rect 19684 5516 24332 5572
rect 24388 5516 24398 5572
rect 200 5460 800 5488
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 200 5404 1932 5460
rect 1988 5404 1998 5460
rect 14130 5404 14140 5460
rect 14196 5404 22092 5460
rect 22148 5404 22158 5460
rect 44706 5404 44716 5460
rect 44772 5404 45388 5460
rect 45444 5404 45454 5460
rect 47730 5404 47740 5460
rect 47796 5404 49868 5460
rect 49924 5404 49934 5460
rect 200 5376 800 5404
rect 1362 5292 1372 5348
rect 1428 5292 6188 5348
rect 6244 5292 7308 5348
rect 7364 5292 7374 5348
rect 12338 5292 12348 5348
rect 12404 5292 16604 5348
rect 16660 5292 16670 5348
rect 16930 5292 16940 5348
rect 16996 5292 18060 5348
rect 18116 5292 20020 5348
rect 19964 5236 20020 5292
rect 26852 5292 41916 5348
rect 41972 5292 41982 5348
rect 45388 5292 45612 5348
rect 45668 5292 45678 5348
rect 47282 5292 47292 5348
rect 47348 5292 52444 5348
rect 52500 5292 53340 5348
rect 53396 5292 53788 5348
rect 53844 5292 54572 5348
rect 54628 5292 54638 5348
rect 26852 5236 26908 5292
rect 2034 5180 2044 5236
rect 2100 5180 2156 5236
rect 2212 5180 2222 5236
rect 3938 5180 3948 5236
rect 4004 5180 4508 5236
rect 4564 5180 4574 5236
rect 4946 5180 4956 5236
rect 5012 5180 5516 5236
rect 5572 5180 5582 5236
rect 5842 5180 5852 5236
rect 5908 5180 9492 5236
rect 9622 5180 9660 5236
rect 9716 5180 9726 5236
rect 10518 5180 10556 5236
rect 10612 5180 10622 5236
rect 11526 5180 11564 5236
rect 11620 5180 11630 5236
rect 11890 5180 11900 5236
rect 11956 5180 14812 5236
rect 14868 5180 14878 5236
rect 15810 5180 15820 5236
rect 15876 5180 16828 5236
rect 16884 5180 16894 5236
rect 19954 5180 19964 5236
rect 20020 5180 20580 5236
rect 21858 5180 21868 5236
rect 21924 5180 22988 5236
rect 23044 5180 26908 5236
rect 28802 5180 28812 5236
rect 28868 5180 31052 5236
rect 31108 5180 31118 5236
rect 32386 5180 32396 5236
rect 32452 5180 36428 5236
rect 36484 5180 37996 5236
rect 38052 5180 38062 5236
rect 4508 5124 4564 5180
rect 9436 5124 9492 5180
rect 20524 5124 20580 5180
rect 2146 5068 2156 5124
rect 2212 5068 2604 5124
rect 2660 5068 2670 5124
rect 4508 5068 5964 5124
rect 6020 5068 6030 5124
rect 6850 5068 6860 5124
rect 6916 5068 8764 5124
rect 8820 5068 8830 5124
rect 9436 5068 11340 5124
rect 11396 5068 11406 5124
rect 19282 5068 19292 5124
rect 19348 5068 20300 5124
rect 20356 5068 20366 5124
rect 20524 5068 27356 5124
rect 27412 5068 27422 5124
rect 28812 5012 28868 5180
rect 33618 5068 33628 5124
rect 33684 5068 33852 5124
rect 33908 5068 34636 5124
rect 34692 5068 34702 5124
rect 36866 5068 36876 5124
rect 36932 5068 37436 5124
rect 37492 5068 40796 5124
rect 40852 5068 40862 5124
rect 45388 5012 45444 5292
rect 49970 5180 49980 5236
rect 50036 5180 56700 5236
rect 56756 5180 56766 5236
rect 45714 5068 45724 5124
rect 45780 5068 52444 5124
rect 52500 5068 52510 5124
rect 7858 4956 7868 5012
rect 7924 4956 10892 5012
rect 10948 4956 10958 5012
rect 16706 4956 16716 5012
rect 16772 4956 23436 5012
rect 23492 4956 23502 5012
rect 23762 4956 23772 5012
rect 23828 4956 24108 5012
rect 24164 4956 24668 5012
rect 24724 4956 24892 5012
rect 24948 4956 24958 5012
rect 28354 4956 28364 5012
rect 28420 4956 28868 5012
rect 43810 4956 43820 5012
rect 43876 4956 45444 5012
rect 45602 4956 45612 5012
rect 45668 4956 46732 5012
rect 46788 4956 46798 5012
rect 56242 4956 56252 5012
rect 56308 4956 58604 5012
rect 58660 4956 58670 5012
rect 45388 4900 45444 4956
rect 7074 4844 7084 4900
rect 7140 4844 25228 4900
rect 25284 4844 25294 4900
rect 45388 4844 47740 4900
rect 47796 4844 47806 4900
rect 48514 4844 48524 4900
rect 48580 4844 51436 4900
rect 51492 4844 58044 4900
rect 58100 4844 58110 4900
rect 14578 4732 14588 4788
rect 14644 4732 15372 4788
rect 15428 4732 15438 4788
rect 15586 4732 15596 4788
rect 15652 4732 17276 4788
rect 17332 4732 17342 4788
rect 41906 4732 41916 4788
rect 41972 4732 43708 4788
rect 43764 4732 47516 4788
rect 47572 4732 47582 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 4946 4620 4956 4676
rect 5012 4620 5404 4676
rect 5460 4620 5470 4676
rect 9090 4620 9100 4676
rect 9156 4620 19684 4676
rect 20178 4620 20188 4676
rect 20244 4620 49644 4676
rect 49700 4620 49710 4676
rect 19628 4564 19684 4620
rect 4610 4508 4620 4564
rect 4676 4508 6636 4564
rect 6692 4508 6702 4564
rect 8642 4508 8652 4564
rect 8708 4508 10108 4564
rect 10164 4508 10174 4564
rect 10658 4508 10668 4564
rect 10724 4508 11228 4564
rect 11284 4508 13020 4564
rect 13076 4508 14140 4564
rect 14196 4508 14206 4564
rect 14578 4508 14588 4564
rect 14644 4508 15148 4564
rect 15204 4508 15214 4564
rect 15372 4508 15820 4564
rect 15876 4508 15886 4564
rect 16482 4508 16492 4564
rect 16548 4508 16940 4564
rect 16996 4508 18172 4564
rect 18228 4508 18238 4564
rect 19628 4508 28140 4564
rect 28196 4508 28206 4564
rect 40114 4508 40124 4564
rect 40180 4508 40460 4564
rect 40516 4508 45948 4564
rect 46004 4508 46014 4564
rect 48066 4508 48076 4564
rect 48132 4508 49980 4564
rect 50036 4508 52332 4564
rect 52388 4508 52398 4564
rect 15372 4452 15428 4508
rect 1026 4396 1036 4452
rect 1092 4396 2716 4452
rect 2772 4396 3612 4452
rect 3668 4396 3678 4452
rect 13794 4396 13804 4452
rect 13860 4396 15428 4452
rect 17714 4396 17724 4452
rect 17780 4396 22316 4452
rect 22372 4396 22382 4452
rect 56130 4396 56140 4452
rect 56196 4396 57484 4452
rect 57540 4396 57550 4452
rect 5058 4284 5068 4340
rect 5124 4284 8204 4340
rect 8260 4284 12684 4340
rect 12740 4284 16492 4340
rect 16548 4284 16558 4340
rect 28354 4284 28364 4340
rect 28420 4284 36204 4340
rect 36260 4284 36270 4340
rect 39554 4284 39564 4340
rect 39620 4284 42140 4340
rect 42196 4284 42206 4340
rect 44258 4284 44268 4340
rect 44324 4284 52556 4340
rect 52612 4284 52622 4340
rect 7186 4172 7196 4228
rect 7252 4172 8988 4228
rect 9044 4172 9054 4228
rect 11330 4172 11340 4228
rect 11396 4172 16156 4228
rect 16212 4172 16222 4228
rect 52882 4172 52892 4228
rect 52948 4172 54124 4228
rect 54180 4172 54908 4228
rect 54964 4172 56700 4228
rect 56756 4172 56766 4228
rect 15138 4060 15148 4116
rect 15204 4060 15596 4116
rect 15652 4060 15662 4116
rect 28252 4060 28980 4116
rect 31042 4060 31052 4116
rect 31108 4060 40236 4116
rect 40292 4060 40302 4116
rect 50372 4060 51996 4116
rect 52052 4060 56588 4116
rect 56644 4060 56654 4116
rect 15362 3948 15372 4004
rect 15428 3948 17948 4004
rect 18004 3948 18014 4004
rect 20178 3948 20188 4004
rect 20244 3948 28028 4004
rect 28084 3948 28094 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 28252 3892 28308 4060
rect 18722 3836 18732 3892
rect 18788 3836 19292 3892
rect 19348 3836 28308 3892
rect 28924 3780 28980 4060
rect 50372 4004 50428 4060
rect 49746 3948 49756 4004
rect 49812 3948 50428 4004
rect 52546 3948 52556 4004
rect 52612 3948 57484 4004
rect 57540 3948 57550 4004
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 37314 3836 37324 3892
rect 37380 3836 38444 3892
rect 38500 3836 38510 3892
rect 45266 3836 45276 3892
rect 45332 3836 46172 3892
rect 46228 3836 48524 3892
rect 48580 3836 48590 3892
rect 49420 3836 50428 3892
rect 50484 3836 51996 3892
rect 52052 3836 52062 3892
rect 49420 3780 49476 3836
rect 10210 3724 10220 3780
rect 10276 3724 23212 3780
rect 23268 3724 23278 3780
rect 24322 3724 24332 3780
rect 24388 3724 25340 3780
rect 25396 3724 28364 3780
rect 28420 3724 28430 3780
rect 28924 3724 48748 3780
rect 48804 3724 49420 3780
rect 49476 3724 49486 3780
rect 49634 3724 49644 3780
rect 49700 3724 50204 3780
rect 50260 3724 57932 3780
rect 57988 3724 57998 3780
rect 8978 3612 8988 3668
rect 9044 3612 10108 3668
rect 10164 3612 10174 3668
rect 13570 3612 13580 3668
rect 13636 3612 16828 3668
rect 16884 3612 16894 3668
rect 24882 3612 24892 3668
rect 24948 3612 39228 3668
rect 39284 3612 40908 3668
rect 40964 3612 41692 3668
rect 41748 3612 41758 3668
rect 46722 3612 46732 3668
rect 46788 3612 48860 3668
rect 48916 3612 49308 3668
rect 49364 3612 51100 3668
rect 51156 3612 52892 3668
rect 52948 3612 52958 3668
rect 55234 3612 55244 3668
rect 55300 3612 57148 3668
rect 57204 3612 57214 3668
rect 12786 3500 12796 3556
rect 12852 3500 20188 3556
rect 20244 3500 20254 3556
rect 30482 3500 30492 3556
rect 30548 3500 31052 3556
rect 31108 3500 31118 3556
rect 48066 3500 48076 3556
rect 48132 3500 49756 3556
rect 49812 3500 49822 3556
rect 50530 3500 50540 3556
rect 50596 3500 52780 3556
rect 52836 3500 52846 3556
rect 4610 3388 4620 3444
rect 4676 3388 5404 3444
rect 5460 3388 5852 3444
rect 5908 3388 5918 3444
rect 28242 3388 28252 3444
rect 28308 3388 29372 3444
rect 29428 3388 29438 3444
rect 38434 3388 38444 3444
rect 38500 3388 42476 3444
rect 42532 3388 43932 3444
rect 43988 3388 43998 3444
rect 51762 3388 51772 3444
rect 51828 3388 53452 3444
rect 53508 3388 53518 3444
rect 11330 3276 11340 3332
rect 11396 3276 27020 3332
rect 27076 3276 27086 3332
rect 37650 3276 37660 3332
rect 37716 3276 57708 3332
rect 57764 3276 58268 3332
rect 58324 3276 58334 3332
rect 8306 3164 8316 3220
rect 8372 3164 13916 3220
rect 13972 3164 13982 3220
rect 15092 3164 16604 3220
rect 16660 3164 16670 3220
rect 15092 3108 15148 3164
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 3826 3052 3836 3108
rect 3892 3052 15148 3108
rect 2930 2940 2940 2996
rect 2996 2940 15652 2996
rect 15810 2940 15820 2996
rect 15876 2940 25676 2996
rect 25732 2940 25742 2996
rect 38994 2940 39004 2996
rect 39060 2940 56476 2996
rect 56532 2940 56542 2996
rect 15596 2884 15652 2940
rect 13906 2828 13916 2884
rect 13972 2828 15540 2884
rect 15596 2828 22988 2884
rect 23044 2828 23054 2884
rect 37090 2828 37100 2884
rect 37156 2828 49476 2884
rect 49634 2828 49644 2884
rect 49700 2828 56252 2884
rect 56308 2828 56318 2884
rect 1586 2716 1596 2772
rect 1652 2716 15260 2772
rect 15316 2716 15326 2772
rect 15484 2660 15540 2828
rect 49420 2772 49476 2828
rect 59200 2772 59800 2800
rect 15698 2716 15708 2772
rect 15764 2716 32844 2772
rect 32900 2716 32910 2772
rect 38098 2716 38108 2772
rect 38164 2716 49196 2772
rect 49252 2716 49262 2772
rect 49420 2716 52220 2772
rect 52276 2716 52286 2772
rect 55346 2716 55356 2772
rect 55412 2716 59800 2772
rect 59200 2688 59800 2716
rect 15484 2604 26348 2660
rect 26404 2604 26414 2660
rect 38322 2604 38332 2660
rect 38388 2604 57820 2660
rect 57876 2604 57886 2660
rect 4162 2492 4172 2548
rect 4228 2492 26012 2548
rect 26068 2492 26078 2548
rect 7186 2268 7196 2324
rect 7252 2268 26908 2324
rect 26964 2268 26974 2324
rect 18 1820 28 1876
rect 84 1820 1932 1876
rect 1988 1820 1998 1876
rect 4834 1596 4844 1652
rect 4900 1596 13692 1652
rect 13748 1596 26348 1652
rect 26404 1596 26414 1652
rect 39890 1596 39900 1652
rect 39956 1596 55468 1652
rect 55524 1596 55534 1652
rect 6178 1484 6188 1540
rect 6244 1484 26572 1540
rect 26628 1484 26638 1540
rect 37874 1484 37884 1540
rect 37940 1484 53900 1540
rect 53956 1484 53966 1540
rect 8306 1372 8316 1428
rect 8372 1372 27580 1428
rect 27636 1372 27646 1428
rect 3042 1260 3052 1316
rect 3108 1260 29148 1316
rect 29204 1260 29214 1316
<< via3 >>
rect 19836 56420 19892 56476
rect 19940 56420 19996 56476
rect 20044 56420 20100 56476
rect 50556 56420 50612 56476
rect 50660 56420 50716 56476
rect 50764 56420 50820 56476
rect 27692 55916 27748 55972
rect 4476 55636 4532 55692
rect 4580 55636 4636 55692
rect 4684 55636 4740 55692
rect 35196 55636 35252 55692
rect 35300 55636 35356 55692
rect 35404 55636 35460 55692
rect 19836 54852 19892 54908
rect 19940 54852 19996 54908
rect 20044 54852 20100 54908
rect 50556 54852 50612 54908
rect 50660 54852 50716 54908
rect 50764 54852 50820 54908
rect 4476 54068 4532 54124
rect 4580 54068 4636 54124
rect 4684 54068 4740 54124
rect 35196 54068 35252 54124
rect 35300 54068 35356 54124
rect 35404 54068 35460 54124
rect 19836 53284 19892 53340
rect 19940 53284 19996 53340
rect 20044 53284 20100 53340
rect 50556 53284 50612 53340
rect 50660 53284 50716 53340
rect 50764 53284 50820 53340
rect 4476 52500 4532 52556
rect 4580 52500 4636 52556
rect 4684 52500 4740 52556
rect 35196 52500 35252 52556
rect 35300 52500 35356 52556
rect 35404 52500 35460 52556
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 34748 49868 34804 49924
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 34748 48636 34804 48692
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 53900 48188 53956 48244
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 34300 46956 34356 47012
rect 55804 46508 55860 46564
rect 57708 46508 57764 46564
rect 20188 46396 20244 46452
rect 41692 46396 41748 46452
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 50316 46060 50372 46116
rect 57708 46060 57764 46116
rect 39452 45724 39508 45780
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 28140 45276 28196 45332
rect 55580 44940 55636 44996
rect 55468 44828 55524 44884
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 54236 44492 54292 44548
rect 34188 44380 34244 44436
rect 54684 44156 54740 44212
rect 55468 44044 55524 44100
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 40012 43708 40068 43764
rect 52556 43596 52612 43652
rect 53340 43372 53396 43428
rect 56700 43372 56756 43428
rect 52556 43260 52612 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 41692 43148 41748 43204
rect 43372 43148 43428 43204
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 26124 43036 26180 43092
rect 35644 42476 35700 42532
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 40012 42252 40068 42308
rect 54012 42140 54068 42196
rect 52444 42028 52500 42084
rect 35756 41916 35812 41972
rect 50316 41916 50372 41972
rect 56140 41804 56196 41860
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 52332 41468 52388 41524
rect 35644 41132 35700 41188
rect 53788 41020 53844 41076
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 52556 40572 52612 40628
rect 53116 40572 53172 40628
rect 53228 40348 53284 40404
rect 35644 40124 35700 40180
rect 52444 40124 52500 40180
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 53900 39900 53956 39956
rect 4060 39788 4116 39844
rect 43372 39676 43428 39732
rect 54236 39676 54292 39732
rect 42140 39564 42196 39620
rect 57708 39564 57764 39620
rect 25228 39340 25284 39396
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 14924 39116 14980 39172
rect 53564 39116 53620 39172
rect 42028 38892 42084 38948
rect 51996 38892 52052 38948
rect 3948 38780 4004 38836
rect 4060 38556 4116 38612
rect 15148 38556 15204 38612
rect 55804 38556 55860 38612
rect 41692 38444 41748 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 53564 38332 53620 38388
rect 3948 38220 4004 38276
rect 16604 38220 16660 38276
rect 54684 38220 54740 38276
rect 53452 38108 53508 38164
rect 16604 37996 16660 38052
rect 34300 37996 34356 38052
rect 41468 37884 41524 37940
rect 44380 37884 44436 37940
rect 50988 37772 51044 37828
rect 40796 37660 40852 37716
rect 51100 37660 51156 37716
rect 53788 37660 53844 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 11564 37436 11620 37492
rect 41468 37436 41524 37492
rect 42028 37324 42084 37380
rect 51212 37100 51268 37156
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 15148 36652 15204 36708
rect 53788 36876 53844 36932
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 38668 36652 38724 36708
rect 38556 36428 38612 36484
rect 53340 36428 53396 36484
rect 55468 36428 55524 36484
rect 11564 36316 11620 36372
rect 53340 36204 53396 36260
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 34188 35980 34244 36036
rect 53788 35868 53844 35924
rect 54012 35868 54068 35924
rect 16716 35644 16772 35700
rect 47180 35532 47236 35588
rect 53228 35532 53284 35588
rect 2268 35420 2324 35476
rect 34972 35420 35028 35476
rect 51996 35308 52052 35364
rect 56028 35308 56084 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 6300 34860 6356 34916
rect 44492 34748 44548 34804
rect 48972 34748 49028 34804
rect 53340 34748 53396 34804
rect 4956 34636 5012 34692
rect 47852 34636 47908 34692
rect 53900 34524 53956 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 9772 34412 9828 34468
rect 43932 34188 43988 34244
rect 7420 34076 7476 34132
rect 56140 34076 56196 34132
rect 56588 34076 56644 34132
rect 14812 33964 14868 34020
rect 44940 33964 44996 34020
rect 11788 33740 11844 33796
rect 12236 33740 12292 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 35644 33628 35700 33684
rect 44156 33628 44212 33684
rect 14924 33516 14980 33572
rect 51212 33516 51268 33572
rect 45948 33404 46004 33460
rect 50988 33292 51044 33348
rect 48076 33180 48132 33236
rect 51212 33180 51268 33236
rect 53564 33180 53620 33236
rect 49980 32956 50036 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 47180 32844 47236 32900
rect 29372 32732 29428 32788
rect 53452 32732 53508 32788
rect 34076 32508 34132 32564
rect 47516 32508 47572 32564
rect 50204 32508 50260 32564
rect 8652 32396 8708 32452
rect 40460 32396 40516 32452
rect 44492 32396 44548 32452
rect 17500 32284 17556 32340
rect 5628 32172 5684 32228
rect 43036 32172 43092 32228
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 8428 32060 8484 32116
rect 17276 32060 17332 32116
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 48636 32060 48692 32116
rect 49644 32060 49700 32116
rect 54012 32060 54068 32116
rect 52108 31948 52164 32004
rect 48636 31836 48692 31892
rect 46844 31724 46900 31780
rect 48860 31724 48916 31780
rect 51212 31724 51268 31780
rect 56476 31724 56532 31780
rect 6524 31612 6580 31668
rect 49980 31612 50036 31668
rect 53676 31612 53732 31668
rect 2380 31500 2436 31556
rect 4844 31500 4900 31556
rect 6412 31500 6468 31556
rect 38780 31500 38836 31556
rect 51212 31500 51268 31556
rect 15036 31388 15092 31444
rect 35756 31388 35812 31444
rect 53452 31388 53508 31444
rect 53676 31388 53732 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 50316 31276 50372 31332
rect 51436 31276 51492 31332
rect 4844 31164 4900 31220
rect 29484 31164 29540 31220
rect 5852 31052 5908 31108
rect 53116 31164 53172 31220
rect 55356 31164 55412 31220
rect 10668 30828 10724 30884
rect 3836 30716 3892 30772
rect 11788 30716 11844 30772
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 38668 30604 38724 30660
rect 49980 30604 50036 30660
rect 56588 30604 56644 30660
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 38444 30492 38500 30548
rect 43596 30492 43652 30548
rect 7756 30380 7812 30436
rect 29932 30380 29988 30436
rect 50372 30380 50428 30436
rect 18620 30268 18676 30324
rect 42252 30268 42308 30324
rect 40460 30156 40516 30212
rect 6412 30044 6468 30100
rect 18732 30044 18788 30100
rect 36652 30044 36708 30100
rect 55580 30044 55636 30100
rect 56588 30044 56644 30100
rect 5628 29932 5684 29988
rect 6300 29932 6356 29988
rect 8652 29932 8708 29988
rect 39116 29932 39172 29988
rect 4956 29820 5012 29876
rect 14476 29820 14532 29876
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 44044 29820 44100 29876
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 8652 29708 8708 29764
rect 55580 29708 55636 29764
rect 47180 29596 47236 29652
rect 48748 29596 48804 29652
rect 7308 29372 7364 29428
rect 44492 29372 44548 29428
rect 6636 29260 6692 29316
rect 7196 29260 7252 29316
rect 36540 29260 36596 29316
rect 19628 29148 19684 29204
rect 41692 29148 41748 29204
rect 49980 29148 50036 29204
rect 51436 29148 51492 29204
rect 7420 29036 7476 29092
rect 46732 29036 46788 29092
rect 49644 29036 49700 29092
rect 49868 29036 49924 29092
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 6524 28924 6580 28980
rect 16604 28924 16660 28980
rect 44156 28924 44212 28980
rect 56028 28924 56084 28980
rect 8428 28812 8484 28868
rect 7308 28700 7364 28756
rect 23100 28700 23156 28756
rect 36540 28700 36596 28756
rect 48860 28700 48916 28756
rect 40572 28588 40628 28644
rect 43596 28588 43652 28644
rect 48636 28588 48692 28644
rect 49644 28476 49700 28532
rect 7084 28364 7140 28420
rect 23436 28364 23492 28420
rect 52668 28364 52724 28420
rect 6636 28252 6692 28308
rect 9772 28252 9828 28308
rect 33628 28252 33684 28308
rect 54348 28252 54404 28308
rect 56252 28252 56308 28308
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 38444 28140 38500 28196
rect 49420 28140 49476 28196
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 19404 28028 19460 28084
rect 34076 28028 34132 28084
rect 39228 28028 39284 28084
rect 22316 27916 22372 27972
rect 40572 27916 40628 27972
rect 7420 27804 7476 27860
rect 4284 27692 4340 27748
rect 8316 27692 8372 27748
rect 11788 27692 11844 27748
rect 49308 27692 49364 27748
rect 54236 27580 54292 27636
rect 14028 27468 14084 27524
rect 14364 27468 14420 27524
rect 26236 27468 26292 27524
rect 43708 27468 43764 27524
rect 50204 27468 50260 27524
rect 54348 27468 54404 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 8428 27356 8484 27412
rect 24780 27356 24836 27412
rect 48524 27356 48580 27412
rect 52668 27356 52724 27412
rect 3500 27132 3556 27188
rect 6076 27132 6132 27188
rect 6860 27020 6916 27076
rect 14252 27244 14308 27300
rect 30940 27244 30996 27300
rect 39116 27244 39172 27300
rect 43372 27244 43428 27300
rect 53564 27244 53620 27300
rect 13804 27132 13860 27188
rect 36428 27132 36484 27188
rect 37212 27132 37268 27188
rect 40348 27132 40404 27188
rect 52332 27132 52388 27188
rect 54348 27132 54404 27188
rect 43260 27020 43316 27076
rect 43596 27020 43652 27076
rect 48524 27020 48580 27076
rect 8092 26908 8148 26964
rect 13804 26908 13860 26964
rect 38332 26908 38388 26964
rect 42588 26908 42644 26964
rect 46844 26908 46900 26964
rect 51548 26908 51604 26964
rect 54236 26908 54292 26964
rect 54908 26908 54964 26964
rect 7868 26796 7924 26852
rect 18620 26796 18676 26852
rect 28476 26796 28532 26852
rect 40908 26796 40964 26852
rect 43260 26796 43316 26852
rect 47852 26796 47908 26852
rect 50204 26796 50260 26852
rect 52220 26796 52276 26852
rect 6972 26684 7028 26740
rect 40684 26684 40740 26740
rect 42252 26684 42308 26740
rect 49532 26684 49588 26740
rect 51548 26684 51604 26740
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 3500 26572 3556 26628
rect 8092 26572 8148 26628
rect 10668 26572 10724 26628
rect 40348 26572 40404 26628
rect 43372 26572 43428 26628
rect 49084 26572 49140 26628
rect 3836 26460 3892 26516
rect 5740 26460 5796 26516
rect 40460 26460 40516 26516
rect 44044 26460 44100 26516
rect 44604 26460 44660 26516
rect 36764 26348 36820 26404
rect 41580 26348 41636 26404
rect 42140 26348 42196 26404
rect 47740 26348 47796 26404
rect 50316 26348 50372 26404
rect 7196 26236 7252 26292
rect 36428 26236 36484 26292
rect 39116 26236 39172 26292
rect 51100 26236 51156 26292
rect 54796 26236 54852 26292
rect 6748 26124 6804 26180
rect 11788 26124 11844 26180
rect 12236 26124 12292 26180
rect 17724 26124 17780 26180
rect 26012 26124 26068 26180
rect 41804 26124 41860 26180
rect 36428 26012 36484 26068
rect 44604 26012 44660 26068
rect 6748 25900 6804 25956
rect 7644 25900 7700 25956
rect 7868 25900 7924 25956
rect 13804 25900 13860 25956
rect 17500 25900 17556 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 49084 26012 49140 26068
rect 52220 26012 52276 26068
rect 56252 26012 56308 26068
rect 51324 25900 51380 25956
rect 12236 25788 12292 25844
rect 19516 25788 19572 25844
rect 55356 25788 55412 25844
rect 44492 25676 44548 25732
rect 48748 25676 48804 25732
rect 2268 25564 2324 25620
rect 6636 25564 6692 25620
rect 7196 25564 7252 25620
rect 9660 25564 9716 25620
rect 19180 25564 19236 25620
rect 52108 25564 52164 25620
rect 9324 25452 9380 25508
rect 11900 25452 11956 25508
rect 17276 25452 17332 25508
rect 40348 25452 40404 25508
rect 41468 25452 41524 25508
rect 44940 25452 44996 25508
rect 48076 25452 48132 25508
rect 48412 25452 48468 25508
rect 53676 25452 53732 25508
rect 56476 25452 56532 25508
rect 7644 25340 7700 25396
rect 14028 25340 14084 25396
rect 17052 25340 17108 25396
rect 49532 25340 49588 25396
rect 3948 25228 4004 25284
rect 33516 25228 33572 25284
rect 35644 25228 35700 25284
rect 41020 25228 41076 25284
rect 41804 25228 41860 25284
rect 42476 25228 42532 25284
rect 43036 25228 43092 25284
rect 3724 25116 3780 25172
rect 6412 25116 6468 25172
rect 7420 25116 7476 25172
rect 25340 25116 25396 25172
rect 30940 25116 30996 25172
rect 36764 25116 36820 25172
rect 37212 25116 37268 25172
rect 43596 25116 43652 25172
rect 46956 25116 47012 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 7308 25004 7364 25060
rect 39228 25004 39284 25060
rect 57484 25004 57540 25060
rect 11900 24892 11956 24948
rect 19180 24892 19236 24948
rect 40908 24892 40964 24948
rect 48188 24892 48244 24948
rect 51212 24892 51268 24948
rect 6076 24780 6132 24836
rect 7308 24780 7364 24836
rect 7532 24780 7588 24836
rect 9772 24780 9828 24836
rect 46732 24780 46788 24836
rect 4844 24668 4900 24724
rect 15260 24668 15316 24724
rect 16716 24668 16772 24724
rect 18732 24668 18788 24724
rect 44156 24668 44212 24724
rect 48860 24668 48916 24724
rect 53116 24668 53172 24724
rect 3948 24556 4004 24612
rect 29260 24556 29316 24612
rect 36876 24556 36932 24612
rect 51884 24556 51940 24612
rect 9324 24444 9380 24500
rect 9996 24444 10052 24500
rect 19516 24444 19572 24500
rect 35756 24444 35812 24500
rect 43484 24444 43540 24500
rect 48636 24444 48692 24500
rect 6636 24332 6692 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 12348 24220 12404 24276
rect 14812 24220 14868 24276
rect 19068 24220 19124 24276
rect 25340 24220 25396 24276
rect 51324 24220 51380 24276
rect 5852 24108 5908 24164
rect 15148 24108 15204 24164
rect 42588 24108 42644 24164
rect 49532 24108 49588 24164
rect 52444 24108 52500 24164
rect 16940 23996 16996 24052
rect 40684 23996 40740 24052
rect 41692 23996 41748 24052
rect 42700 23996 42756 24052
rect 49308 23996 49364 24052
rect 6524 23884 6580 23940
rect 6748 23884 6804 23940
rect 7196 23884 7252 23940
rect 7420 23884 7476 23940
rect 10668 23884 10724 23940
rect 11676 23884 11732 23940
rect 3724 23772 3780 23828
rect 5964 23660 6020 23716
rect 48188 23884 48244 23940
rect 9772 23772 9828 23828
rect 42588 23772 42644 23828
rect 49308 23772 49364 23828
rect 4284 23548 4340 23604
rect 6748 23548 6804 23604
rect 7532 23660 7588 23716
rect 14476 23660 14532 23716
rect 15596 23660 15652 23716
rect 20300 23660 20356 23716
rect 35644 23660 35700 23716
rect 38108 23660 38164 23716
rect 38332 23660 38388 23716
rect 38780 23660 38836 23716
rect 48076 23660 48132 23716
rect 48636 23660 48692 23716
rect 50204 23660 50260 23716
rect 51324 23660 51380 23716
rect 9996 23548 10052 23604
rect 15036 23548 15092 23604
rect 36652 23548 36708 23604
rect 36988 23548 37044 23604
rect 47852 23548 47908 23604
rect 7420 23436 7476 23492
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 18956 23436 19012 23492
rect 40348 23436 40404 23492
rect 42700 23436 42756 23492
rect 49084 23436 49140 23492
rect 13468 23324 13524 23380
rect 19516 23324 19572 23380
rect 43036 23324 43092 23380
rect 48524 23324 48580 23380
rect 33404 23212 33460 23268
rect 28476 23100 28532 23156
rect 40124 23212 40180 23268
rect 42476 23100 42532 23156
rect 47404 23100 47460 23156
rect 50204 23436 50260 23492
rect 56924 23436 56980 23492
rect 57484 23436 57540 23492
rect 55244 23324 55300 23380
rect 52444 23212 52500 23268
rect 56028 23212 56084 23268
rect 50204 23100 50260 23156
rect 16492 22988 16548 23044
rect 17724 22988 17780 23044
rect 43820 22988 43876 23044
rect 49308 22988 49364 23044
rect 49532 22988 49588 23044
rect 50092 22988 50148 23044
rect 53228 22988 53284 23044
rect 7420 22876 7476 22932
rect 11900 22876 11956 22932
rect 24332 22876 24388 22932
rect 40124 22876 40180 22932
rect 47068 22876 47124 22932
rect 49644 22876 49700 22932
rect 52332 22876 52388 22932
rect 56924 22876 56980 22932
rect 23548 22764 23604 22820
rect 25900 22764 25956 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 15372 22652 15428 22708
rect 26460 22652 26516 22708
rect 36988 22652 37044 22708
rect 38444 22652 38500 22708
rect 41692 22652 41748 22708
rect 19180 22540 19236 22596
rect 27020 22540 27076 22596
rect 49756 22540 49812 22596
rect 51436 22540 51492 22596
rect 55468 22540 55524 22596
rect 15036 22428 15092 22484
rect 17724 22428 17780 22484
rect 18732 22428 18788 22484
rect 26572 22428 26628 22484
rect 40236 22428 40292 22484
rect 55804 22428 55860 22484
rect 2380 22316 2436 22372
rect 6412 22316 6468 22372
rect 16492 22316 16548 22372
rect 48636 22316 48692 22372
rect 51436 22316 51492 22372
rect 52556 22316 52612 22372
rect 55020 22316 55076 22372
rect 28812 22204 28868 22260
rect 33516 22204 33572 22260
rect 37996 22204 38052 22260
rect 38556 22204 38612 22260
rect 46620 22204 46676 22260
rect 48524 22204 48580 22260
rect 49308 22204 49364 22260
rect 56924 22204 56980 22260
rect 18508 22092 18564 22148
rect 13244 21980 13300 22036
rect 19180 21980 19236 22036
rect 24220 21980 24276 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 38108 22092 38164 22148
rect 40012 22092 40068 22148
rect 41692 22092 41748 22148
rect 49756 22092 49812 22148
rect 50092 22092 50148 22148
rect 51212 22092 51268 22148
rect 51660 21980 51716 22036
rect 51996 21980 52052 22036
rect 57372 21980 57428 22036
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 40572 21868 40628 21924
rect 41692 21868 41748 21924
rect 48188 21868 48244 21924
rect 51100 21868 51156 21924
rect 8316 21756 8372 21812
rect 18732 21756 18788 21812
rect 24444 21756 24500 21812
rect 32732 21756 32788 21812
rect 35980 21756 36036 21812
rect 44156 21756 44212 21812
rect 47404 21756 47460 21812
rect 48300 21756 48356 21812
rect 18508 21644 18564 21700
rect 22316 21644 22372 21700
rect 30044 21644 30100 21700
rect 47964 21644 48020 21700
rect 53228 21644 53284 21700
rect 55244 21644 55300 21700
rect 56364 21644 56420 21700
rect 7980 21532 8036 21588
rect 13356 21532 13412 21588
rect 24332 21532 24388 21588
rect 29260 21532 29316 21588
rect 44044 21532 44100 21588
rect 47516 21532 47572 21588
rect 48300 21532 48356 21588
rect 49308 21532 49364 21588
rect 50204 21532 50260 21588
rect 16604 21420 16660 21476
rect 18732 21420 18788 21476
rect 39004 21420 39060 21476
rect 48188 21420 48244 21476
rect 48636 21420 48692 21476
rect 53340 21420 53396 21476
rect 53676 21420 53732 21476
rect 54684 21420 54740 21476
rect 6972 21308 7028 21364
rect 20300 21308 20356 21364
rect 40572 21308 40628 21364
rect 49644 21308 49700 21364
rect 51436 21308 51492 21364
rect 23772 21196 23828 21252
rect 33516 21196 33572 21252
rect 46620 21196 46676 21252
rect 47068 21196 47124 21252
rect 53228 21196 53284 21252
rect 55468 21196 55524 21252
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 18396 21084 18452 21140
rect 54124 21084 54180 21140
rect 35644 20972 35700 21028
rect 40348 20972 40404 21028
rect 44156 20972 44212 21028
rect 45836 20972 45892 21028
rect 49756 20972 49812 21028
rect 25228 20860 25284 20916
rect 41132 20860 41188 20916
rect 43708 20860 43764 20916
rect 45612 20860 45668 20916
rect 46956 20860 47012 20916
rect 51100 20860 51156 20916
rect 40908 20748 40964 20804
rect 41468 20748 41524 20804
rect 42812 20748 42868 20804
rect 51884 20748 51940 20804
rect 53900 20748 53956 20804
rect 57708 20748 57764 20804
rect 38556 20636 38612 20692
rect 40460 20636 40516 20692
rect 47404 20636 47460 20692
rect 48300 20636 48356 20692
rect 22876 20524 22932 20580
rect 37436 20524 37492 20580
rect 43932 20524 43988 20580
rect 48636 20524 48692 20580
rect 48860 20524 48916 20580
rect 49980 20524 50036 20580
rect 3612 20412 3668 20468
rect 16716 20412 16772 20468
rect 20748 20412 20804 20468
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 35756 20412 35812 20468
rect 36876 20412 36932 20468
rect 41468 20412 41524 20468
rect 45612 20412 45668 20468
rect 48748 20412 48804 20468
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 25900 20300 25956 20356
rect 40684 20300 40740 20356
rect 50316 20300 50372 20356
rect 19404 20188 19460 20244
rect 24444 20188 24500 20244
rect 43484 20188 43540 20244
rect 51212 20188 51268 20244
rect 51884 20188 51940 20244
rect 4956 20076 5012 20132
rect 29820 20076 29876 20132
rect 49420 20076 49476 20132
rect 19068 19964 19124 20020
rect 19292 19964 19348 20020
rect 31724 19964 31780 20020
rect 41020 19964 41076 20020
rect 44268 19964 44324 20020
rect 50204 19964 50260 20020
rect 51660 19964 51716 20020
rect 5740 19852 5796 19908
rect 13580 19852 13636 19908
rect 13916 19852 13972 19908
rect 24332 19852 24388 19908
rect 37996 19852 38052 19908
rect 40236 19852 40292 19908
rect 43372 19740 43428 19796
rect 49532 19740 49588 19796
rect 51548 19740 51604 19796
rect 51996 19740 52052 19796
rect 23548 19628 23604 19684
rect 23772 19628 23828 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 15820 19516 15876 19572
rect 24556 19516 24612 19572
rect 40012 19516 40068 19572
rect 44044 19516 44100 19572
rect 54908 19516 54964 19572
rect 13356 19404 13412 19460
rect 13580 19404 13636 19460
rect 30044 19404 30100 19460
rect 38668 19404 38724 19460
rect 49644 19404 49700 19460
rect 53116 19404 53172 19460
rect 54012 19404 54068 19460
rect 10332 19292 10388 19348
rect 19628 19292 19684 19348
rect 26460 19292 26516 19348
rect 45948 19292 46004 19348
rect 48972 19292 49028 19348
rect 55132 19292 55188 19348
rect 13692 19180 13748 19236
rect 15260 19180 15316 19236
rect 42812 19180 42868 19236
rect 47404 19180 47460 19236
rect 15148 19068 15204 19124
rect 57260 19068 57316 19124
rect 3724 18956 3780 19012
rect 17164 18956 17220 19012
rect 18172 18956 18228 19012
rect 22876 18956 22932 19012
rect 24220 18956 24276 19012
rect 26460 18956 26516 19012
rect 55132 18956 55188 19012
rect 55468 18956 55524 19012
rect 56476 18956 56532 19012
rect 18508 18844 18564 18900
rect 40796 18844 40852 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 52444 18844 52500 18900
rect 11676 18732 11732 18788
rect 12124 18732 12180 18788
rect 12348 18732 12404 18788
rect 18172 18732 18228 18788
rect 37100 18732 37156 18788
rect 49308 18732 49364 18788
rect 49756 18732 49812 18788
rect 52108 18732 52164 18788
rect 52892 18732 52948 18788
rect 54460 18732 54516 18788
rect 12460 18620 12516 18676
rect 15708 18620 15764 18676
rect 23324 18620 23380 18676
rect 26236 18620 26292 18676
rect 43484 18620 43540 18676
rect 6636 18508 6692 18564
rect 12124 18508 12180 18564
rect 15820 18508 15876 18564
rect 39116 18508 39172 18564
rect 56476 18620 56532 18676
rect 47404 18508 47460 18564
rect 3724 18396 3780 18452
rect 3948 18396 4004 18452
rect 16940 18396 16996 18452
rect 18956 18396 19012 18452
rect 19180 18396 19236 18452
rect 40684 18396 40740 18452
rect 43036 18396 43092 18452
rect 49532 18396 49588 18452
rect 52108 18396 52164 18452
rect 4284 18284 4340 18340
rect 21868 18284 21924 18340
rect 25676 18284 25732 18340
rect 40908 18284 40964 18340
rect 51100 18284 51156 18340
rect 13244 18172 13300 18228
rect 13468 18172 13524 18228
rect 15708 18172 15764 18228
rect 23548 18172 23604 18228
rect 36876 18172 36932 18228
rect 37100 18172 37156 18228
rect 47964 18172 48020 18228
rect 48636 18172 48692 18228
rect 52220 18172 52276 18228
rect 53564 18172 53620 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 7196 18060 7252 18116
rect 16828 18060 16884 18116
rect 19068 18060 19124 18116
rect 21868 18060 21924 18116
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 11676 17948 11732 18004
rect 13356 17948 13412 18004
rect 19180 17948 19236 18004
rect 26012 17948 26068 18004
rect 43820 17948 43876 18004
rect 50092 17948 50148 18004
rect 52108 17948 52164 18004
rect 52444 17948 52500 18004
rect 4060 17724 4116 17780
rect 8204 17724 8260 17780
rect 17164 17836 17220 17892
rect 18844 17836 18900 17892
rect 19516 17836 19572 17892
rect 40348 17836 40404 17892
rect 54124 17836 54180 17892
rect 9660 17724 9716 17780
rect 16268 17724 16324 17780
rect 23660 17724 23716 17780
rect 37436 17724 37492 17780
rect 43596 17724 43652 17780
rect 47180 17724 47236 17780
rect 52108 17724 52164 17780
rect 52332 17724 52388 17780
rect 4172 17612 4228 17668
rect 5068 17612 5124 17668
rect 8316 17612 8372 17668
rect 13468 17612 13524 17668
rect 9660 17500 9716 17556
rect 26684 17612 26740 17668
rect 45836 17612 45892 17668
rect 46844 17612 46900 17668
rect 49644 17612 49700 17668
rect 18396 17500 18452 17556
rect 21420 17500 21476 17556
rect 34972 17500 35028 17556
rect 44044 17500 44100 17556
rect 46172 17500 46228 17556
rect 4844 17388 4900 17444
rect 23324 17388 23380 17444
rect 35644 17388 35700 17444
rect 44268 17388 44324 17444
rect 45276 17388 45332 17444
rect 54908 17388 54964 17444
rect 57260 17388 57316 17444
rect 18956 17276 19012 17332
rect 41580 17276 41636 17332
rect 46396 17276 46452 17332
rect 49084 17276 49140 17332
rect 7308 17164 7364 17220
rect 6412 17052 6468 17108
rect 11900 17052 11956 17108
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 26348 17052 26404 17108
rect 35980 17052 36036 17108
rect 41804 17052 41860 17108
rect 43036 17052 43092 17108
rect 47964 17052 48020 17108
rect 49980 17052 50036 17108
rect 53564 17052 53620 17108
rect 54460 17052 54516 17108
rect 5404 16940 5460 16996
rect 6860 16940 6916 16996
rect 40012 16940 40068 16996
rect 43596 16940 43652 16996
rect 50316 16940 50372 16996
rect 13244 16828 13300 16884
rect 18844 16828 18900 16884
rect 19628 16828 19684 16884
rect 25228 16828 25284 16884
rect 40572 16828 40628 16884
rect 41132 16828 41188 16884
rect 5852 16716 5908 16772
rect 16268 16716 16324 16772
rect 3612 16604 3668 16660
rect 7420 16604 7476 16660
rect 8204 16604 8260 16660
rect 15372 16604 15428 16660
rect 16156 16604 16212 16660
rect 23436 16604 23492 16660
rect 26572 16604 26628 16660
rect 43372 16604 43428 16660
rect 43820 16604 43876 16660
rect 7532 16492 7588 16548
rect 38444 16492 38500 16548
rect 51884 16492 51940 16548
rect 52668 16492 52724 16548
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 28812 16380 28868 16436
rect 48748 16380 48804 16436
rect 51324 16380 51380 16436
rect 11788 16268 11844 16324
rect 16044 16268 16100 16324
rect 23548 16268 23604 16324
rect 51436 16268 51492 16324
rect 57372 16268 57428 16324
rect 4172 16044 4228 16100
rect 23660 16156 23716 16212
rect 39564 16156 39620 16212
rect 46844 16156 46900 16212
rect 18732 16044 18788 16100
rect 24556 16044 24612 16100
rect 26460 16044 26516 16100
rect 29932 16044 29988 16100
rect 30828 16044 30884 16100
rect 23324 15932 23380 15988
rect 25228 15932 25284 15988
rect 43932 16044 43988 16100
rect 49644 16044 49700 16100
rect 44156 15932 44212 15988
rect 53676 15932 53732 15988
rect 54460 15932 54516 15988
rect 7532 15820 7588 15876
rect 19404 15820 19460 15876
rect 39900 15820 39956 15876
rect 8092 15708 8148 15764
rect 26684 15708 26740 15764
rect 37100 15708 37156 15764
rect 38668 15708 38724 15764
rect 49756 15708 49812 15764
rect 51996 15708 52052 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 10220 15596 10276 15652
rect 16716 15596 16772 15652
rect 18732 15596 18788 15652
rect 20524 15596 20580 15652
rect 35644 15596 35700 15652
rect 46284 15596 46340 15652
rect 47740 15596 47796 15652
rect 53452 15596 53508 15652
rect 55468 15596 55524 15652
rect 5292 15484 5348 15540
rect 6412 15484 6468 15540
rect 18172 15484 18228 15540
rect 23548 15484 23604 15540
rect 24780 15484 24836 15540
rect 31724 15484 31780 15540
rect 39564 15484 39620 15540
rect 40460 15484 40516 15540
rect 44380 15484 44436 15540
rect 46508 15484 46564 15540
rect 51884 15484 51940 15540
rect 56588 15484 56644 15540
rect 6860 15372 6916 15428
rect 9660 15372 9716 15428
rect 18844 15372 18900 15428
rect 19516 15372 19572 15428
rect 20300 15372 20356 15428
rect 43708 15372 43764 15428
rect 11676 15260 11732 15316
rect 29820 15260 29876 15316
rect 46844 15260 46900 15316
rect 48524 15260 48580 15316
rect 52668 15260 52724 15316
rect 57708 15260 57764 15316
rect 4172 15148 4228 15204
rect 23436 15148 23492 15204
rect 23772 15148 23828 15204
rect 42028 15148 42084 15204
rect 47740 15148 47796 15204
rect 49756 15148 49812 15204
rect 50988 15148 51044 15204
rect 7420 15036 7476 15092
rect 11900 15036 11956 15092
rect 19068 15036 19124 15092
rect 46284 15036 46340 15092
rect 51100 15036 51156 15092
rect 4172 14924 4228 14980
rect 6524 14924 6580 14980
rect 37100 14924 37156 14980
rect 39564 14924 39620 14980
rect 48524 14924 48580 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 5740 14812 5796 14868
rect 8540 14812 8596 14868
rect 21420 14812 21476 14868
rect 9660 14700 9716 14756
rect 48412 14700 48468 14756
rect 7644 14588 7700 14644
rect 8652 14588 8708 14644
rect 13916 14588 13972 14644
rect 18620 14588 18676 14644
rect 23100 14588 23156 14644
rect 27020 14588 27076 14644
rect 39116 14588 39172 14644
rect 47852 14588 47908 14644
rect 49868 14588 49924 14644
rect 53340 14588 53396 14644
rect 3612 14476 3668 14532
rect 6188 14476 6244 14532
rect 6972 14476 7028 14532
rect 8876 14476 8932 14532
rect 16604 14476 16660 14532
rect 20524 14476 20580 14532
rect 39452 14476 39508 14532
rect 53676 14476 53732 14532
rect 41692 14364 41748 14420
rect 48636 14364 48692 14420
rect 3612 14252 3668 14308
rect 4060 14252 4116 14308
rect 7980 14252 8036 14308
rect 11564 14252 11620 14308
rect 23436 14252 23492 14308
rect 49532 14252 49588 14308
rect 56028 14252 56084 14308
rect 3500 14140 3556 14196
rect 23324 14140 23380 14196
rect 46620 14140 46676 14196
rect 49644 14140 49700 14196
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 5292 14028 5348 14084
rect 6860 14028 6916 14084
rect 10332 14028 10388 14084
rect 15596 14028 15652 14084
rect 19068 14028 19124 14084
rect 5068 13916 5124 13972
rect 15932 13916 15988 13972
rect 16380 13916 16436 13972
rect 23660 13916 23716 13972
rect 24220 13916 24276 13972
rect 33404 13916 33460 13972
rect 44156 13916 44212 13972
rect 45276 13916 45332 13972
rect 46396 13916 46452 13972
rect 51100 13916 51156 13972
rect 6524 13804 6580 13860
rect 7644 13804 7700 13860
rect 8652 13804 8708 13860
rect 19180 13804 19236 13860
rect 52108 13804 52164 13860
rect 53228 13804 53284 13860
rect 6636 13692 6692 13748
rect 8204 13692 8260 13748
rect 26348 13692 26404 13748
rect 4956 13468 5012 13524
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 13468 13580 13524 13636
rect 17052 13580 17108 13636
rect 18732 13580 18788 13636
rect 23436 13580 23492 13636
rect 41580 13580 41636 13636
rect 41916 13580 41972 13636
rect 47068 13580 47124 13636
rect 53900 13580 53956 13636
rect 43820 13468 43876 13524
rect 50204 13356 50260 13412
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 21868 13244 21924 13300
rect 41692 13244 41748 13300
rect 51100 13244 51156 13300
rect 3500 13132 3556 13188
rect 5852 13132 5908 13188
rect 18956 13132 19012 13188
rect 19628 13132 19684 13188
rect 42140 13132 42196 13188
rect 56364 13132 56420 13188
rect 7756 13020 7812 13076
rect 8092 13020 8148 13076
rect 16380 13020 16436 13076
rect 30828 13020 30884 13076
rect 51996 13020 52052 13076
rect 2044 12908 2100 12964
rect 4956 12908 5012 12964
rect 7196 12908 7252 12964
rect 20300 12908 20356 12964
rect 20524 12908 20580 12964
rect 40236 12908 40292 12964
rect 40572 12908 40628 12964
rect 51100 12908 51156 12964
rect 4284 12796 4340 12852
rect 6188 12796 6244 12852
rect 15036 12796 15092 12852
rect 19404 12796 19460 12852
rect 39452 12796 39508 12852
rect 49644 12796 49700 12852
rect 9324 12684 9380 12740
rect 10108 12684 10164 12740
rect 15820 12684 15876 12740
rect 16268 12684 16324 12740
rect 19628 12684 19684 12740
rect 21420 12684 21476 12740
rect 23324 12684 23380 12740
rect 18508 12572 18564 12628
rect 49532 12572 49588 12628
rect 49756 12572 49812 12628
rect 52556 12572 52612 12628
rect 3724 12460 3780 12516
rect 18956 12460 19012 12516
rect 3948 12348 4004 12404
rect 4956 12348 5012 12404
rect 15148 12348 15204 12404
rect 16828 12348 16884 12404
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 19404 12460 19460 12516
rect 43932 12460 43988 12516
rect 46172 12460 46228 12516
rect 48748 12348 48804 12404
rect 55132 12348 55188 12404
rect 50316 12236 50372 12292
rect 18172 12124 18228 12180
rect 24220 12124 24276 12180
rect 54908 12124 54964 12180
rect 7308 12012 7364 12068
rect 10108 12012 10164 12068
rect 17052 12012 17108 12068
rect 47180 11900 47236 11956
rect 12460 11788 12516 11844
rect 19628 11788 19684 11844
rect 29484 11788 29540 11844
rect 49532 11788 49588 11844
rect 55020 11788 55076 11844
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 8316 11676 8372 11732
rect 16604 11676 16660 11732
rect 16828 11676 16884 11732
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 50316 11676 50372 11732
rect 8204 11564 8260 11620
rect 14924 11564 14980 11620
rect 48076 11564 48132 11620
rect 52108 11564 52164 11620
rect 54908 11564 54964 11620
rect 22764 11452 22820 11508
rect 43036 11452 43092 11508
rect 53564 11452 53620 11508
rect 14924 11340 14980 11396
rect 16604 11340 16660 11396
rect 20748 11340 20804 11396
rect 8316 11228 8372 11284
rect 41804 11116 41860 11172
rect 54796 11116 54852 11172
rect 46508 11004 46564 11060
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 43596 10892 43652 10948
rect 7420 10780 7476 10836
rect 35756 10780 35812 10836
rect 2156 10668 2212 10724
rect 2380 10668 2436 10724
rect 4956 10556 5012 10612
rect 7644 10556 7700 10612
rect 28140 10556 28196 10612
rect 17724 10444 17780 10500
rect 56476 10444 56532 10500
rect 20300 10332 20356 10388
rect 13916 10220 13972 10276
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 5404 10108 5460 10164
rect 51548 10108 51604 10164
rect 10556 9996 10612 10052
rect 48860 9996 48916 10052
rect 56924 9996 56980 10052
rect 15932 9884 15988 9940
rect 43484 9772 43540 9828
rect 54684 9772 54740 9828
rect 6636 9436 6692 9492
rect 14812 9436 14868 9492
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 15932 9324 15988 9380
rect 16604 9324 16660 9380
rect 10220 9212 10276 9268
rect 11676 9212 11732 9268
rect 13692 9212 13748 9268
rect 15148 9212 15204 9268
rect 16156 9212 16212 9268
rect 3948 9100 4004 9156
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 48300 9212 48356 9268
rect 51884 9212 51940 9268
rect 51100 8988 51156 9044
rect 5628 8876 5684 8932
rect 14812 8876 14868 8932
rect 50316 8876 50372 8932
rect 19068 8764 19124 8820
rect 56924 8764 56980 8820
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 4956 8428 5012 8484
rect 12236 8428 12292 8484
rect 16044 8316 16100 8372
rect 32732 8316 32788 8372
rect 52892 8316 52948 8372
rect 49980 8204 50036 8260
rect 51436 8204 51492 8260
rect 27692 7868 27748 7924
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 41916 7756 41972 7812
rect 53788 7756 53844 7812
rect 19516 7644 19572 7700
rect 47964 7644 48020 7700
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 15036 6860 15092 6916
rect 17276 6748 17332 6804
rect 29372 6748 29428 6804
rect 22764 6524 22820 6580
rect 47740 6524 47796 6580
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 5628 6188 5684 6244
rect 3948 6076 4004 6132
rect 56028 6076 56084 6132
rect 9660 5740 9716 5796
rect 19068 5740 19124 5796
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 47740 5404 47796 5460
rect 2044 5180 2100 5236
rect 3948 5180 4004 5236
rect 9660 5180 9716 5236
rect 10556 5180 10612 5236
rect 11564 5180 11620 5236
rect 22988 5180 23044 5236
rect 2156 5068 2212 5124
rect 33628 5068 33684 5124
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 20188 4620 20244 4676
rect 10108 4508 10164 4564
rect 28364 4284 28420 4340
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 10220 3724 10276 3780
rect 28364 3724 28420 3780
rect 8316 3164 8372 3220
rect 16604 3164 16660 3220
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 15820 2940 15876 2996
rect 25676 2940 25732 2996
rect 39004 2940 39060 2996
rect 56476 2940 56532 2996
rect 22988 2828 23044 2884
rect 49644 2828 49700 2884
rect 15260 2716 15316 2772
rect 15708 2716 15764 2772
rect 49196 2716 49252 2772
rect 38332 2604 38388 2660
rect 4844 1596 4900 1652
rect 13692 1596 13748 1652
rect 26348 1596 26404 1652
rect 39900 1596 39956 1652
rect 26572 1484 26628 1540
<< metal4 >>
rect 4448 55692 4768 56508
rect 4448 55636 4476 55692
rect 4532 55636 4580 55692
rect 4636 55636 4684 55692
rect 4740 55636 4768 55692
rect 4448 54124 4768 55636
rect 4448 54068 4476 54124
rect 4532 54068 4580 54124
rect 4636 54068 4684 54124
rect 4740 54068 4768 54124
rect 4448 52556 4768 54068
rect 4448 52500 4476 52556
rect 4532 52500 4580 52556
rect 4636 52500 4684 52556
rect 4740 52500 4768 52556
rect 4448 50988 4768 52500
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4060 39844 4116 39854
rect 3948 38836 4004 38846
rect 3948 38276 4004 38780
rect 4060 38612 4116 39788
rect 4060 38546 4116 38556
rect 3948 38210 4004 38220
rect 4448 38444 4768 39956
rect 19808 56476 20128 56508
rect 19808 56420 19836 56476
rect 19892 56420 19940 56476
rect 19996 56420 20044 56476
rect 20100 56420 20128 56476
rect 19808 54908 20128 56420
rect 19808 54852 19836 54908
rect 19892 54852 19940 54908
rect 19996 54852 20044 54908
rect 20100 54852 20128 54908
rect 19808 53340 20128 54852
rect 19808 53284 19836 53340
rect 19892 53284 19940 53340
rect 19996 53284 20044 53340
rect 20100 53284 20128 53340
rect 19808 51772 20128 53284
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 19808 45500 20128 47012
rect 27692 55972 27748 55982
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 14924 39172 14980 39182
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 2268 35476 2324 35486
rect 2268 25620 2324 35420
rect 4448 35308 4768 36820
rect 11564 37492 11620 37502
rect 11564 36372 11620 37436
rect 11564 36306 11620 36316
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 6300 34916 6356 34926
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 2268 25554 2324 25564
rect 2380 31556 2436 31566
rect 2380 22372 2436 31500
rect 3836 30772 3892 30782
rect 3500 27188 3556 27198
rect 3500 26628 3556 27132
rect 3500 26562 3556 26572
rect 3836 26516 3892 30716
rect 4448 30604 4768 32116
rect 4956 34692 5012 34702
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 3836 26450 3892 26460
rect 4284 27748 4340 27758
rect 3948 25284 4004 25294
rect 3724 25172 3780 25182
rect 3724 23828 3780 25116
rect 3948 24612 4004 25228
rect 3948 24546 4004 24556
rect 3724 23762 3780 23772
rect 4284 23604 4340 27692
rect 4284 23538 4340 23548
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4844 31556 4900 31566
rect 4844 31220 4900 31500
rect 4844 24724 4900 31164
rect 4956 29876 5012 34636
rect 5628 32228 5684 32238
rect 5628 29988 5684 32172
rect 5628 29922 5684 29932
rect 5852 31108 5908 31118
rect 4956 29810 5012 29820
rect 4844 24658 4900 24668
rect 5740 26516 5796 26526
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 2044 12964 2100 12974
rect 2044 5236 2100 12908
rect 2044 5170 2100 5180
rect 2156 10724 2212 10734
rect 2156 5124 2212 10668
rect 2380 10724 2436 22316
rect 4448 22764 4768 24276
rect 5740 23548 5796 26460
rect 5852 24164 5908 31052
rect 6300 29988 6356 34860
rect 9772 34468 9828 34478
rect 7420 34132 7476 34142
rect 6524 31668 6580 31678
rect 6300 29922 6356 29932
rect 6412 31556 6468 31566
rect 6412 30100 6468 31500
rect 6076 27188 6132 27198
rect 6076 24836 6132 27132
rect 6412 25172 6468 30044
rect 6524 28980 6580 31612
rect 7308 29428 7364 29438
rect 6524 25284 6580 28924
rect 6636 29316 6692 29326
rect 6636 28308 6692 29260
rect 7196 29316 7252 29326
rect 6636 25620 6692 28252
rect 7084 28420 7140 28430
rect 6860 27076 6916 27086
rect 6748 26180 6804 26190
rect 6748 25956 6804 26124
rect 6748 25890 6804 25900
rect 6636 25554 6692 25564
rect 6524 25228 6804 25284
rect 6412 25106 6468 25116
rect 6076 24770 6132 24780
rect 6636 24388 6692 24398
rect 5852 24098 5908 24108
rect 6300 24332 6636 24388
rect 6300 24052 6356 24332
rect 6636 24322 6692 24332
rect 6748 24164 6804 25228
rect 5964 23996 6356 24052
rect 6412 24108 6804 24164
rect 5964 23716 6020 23996
rect 5964 23650 6020 23660
rect 5740 23492 6244 23548
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 3612 20468 3668 20478
rect 3612 16660 3668 20412
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 3612 16594 3668 16604
rect 3724 19012 3780 19022
rect 3724 18452 3780 18956
rect 3612 14532 3668 14542
rect 3612 14308 3668 14476
rect 3612 14242 3668 14252
rect 3500 14196 3556 14206
rect 3500 13188 3556 14140
rect 3500 13122 3556 13132
rect 3724 12516 3780 18396
rect 3724 12450 3780 12460
rect 3948 18452 4004 18462
rect 3948 12404 4004 18396
rect 4284 18340 4340 18350
rect 4060 17780 4116 17790
rect 4060 14308 4116 17724
rect 4172 17668 4228 17678
rect 4172 16100 4228 17612
rect 4172 16034 4228 16044
rect 4172 15204 4228 15214
rect 4172 14980 4228 15148
rect 4172 14914 4228 14924
rect 4060 14242 4116 14252
rect 4284 12852 4340 18284
rect 4284 12786 4340 12796
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4956 20132 5012 20142
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 3948 12338 4004 12348
rect 2380 10658 2436 10668
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 3948 9156 4004 9166
rect 3948 6132 4004 9100
rect 3948 5236 4004 6076
rect 3948 5170 4004 5180
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 2156 5058 2212 5068
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 4844 17444 4900 17454
rect 4844 1652 4900 17388
rect 4956 13524 5012 20076
rect 5740 19908 5796 19918
rect 5068 17668 5124 17678
rect 5068 13972 5124 17612
rect 5404 16996 5460 17006
rect 5292 15540 5348 15550
rect 5292 14084 5348 15484
rect 5292 14018 5348 14028
rect 5068 13906 5124 13916
rect 4956 12964 5012 13468
rect 4956 12898 5012 12908
rect 4956 12404 5012 12414
rect 4956 10612 5012 12348
rect 4956 8484 5012 10556
rect 5404 10164 5460 16940
rect 5740 14868 5796 19852
rect 5740 14802 5796 14812
rect 5852 16772 5908 16782
rect 5852 13188 5908 16716
rect 5852 13122 5908 13132
rect 6188 14532 6244 23492
rect 6412 22372 6468 24108
rect 6524 23940 6580 23950
rect 6748 23940 6804 23950
rect 6580 23884 6748 23940
rect 6524 23874 6580 23884
rect 6748 23604 6804 23884
rect 6748 23538 6804 23548
rect 6412 17108 6468 22316
rect 6412 15540 6468 17052
rect 6412 15474 6468 15484
rect 6636 18564 6692 18574
rect 6188 12852 6244 14476
rect 6524 14980 6580 14990
rect 6524 13860 6580 14924
rect 6524 13794 6580 13804
rect 6188 12786 6244 12796
rect 6636 13748 6692 18508
rect 6860 16996 6916 27020
rect 6972 26740 7028 26750
rect 6972 21364 7028 26684
rect 7084 23716 7140 28364
rect 7196 26292 7252 29260
rect 7308 28756 7364 29372
rect 7308 28690 7364 28700
rect 7420 29092 7476 34076
rect 8652 32452 8708 32462
rect 8428 32116 8484 32126
rect 7420 27860 7476 29036
rect 7420 27794 7476 27804
rect 7756 30436 7812 30446
rect 7196 26226 7252 26236
rect 7644 25956 7700 25966
rect 7196 25620 7252 25630
rect 7196 23940 7252 25564
rect 7644 25396 7700 25900
rect 7420 25172 7476 25182
rect 7308 25060 7364 25070
rect 7308 24836 7364 25004
rect 7308 24770 7364 24780
rect 7196 23874 7252 23884
rect 7420 23940 7476 25116
rect 7420 23874 7476 23884
rect 7532 24836 7588 24846
rect 7532 23716 7588 24780
rect 7084 23660 7364 23716
rect 7308 23548 7364 23660
rect 7532 23650 7588 23660
rect 6972 21298 7028 21308
rect 7084 23492 7364 23548
rect 7420 23492 7476 23502
rect 6860 16930 6916 16940
rect 6860 15428 6916 15438
rect 6860 14084 6916 15372
rect 6972 14532 7028 14542
rect 7084 14532 7140 23492
rect 7420 22932 7476 23436
rect 7420 22866 7476 22876
rect 7028 14476 7140 14532
rect 7196 18116 7252 18126
rect 6972 14466 7028 14476
rect 6860 14018 6916 14028
rect 5404 10098 5460 10108
rect 6636 9492 6692 13692
rect 7196 12964 7252 18060
rect 7196 12898 7252 12908
rect 7308 17220 7364 17230
rect 7308 12068 7364 17164
rect 7308 12002 7364 12012
rect 7420 16660 7476 16670
rect 7420 15092 7476 16604
rect 7532 16548 7588 16558
rect 7532 15876 7588 16492
rect 7532 15810 7588 15820
rect 7420 10836 7476 15036
rect 7644 14644 7700 25340
rect 7644 14578 7700 14588
rect 7420 10770 7476 10780
rect 7644 13860 7700 13870
rect 7644 10612 7700 13804
rect 7756 13076 7812 30380
rect 8428 28868 8484 32060
rect 8652 29988 8708 32396
rect 8652 29764 8708 29932
rect 8652 29698 8708 29708
rect 8316 27748 8372 27758
rect 8092 26964 8148 26974
rect 7868 26852 7924 26862
rect 7868 25956 7924 26796
rect 8092 26628 8148 26908
rect 8092 26562 8148 26572
rect 7868 25890 7924 25900
rect 8316 21812 8372 27692
rect 8428 27412 8484 28812
rect 9772 28308 9828 34412
rect 14812 34020 14868 34030
rect 11788 33796 11844 33806
rect 12236 33796 12292 33806
rect 11844 33740 12236 33796
rect 11788 33730 11844 33740
rect 12236 33730 12292 33740
rect 9772 28242 9828 28252
rect 10668 30884 10724 30894
rect 8428 27346 8484 27356
rect 10668 26628 10724 30828
rect 11788 30772 11844 30782
rect 11788 27748 11844 30716
rect 11788 27682 11844 27692
rect 14476 29876 14532 29886
rect 14028 27524 14084 27534
rect 9660 25620 9716 25630
rect 8316 21746 8372 21756
rect 9324 25508 9380 25518
rect 9324 24500 9380 25452
rect 7980 21588 8036 21598
rect 7980 14308 8036 21532
rect 8204 17780 8260 17790
rect 8204 16660 8260 17724
rect 8204 16594 8260 16604
rect 8316 17668 8372 17678
rect 7980 14242 8036 14252
rect 8092 15764 8148 15774
rect 7756 13010 7812 13020
rect 8092 13076 8148 15708
rect 8316 15148 8372 17612
rect 8092 13010 8148 13020
rect 8204 15092 8372 15148
rect 8204 13748 8260 15092
rect 8540 14868 8596 14878
rect 8540 14644 8596 14812
rect 8652 14644 8708 14654
rect 8540 14588 8652 14644
rect 8652 14578 8708 14588
rect 8876 14532 8932 14542
rect 8652 13860 8708 13870
rect 8876 13860 8932 14476
rect 8708 13804 8932 13860
rect 8652 13794 8708 13804
rect 8204 11620 8260 13692
rect 9324 12740 9380 24444
rect 9660 17780 9716 25564
rect 9772 24836 9828 24846
rect 9772 23828 9828 24780
rect 9772 23762 9828 23772
rect 9996 24500 10052 24510
rect 9996 23604 10052 24444
rect 10668 23940 10724 26572
rect 13804 27188 13860 27198
rect 13804 26964 13860 27132
rect 11788 26180 11844 26190
rect 10668 23874 10724 23884
rect 11676 23940 11732 23950
rect 9996 23538 10052 23548
rect 9660 17556 9716 17724
rect 9660 17490 9716 17500
rect 10332 19348 10388 19358
rect 10220 15652 10276 15662
rect 9324 12674 9380 12684
rect 9660 15428 9716 15438
rect 9660 14756 9716 15372
rect 8204 11554 8260 11564
rect 8316 11732 8372 11742
rect 7644 10546 7700 10556
rect 8316 11284 8372 11676
rect 6636 9426 6692 9436
rect 4956 8418 5012 8428
rect 5628 8932 5684 8942
rect 5628 6244 5684 8876
rect 5628 6178 5684 6188
rect 8316 3220 8372 11228
rect 9660 5796 9716 14700
rect 9660 5236 9716 5740
rect 9660 5170 9716 5180
rect 10108 12740 10164 12750
rect 10108 12068 10164 12684
rect 10108 4564 10164 12012
rect 10108 4498 10164 4508
rect 10220 9268 10276 15596
rect 10332 14084 10388 19292
rect 11676 18788 11732 23884
rect 11676 18004 11732 18732
rect 11676 15316 11732 17948
rect 11788 16324 11844 26124
rect 12236 26180 12292 26190
rect 12236 25844 12292 26124
rect 13804 25956 13860 26908
rect 13804 25890 13860 25900
rect 11900 25508 11956 25518
rect 11900 24948 11956 25452
rect 11900 24882 11956 24892
rect 11900 22932 11956 22942
rect 11900 17108 11956 22876
rect 12124 18788 12180 18798
rect 12124 18564 12180 18732
rect 12124 18498 12180 18508
rect 11900 17042 11956 17052
rect 11788 16258 11844 16268
rect 10332 14018 10388 14028
rect 11564 14308 11620 14318
rect 10220 3780 10276 9212
rect 10556 10052 10612 10062
rect 10556 5236 10612 9996
rect 10556 5170 10612 5180
rect 11564 5236 11620 14252
rect 11676 9268 11732 15260
rect 11900 15092 11956 15102
rect 12236 15092 12292 25788
rect 14028 25396 14084 27468
rect 14364 27524 14420 27534
rect 14252 27300 14308 27310
rect 14364 27300 14420 27468
rect 14308 27244 14420 27300
rect 14252 27234 14308 27244
rect 14028 25330 14084 25340
rect 12348 24276 12404 24286
rect 12348 18788 12404 24220
rect 14476 23716 14532 29820
rect 14812 24276 14868 33964
rect 14924 33572 14980 39116
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 15148 38612 15204 38622
rect 15148 36708 15204 38556
rect 16604 38276 16660 38286
rect 16604 38052 16660 38220
rect 16604 37986 16660 37996
rect 15148 36642 15204 36652
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 14924 33506 14980 33516
rect 16716 35700 16772 35710
rect 14812 24210 14868 24220
rect 15036 31444 15092 31454
rect 14476 23650 14532 23660
rect 15036 23604 15092 31388
rect 16604 28980 16660 28990
rect 15260 24724 15316 24734
rect 15036 23538 15092 23548
rect 15148 24164 15204 24174
rect 13468 23380 13524 23390
rect 12348 18722 12404 18732
rect 13244 22036 13300 22046
rect 11956 15036 12292 15092
rect 11900 15026 11956 15036
rect 11676 9202 11732 9212
rect 12236 8484 12292 15036
rect 12460 18676 12516 18686
rect 12460 11844 12516 18620
rect 13244 18228 13300 21980
rect 13244 16884 13300 18172
rect 13356 21588 13412 21598
rect 13356 19460 13412 21532
rect 13356 18004 13412 19404
rect 13468 18228 13524 23324
rect 15036 22484 15092 22494
rect 15148 22484 15204 24108
rect 15092 22428 15204 22484
rect 15036 22418 15092 22428
rect 13580 19908 13636 19918
rect 13580 19460 13636 19852
rect 13580 19394 13636 19404
rect 13916 19908 13972 19918
rect 13468 18162 13524 18172
rect 13692 19236 13748 19246
rect 13356 17938 13412 17948
rect 13244 16818 13300 16828
rect 13468 17668 13524 17678
rect 13468 13636 13524 17612
rect 13468 13570 13524 13580
rect 12460 11778 12516 11788
rect 12236 8418 12292 8428
rect 13692 9268 13748 19180
rect 13916 14644 13972 19852
rect 15260 19236 15316 24668
rect 15596 23716 15652 23726
rect 15260 19170 15316 19180
rect 15372 22708 15428 22718
rect 13916 10276 13972 14588
rect 15148 19124 15204 19134
rect 15036 12852 15092 12862
rect 14924 11620 14980 11630
rect 14924 11396 14980 11564
rect 14924 11330 14980 11340
rect 13916 10210 13972 10220
rect 11564 5170 11620 5180
rect 10220 3714 10276 3724
rect 8316 3154 8372 3164
rect 4844 1586 4900 1596
rect 13692 1652 13748 9212
rect 14812 9492 14868 9502
rect 14812 8932 14868 9436
rect 14812 8866 14868 8876
rect 15036 6916 15092 12796
rect 15148 12404 15204 19068
rect 15372 16660 15428 22652
rect 15372 16594 15428 16604
rect 15596 14084 15652 23660
rect 16492 23044 16548 23054
rect 16492 22372 16548 22988
rect 16492 22306 16548 22316
rect 16604 21476 16660 28924
rect 16716 24724 16772 35644
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 17500 32340 17556 32350
rect 17276 32116 17332 32126
rect 17276 25508 17332 32060
rect 17500 25956 17556 32284
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 18620 30324 18676 30334
rect 18620 26852 18676 30268
rect 18620 26786 18676 26796
rect 18732 30100 18788 30110
rect 17500 25890 17556 25900
rect 17724 26180 17780 26190
rect 16716 24658 16772 24668
rect 17052 25396 17108 25406
rect 16604 21410 16660 21420
rect 16940 24052 16996 24062
rect 16716 20468 16772 20478
rect 15820 19572 15876 19582
rect 15708 18676 15764 18686
rect 15708 18228 15764 18620
rect 15708 18162 15764 18172
rect 15820 18564 15876 19516
rect 15596 14018 15652 14028
rect 15148 9268 15204 12348
rect 15148 9202 15204 9212
rect 15820 12740 15876 18508
rect 16268 17780 16324 17790
rect 16268 16772 16324 17724
rect 16156 16660 16212 16670
rect 16044 16324 16100 16334
rect 15036 6850 15092 6860
rect 15820 2996 15876 12684
rect 15932 13972 15988 13982
rect 15932 9940 15988 13916
rect 15932 9380 15988 9884
rect 15932 9314 15988 9324
rect 16044 8372 16100 16268
rect 16156 9268 16212 16604
rect 16268 12740 16324 16716
rect 16716 15652 16772 20412
rect 16940 18452 16996 23996
rect 16940 18386 16996 18396
rect 16716 15586 16772 15596
rect 16828 18116 16884 18126
rect 16604 14532 16660 14542
rect 16380 13972 16436 13982
rect 16380 13076 16436 13916
rect 16380 13010 16436 13020
rect 16268 12674 16324 12684
rect 16604 11732 16660 14476
rect 16828 12404 16884 18060
rect 16828 12338 16884 12348
rect 17052 13636 17108 25340
rect 17164 19012 17220 19022
rect 17164 17892 17220 18956
rect 17164 17826 17220 17836
rect 17052 12068 17108 13580
rect 17052 12002 17108 12012
rect 16604 11666 16660 11676
rect 16828 11732 16884 11742
rect 16604 11396 16660 11406
rect 16828 11396 16884 11676
rect 16660 11340 16884 11396
rect 16604 11330 16660 11340
rect 16156 9202 16212 9212
rect 16604 9380 16660 9390
rect 16044 8306 16100 8316
rect 16604 3220 16660 9324
rect 17276 6804 17332 25452
rect 17724 23044 17780 26124
rect 18732 24724 18788 30044
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19628 29204 19684 29214
rect 19404 28084 19460 28094
rect 19180 25620 19236 25630
rect 18732 24658 18788 24668
rect 19068 25564 19180 25620
rect 19068 24276 19124 25564
rect 19180 25554 19236 25564
rect 17724 22484 17780 22988
rect 18956 23492 19012 23502
rect 17724 10500 17780 22428
rect 18732 22484 18788 22494
rect 18508 22148 18564 22158
rect 18508 21700 18564 22092
rect 18732 21812 18788 22428
rect 18732 21746 18788 21756
rect 18396 21140 18452 21150
rect 18172 19012 18228 19022
rect 18172 18788 18228 18956
rect 18172 15540 18228 18732
rect 18396 17556 18452 21084
rect 18396 17490 18452 17500
rect 18508 18900 18564 21644
rect 18172 12180 18228 15484
rect 18508 12628 18564 18844
rect 18732 21476 18788 21486
rect 18732 16100 18788 21420
rect 18956 19796 19012 23436
rect 19068 20020 19124 24220
rect 19180 24948 19236 24958
rect 19180 22596 19236 24892
rect 19180 22036 19236 22540
rect 19180 21970 19236 21980
rect 19404 20244 19460 28028
rect 19516 25844 19572 25854
rect 19516 24500 19572 25788
rect 19516 24434 19572 24444
rect 19404 20178 19460 20188
rect 19516 23380 19572 23390
rect 19068 19954 19124 19964
rect 19292 20020 19348 20030
rect 19292 19796 19348 19964
rect 18956 19740 19348 19796
rect 18956 18452 19012 19740
rect 18620 16044 18732 16100
rect 18620 14644 18676 16044
rect 18732 16034 18788 16044
rect 18844 17892 18900 17902
rect 18844 16884 18900 17836
rect 18956 17332 19012 18396
rect 19180 18452 19236 18462
rect 18956 17266 19012 17276
rect 19068 18116 19124 18126
rect 18620 14578 18676 14588
rect 18732 15652 18788 15662
rect 18732 13636 18788 15596
rect 18844 15428 18900 16828
rect 18844 15362 18900 15372
rect 19068 15092 19124 18060
rect 19068 14084 19124 15036
rect 19068 14018 19124 14028
rect 19180 18004 19236 18396
rect 19180 13860 19236 17948
rect 19516 17892 19572 23324
rect 19628 19348 19684 29148
rect 19628 19282 19684 19292
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19516 17826 19572 17836
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19628 16884 19684 16894
rect 19180 13794 19236 13804
rect 19404 15876 19460 15886
rect 18732 13570 18788 13580
rect 18508 12562 18564 12572
rect 18956 13188 19012 13198
rect 18956 12516 19012 13132
rect 18956 12450 19012 12460
rect 19404 12852 19460 15820
rect 19404 12516 19460 12796
rect 19404 12450 19460 12460
rect 19516 15428 19572 15438
rect 18172 12114 18228 12124
rect 17724 10434 17780 10444
rect 17276 6738 17332 6748
rect 19068 8820 19124 8830
rect 19068 5796 19124 8764
rect 19516 7700 19572 15372
rect 19628 13188 19684 16828
rect 19628 13122 19684 13132
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19628 12740 19684 12750
rect 19628 11844 19684 12684
rect 19628 11778 19684 11788
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19516 7634 19572 7644
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19068 5730 19124 5740
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 16604 3154 16660 3164
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 20188 46452 20244 46462
rect 20188 4676 20244 46396
rect 26124 43092 26180 43102
rect 25228 39396 25284 39406
rect 23100 28756 23156 28766
rect 22316 27972 22372 27982
rect 20300 23716 20356 23726
rect 20300 21364 20356 23660
rect 22316 21700 22372 27916
rect 22316 21634 22372 21644
rect 20300 21298 20356 21308
rect 22876 20580 22932 20590
rect 20748 20468 20804 20478
rect 20524 15652 20580 15662
rect 20300 15428 20356 15438
rect 20300 12964 20356 15372
rect 20300 10388 20356 12908
rect 20524 14532 20580 15596
rect 20524 12964 20580 14476
rect 20524 12898 20580 12908
rect 20748 11396 20804 20412
rect 22876 19012 22932 20524
rect 22876 18946 22932 18956
rect 21868 18340 21924 18350
rect 21868 18116 21924 18284
rect 21420 17556 21476 17566
rect 21420 14868 21476 17500
rect 21420 12740 21476 14812
rect 21868 13300 21924 18060
rect 23100 14644 23156 28700
rect 23436 28420 23492 28430
rect 23324 18676 23380 18686
rect 23324 17444 23380 18620
rect 23324 17378 23380 17388
rect 23436 16660 23492 28364
rect 24780 27412 24836 27422
rect 24332 22932 24388 22942
rect 23548 22820 23604 22830
rect 23548 19684 23604 22764
rect 24220 22036 24276 22046
rect 23548 18228 23604 19628
rect 23548 18162 23604 18172
rect 23772 21252 23828 21262
rect 23772 19684 23828 21196
rect 23436 16594 23492 16604
rect 23660 17780 23716 17790
rect 23548 16324 23604 16334
rect 23100 14578 23156 14588
rect 23324 15988 23380 15998
rect 21868 13234 21924 13244
rect 23324 14196 23380 15932
rect 23548 15540 23604 16268
rect 23548 15474 23604 15484
rect 23660 16212 23716 17724
rect 21420 12674 21476 12684
rect 23324 12740 23380 14140
rect 23436 15204 23492 15214
rect 23436 14308 23492 15148
rect 23436 13636 23492 14252
rect 23660 13972 23716 16156
rect 23772 15204 23828 19628
rect 24220 19012 24276 21980
rect 24332 21588 24388 22876
rect 24332 19908 24388 21532
rect 24444 21812 24500 21822
rect 24444 20244 24500 21756
rect 24444 20178 24500 20188
rect 24332 19842 24388 19852
rect 24220 18946 24276 18956
rect 24556 19572 24612 19582
rect 24556 16100 24612 19516
rect 24556 16034 24612 16044
rect 24780 15540 24836 27356
rect 25228 20916 25284 39340
rect 26124 26908 26180 43036
rect 26012 26852 26180 26908
rect 26236 27524 26292 27534
rect 26012 26180 26068 26852
rect 25340 25172 25396 25182
rect 25340 24276 25396 25116
rect 25340 24210 25396 24220
rect 25228 20850 25284 20860
rect 25900 22820 25956 22830
rect 25900 20356 25956 22764
rect 25900 20290 25956 20300
rect 25676 18340 25732 18350
rect 25228 16884 25284 16894
rect 25228 15988 25284 16828
rect 25228 15922 25284 15932
rect 24780 15474 24836 15484
rect 23772 15138 23828 15148
rect 23660 13906 23716 13916
rect 24220 13972 24276 13982
rect 23436 13570 23492 13580
rect 23324 12674 23380 12684
rect 24220 12180 24276 13916
rect 24220 12114 24276 12124
rect 20748 11330 20804 11340
rect 22764 11508 22820 11518
rect 20300 10322 20356 10332
rect 22764 6580 22820 11452
rect 22764 6514 22820 6524
rect 20188 4610 20244 4620
rect 22988 5236 23044 5246
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 15820 2930 15876 2940
rect 22988 2884 23044 5180
rect 25676 2996 25732 18284
rect 26012 18004 26068 26124
rect 26236 18676 26292 27468
rect 26460 22708 26516 22718
rect 26460 19348 26516 22652
rect 27020 22596 27076 22606
rect 26460 19282 26516 19292
rect 26572 22484 26628 22494
rect 26236 18610 26292 18620
rect 26460 19012 26516 19022
rect 26012 17938 26068 17948
rect 25676 2930 25732 2940
rect 26348 17108 26404 17118
rect 26348 13748 26404 17052
rect 26460 16100 26516 18956
rect 26460 16034 26516 16044
rect 26572 16660 26628 22428
rect 22988 2818 23044 2828
rect 15260 2772 15316 2782
rect 15708 2772 15764 2782
rect 15316 2716 15708 2772
rect 15260 2706 15316 2716
rect 15708 2706 15764 2716
rect 13692 1586 13748 1596
rect 26348 1652 26404 13692
rect 26348 1586 26404 1596
rect 26572 1540 26628 16604
rect 26684 17668 26740 17678
rect 26684 15764 26740 17612
rect 26684 15698 26740 15708
rect 27020 14644 27076 22540
rect 27020 14578 27076 14588
rect 27692 7924 27748 55916
rect 35168 55692 35488 56508
rect 35168 55636 35196 55692
rect 35252 55636 35300 55692
rect 35356 55636 35404 55692
rect 35460 55636 35488 55692
rect 35168 54124 35488 55636
rect 35168 54068 35196 54124
rect 35252 54068 35300 54124
rect 35356 54068 35404 54124
rect 35460 54068 35488 54124
rect 35168 52556 35488 54068
rect 35168 52500 35196 52556
rect 35252 52500 35300 52556
rect 35356 52500 35404 52556
rect 35460 52500 35488 52556
rect 35168 50988 35488 52500
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 34748 49924 34804 49934
rect 34748 48692 34804 49868
rect 34748 48626 34804 48636
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 34300 47012 34356 47022
rect 28140 45332 28196 45342
rect 28140 10612 28196 45276
rect 34188 44436 34244 44446
rect 34188 36036 34244 44380
rect 34300 38052 34356 46956
rect 34300 37986 34356 37996
rect 35168 46284 35488 47796
rect 50528 56476 50848 56508
rect 50528 56420 50556 56476
rect 50612 56420 50660 56476
rect 50716 56420 50764 56476
rect 50820 56420 50848 56476
rect 50528 54908 50848 56420
rect 50528 54852 50556 54908
rect 50612 54852 50660 54908
rect 50716 54852 50764 54908
rect 50820 54852 50848 54908
rect 50528 53340 50848 54852
rect 50528 53284 50556 53340
rect 50612 53284 50660 53340
rect 50716 53284 50764 53340
rect 50820 53284 50848 53340
rect 50528 51772 50848 53284
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 41692 46452 41748 46462
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 39452 45780 39508 45790
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35644 42532 35700 42542
rect 35644 41188 35700 42476
rect 35644 41122 35700 41132
rect 35756 41972 35812 41982
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 34188 35970 34244 35980
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 34972 35476 35028 35486
rect 29372 32788 29428 32798
rect 28476 26852 28532 26862
rect 28476 23156 28532 26796
rect 28476 23090 28532 23100
rect 29260 24612 29316 24622
rect 28812 22260 28868 22270
rect 28812 16436 28868 22204
rect 29260 21588 29316 24556
rect 29260 21522 29316 21532
rect 28812 16370 28868 16380
rect 28140 10546 28196 10556
rect 27692 7858 27748 7868
rect 29372 6804 29428 32732
rect 34076 32564 34132 32574
rect 29484 31220 29540 31230
rect 29484 11844 29540 31164
rect 29932 30436 29988 30446
rect 29820 20132 29876 20142
rect 29820 15316 29876 20076
rect 29932 16100 29988 30380
rect 33628 28308 33684 28318
rect 30940 27300 30996 27310
rect 30940 25172 30996 27244
rect 30940 25106 30996 25116
rect 33516 25284 33572 25294
rect 33404 23268 33460 23278
rect 32732 21812 32788 21822
rect 30044 21700 30100 21710
rect 30044 19460 30100 21644
rect 30044 19394 30100 19404
rect 31724 20020 31780 20030
rect 29932 16034 29988 16044
rect 30828 16100 30884 16110
rect 29820 15250 29876 15260
rect 30828 13076 30884 16044
rect 31724 15540 31780 19964
rect 31724 15474 31780 15484
rect 30828 13010 30884 13020
rect 29484 11778 29540 11788
rect 32732 8372 32788 21756
rect 33404 13972 33460 23212
rect 33516 22260 33572 25228
rect 33516 21252 33572 22204
rect 33516 21186 33572 21196
rect 33404 13906 33460 13916
rect 32732 8306 32788 8316
rect 29372 6738 29428 6748
rect 33628 5124 33684 28252
rect 34076 28084 34132 32508
rect 34076 28018 34132 28028
rect 34972 17556 35028 35420
rect 34972 17490 35028 17500
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35644 40180 35700 40190
rect 35756 40180 35812 41916
rect 35700 40124 35812 40180
rect 35644 33684 35700 40124
rect 38668 36708 38724 36718
rect 38556 36484 38612 36494
rect 38668 36484 38724 36652
rect 38612 36428 38724 36484
rect 38556 36418 38612 36428
rect 35644 33618 35700 33628
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 38780 31556 38836 31566
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35756 31444 35812 31454
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35644 25284 35700 25294
rect 35644 23716 35700 25228
rect 35756 24500 35812 31388
rect 38668 30660 38724 30670
rect 38444 30548 38500 30558
rect 36652 30100 36708 30110
rect 36540 29316 36596 29326
rect 36540 28756 36596 29260
rect 36540 28690 36596 28700
rect 36428 27188 36484 27198
rect 36428 26292 36484 27132
rect 36428 26068 36484 26236
rect 36428 26002 36484 26012
rect 35756 24434 35812 24444
rect 35644 21028 35700 23660
rect 36652 23604 36708 30044
rect 38444 28196 38500 30492
rect 38444 28130 38500 28140
rect 37212 27188 37268 27198
rect 36764 26404 36820 26414
rect 36764 25172 36820 26348
rect 36764 25106 36820 25116
rect 37212 25172 37268 27132
rect 37212 25106 37268 25116
rect 38332 26964 38388 26974
rect 36652 23538 36708 23548
rect 36876 24612 36932 24622
rect 35644 20962 35700 20972
rect 35980 21812 36036 21822
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 33628 5058 33684 5068
rect 35168 16492 35488 18004
rect 35756 20468 35812 20478
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35644 17444 35700 17454
rect 35644 15652 35700 17388
rect 35644 15586 35700 15596
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35756 10836 35812 20412
rect 35980 17108 36036 21756
rect 36876 20468 36932 24556
rect 38108 23716 38164 23726
rect 36988 23604 37044 23614
rect 36988 22708 37044 23548
rect 36988 22642 37044 22652
rect 37996 22260 38052 22270
rect 36876 18228 36932 20412
rect 37436 20580 37492 20590
rect 36876 18162 36932 18172
rect 37100 18788 37156 18798
rect 37100 18228 37156 18732
rect 37100 18162 37156 18172
rect 37436 17780 37492 20524
rect 37996 19908 38052 22204
rect 38108 22148 38164 23660
rect 38108 22082 38164 22092
rect 38332 23716 38388 26908
rect 37996 19842 38052 19852
rect 37436 17714 37492 17724
rect 35980 17042 36036 17052
rect 37100 15764 37156 15774
rect 37100 14980 37156 15708
rect 37100 14914 37156 14924
rect 35756 10770 35812 10780
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 28364 4340 28420 4350
rect 28364 3780 28420 4284
rect 28364 3714 28420 3724
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 38332 2660 38388 23660
rect 38444 22708 38500 22718
rect 38444 16548 38500 22652
rect 38556 22260 38612 22270
rect 38556 20692 38612 22204
rect 38556 20626 38612 20636
rect 38444 16482 38500 16492
rect 38668 19460 38724 30604
rect 38780 23716 38836 31500
rect 39116 29988 39172 29998
rect 39116 27300 39172 29932
rect 39116 26292 39172 27244
rect 39116 26226 39172 26236
rect 39228 28084 39284 28094
rect 39228 25060 39284 28028
rect 39228 24994 39284 25004
rect 38780 23650 38836 23660
rect 38668 15764 38724 19404
rect 38668 15698 38724 15708
rect 39004 21476 39060 21486
rect 39004 2996 39060 21420
rect 39116 18564 39172 18574
rect 39116 14644 39172 18508
rect 39116 14578 39172 14588
rect 39452 14532 39508 45724
rect 40012 43764 40068 43774
rect 40012 42308 40068 43708
rect 40012 42242 40068 42252
rect 41692 43204 41748 46396
rect 50316 46116 50372 46126
rect 41692 38500 41748 43148
rect 43372 43204 43428 43214
rect 43372 39732 43428 43148
rect 50316 41972 50372 46060
rect 50316 41906 50372 41916
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 53900 48244 53956 48254
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 43372 39666 43428 39676
rect 50528 40796 50848 42308
rect 52556 43652 52612 43662
rect 52556 43316 52612 43596
rect 52444 42084 52500 42094
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 42140 39620 42196 39630
rect 41692 38434 41748 38444
rect 42028 38948 42084 38958
rect 41468 37940 41524 37950
rect 40796 37716 40852 37726
rect 40460 32452 40516 32462
rect 40460 30212 40516 32396
rect 40348 27188 40404 27198
rect 40348 26628 40404 27132
rect 40348 26562 40404 26572
rect 40460 26516 40516 30156
rect 40572 28644 40628 28654
rect 40572 27972 40628 28588
rect 40572 27906 40628 27916
rect 40460 26450 40516 26460
rect 40684 26740 40740 26750
rect 40348 25508 40404 25518
rect 40348 23492 40404 25452
rect 40684 24052 40740 26684
rect 40684 23986 40740 23996
rect 40348 23426 40404 23436
rect 40124 23268 40180 23278
rect 40124 22932 40180 23212
rect 40124 22866 40180 22876
rect 40236 22484 40292 22494
rect 40012 22148 40068 22158
rect 40012 19572 40068 22092
rect 40012 16996 40068 19516
rect 40012 16930 40068 16940
rect 40236 19908 40292 22428
rect 40572 21924 40628 21934
rect 40572 21364 40628 21868
rect 39564 16212 39620 16222
rect 39564 15540 39620 16156
rect 39564 14980 39620 15484
rect 39564 14914 39620 14924
rect 39900 15876 39956 15886
rect 39452 12852 39508 14476
rect 39452 12786 39508 12796
rect 39004 2930 39060 2940
rect 38332 2594 38388 2604
rect 39900 1652 39956 15820
rect 40236 12964 40292 19852
rect 40348 21028 40404 21038
rect 40348 17892 40404 20972
rect 40348 17826 40404 17836
rect 40460 20692 40516 20702
rect 40460 15540 40516 20636
rect 40460 15474 40516 15484
rect 40572 16884 40628 21308
rect 40684 20356 40740 20366
rect 40684 18452 40740 20300
rect 40796 18900 40852 37660
rect 41468 37492 41524 37884
rect 40908 26852 40964 26862
rect 40908 24948 40964 26796
rect 41468 25508 41524 37436
rect 42028 37380 42084 38892
rect 42028 37314 42084 37324
rect 41692 29204 41748 29214
rect 41468 25442 41524 25452
rect 41580 26404 41636 26414
rect 40908 24882 40964 24892
rect 41020 25284 41076 25294
rect 40796 18834 40852 18844
rect 40908 20804 40964 20814
rect 40684 18386 40740 18396
rect 40908 18340 40964 20748
rect 41020 20020 41076 25228
rect 41020 19954 41076 19964
rect 41132 20916 41188 20926
rect 40908 18274 40964 18284
rect 40236 12898 40292 12908
rect 40572 12964 40628 16828
rect 41132 16884 41188 20860
rect 41132 16818 41188 16828
rect 41468 20804 41524 20814
rect 41468 20468 41524 20748
rect 41468 15148 41524 20412
rect 41580 17332 41636 26348
rect 41692 24052 41748 29148
rect 42140 26908 42196 39564
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 44380 37940 44436 37950
rect 43932 34244 43988 34254
rect 43036 32228 43092 32238
rect 42028 26852 42196 26908
rect 42252 30324 42308 30334
rect 41804 26180 41860 26190
rect 41804 25284 41860 26124
rect 41804 25218 41860 25228
rect 41692 23986 41748 23996
rect 41692 22708 41748 22718
rect 41692 22148 41748 22652
rect 41692 21924 41748 22092
rect 41692 21858 41748 21868
rect 41580 17266 41636 17276
rect 41804 17108 41860 17118
rect 41468 15092 41636 15148
rect 41580 13636 41636 15092
rect 41580 13570 41636 13580
rect 41692 14420 41748 14430
rect 41692 13300 41748 14364
rect 41692 13234 41748 13244
rect 40572 12898 40628 12908
rect 41804 11172 41860 17052
rect 42028 15204 42084 26852
rect 42252 26740 42308 30268
rect 42252 26674 42308 26684
rect 42588 26964 42644 26974
rect 42028 15138 42084 15148
rect 42140 26404 42196 26414
rect 41804 11106 41860 11116
rect 41916 13636 41972 13646
rect 41916 7812 41972 13580
rect 42140 13188 42196 26348
rect 42476 25284 42532 25294
rect 42476 23156 42532 25228
rect 42588 24164 42644 26908
rect 42588 23828 42644 24108
rect 43036 25284 43092 32172
rect 43596 30548 43652 30558
rect 43596 28644 43652 30492
rect 43596 28578 43652 28588
rect 43708 27524 43764 27534
rect 43372 27300 43428 27310
rect 43260 27076 43316 27086
rect 43260 26852 43316 27020
rect 43260 26786 43316 26796
rect 43372 26628 43428 27244
rect 43372 26562 43428 26572
rect 43596 27076 43652 27086
rect 42588 23762 42644 23772
rect 42700 24052 42756 24062
rect 42700 23492 42756 23996
rect 42700 23426 42756 23436
rect 43036 23380 43092 25228
rect 43596 25172 43652 27020
rect 43596 25106 43652 25116
rect 43484 24500 43540 24510
rect 43484 23548 43540 24444
rect 43036 23314 43092 23324
rect 43372 23492 43540 23548
rect 42476 23090 42532 23100
rect 42812 20804 42868 20814
rect 42812 19236 42868 20748
rect 42812 19170 42868 19180
rect 43372 19796 43428 23492
rect 43708 20916 43764 27468
rect 43596 20860 43708 20916
rect 42140 13122 42196 13132
rect 43036 18452 43092 18462
rect 43036 17108 43092 18396
rect 43036 11508 43092 17052
rect 43372 16660 43428 19740
rect 43484 20244 43540 20254
rect 43484 18676 43540 20188
rect 43484 18610 43540 18620
rect 43596 17780 43652 20860
rect 43708 20850 43764 20860
rect 43820 23044 43876 23054
rect 43820 18004 43876 22988
rect 43932 20580 43988 34188
rect 44156 33684 44212 33694
rect 44044 29876 44100 29886
rect 44044 26516 44100 29820
rect 44156 28980 44212 33628
rect 44156 28914 44212 28924
rect 44044 26450 44100 26460
rect 44156 24724 44212 24734
rect 44156 21812 44212 24668
rect 44156 21746 44212 21756
rect 43932 20514 43988 20524
rect 44044 21588 44100 21598
rect 43820 17938 43876 17948
rect 44044 19572 44100 21532
rect 43596 17714 43652 17724
rect 44044 17556 44100 19516
rect 44044 17490 44100 17500
rect 44156 21028 44212 21038
rect 43372 16594 43428 16604
rect 43596 16996 43652 17006
rect 43596 15148 43652 16940
rect 43820 16660 43876 16670
rect 43036 11442 43092 11452
rect 43484 15092 43652 15148
rect 43708 15428 43764 15438
rect 43484 9828 43540 15092
rect 43708 14980 43764 15372
rect 43596 14924 43764 14980
rect 43596 10948 43652 14924
rect 43820 13524 43876 16604
rect 43820 13458 43876 13468
rect 43932 16100 43988 16110
rect 43932 12516 43988 16044
rect 44156 15988 44212 20972
rect 44268 20020 44324 20030
rect 44268 17444 44324 19964
rect 44268 17378 44324 17388
rect 44156 13972 44212 15932
rect 44380 15540 44436 37884
rect 50528 37660 50848 39172
rect 52332 41524 52388 41534
rect 51996 38948 52052 38958
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 47180 35588 47236 35598
rect 44492 34804 44548 34814
rect 44492 32452 44548 34748
rect 44492 32386 44548 32396
rect 44940 34020 44996 34030
rect 44492 29428 44548 29438
rect 44492 25732 44548 29372
rect 44604 26516 44660 26526
rect 44604 26068 44660 26460
rect 44604 26002 44660 26012
rect 44492 25666 44548 25676
rect 44940 25508 44996 33964
rect 44940 25442 44996 25452
rect 45948 33460 46004 33470
rect 45836 21028 45892 21038
rect 45612 20916 45668 20926
rect 45612 20468 45668 20860
rect 45612 20402 45668 20412
rect 45836 17668 45892 20972
rect 45948 19348 46004 33404
rect 47180 32900 47236 35532
rect 48972 34804 49028 34814
rect 46844 31780 46900 31790
rect 46732 29092 46788 29102
rect 46732 24836 46788 29036
rect 46844 26964 46900 31724
rect 47180 29652 47236 32844
rect 47852 34692 47908 34702
rect 47180 29586 47236 29596
rect 47516 32564 47572 32574
rect 46844 26898 46900 26908
rect 46732 24770 46788 24780
rect 46956 25172 47012 25182
rect 45948 19282 46004 19292
rect 46620 22260 46676 22270
rect 46620 21252 46676 22204
rect 45836 17602 45892 17612
rect 46172 17556 46228 17566
rect 44380 15474 44436 15484
rect 45276 17444 45332 17454
rect 44156 13906 44212 13916
rect 45276 13972 45332 17388
rect 45276 13906 45332 13916
rect 43932 12450 43988 12460
rect 46172 12516 46228 17500
rect 46396 17332 46452 17342
rect 46284 15652 46340 15662
rect 46284 15092 46340 15596
rect 46284 15026 46340 15036
rect 46396 13972 46452 17276
rect 46396 13906 46452 13916
rect 46508 15540 46564 15550
rect 46172 12450 46228 12460
rect 46508 11060 46564 15484
rect 46620 14196 46676 21196
rect 46956 20916 47012 25116
rect 47404 23156 47460 23166
rect 46956 20850 47012 20860
rect 47068 22932 47124 22942
rect 47068 21252 47124 22876
rect 47404 21812 47460 23100
rect 47404 21746 47460 21756
rect 47516 21588 47572 32508
rect 47852 26852 47908 34636
rect 47852 26786 47908 26796
rect 48076 33236 48132 33246
rect 47516 21522 47572 21532
rect 47740 26404 47796 26414
rect 46844 17668 46900 17678
rect 46844 16212 46900 17612
rect 46844 15316 46900 16156
rect 46844 15250 46900 15260
rect 46620 14130 46676 14140
rect 47068 13636 47124 21196
rect 47404 20692 47460 20702
rect 47404 19236 47460 20636
rect 47404 18564 47460 19180
rect 47404 18498 47460 18508
rect 47068 13570 47124 13580
rect 47180 17780 47236 17790
rect 47180 11956 47236 17724
rect 47180 11890 47236 11900
rect 47740 15652 47796 26348
rect 48076 25508 48132 33180
rect 48636 32116 48692 32126
rect 48636 31892 48692 32060
rect 48636 28644 48692 31836
rect 48860 31780 48916 31790
rect 48636 28578 48692 28588
rect 48748 29652 48804 29662
rect 48524 27412 48580 27422
rect 48524 27076 48580 27356
rect 48076 25442 48132 25452
rect 48412 25508 48468 25518
rect 48188 24948 48244 24958
rect 48188 23940 48244 24892
rect 48188 23874 48244 23884
rect 48076 23716 48132 23726
rect 47740 15204 47796 15596
rect 46508 10994 46564 11004
rect 43596 10882 43652 10892
rect 43484 9762 43540 9772
rect 41916 7746 41972 7756
rect 47740 6580 47796 15148
rect 47852 23604 47908 23614
rect 47852 21700 47908 23548
rect 47964 21700 48020 21710
rect 47852 21644 47964 21700
rect 47852 14644 47908 21644
rect 47964 21634 48020 21644
rect 47852 14578 47908 14588
rect 47964 18228 48020 18238
rect 47964 17108 48020 18172
rect 47964 7700 48020 17052
rect 48076 11620 48132 23660
rect 48188 21924 48244 21934
rect 48188 21476 48244 21868
rect 48188 21410 48244 21420
rect 48300 21812 48356 21822
rect 48300 21588 48356 21756
rect 48076 11554 48132 11564
rect 48300 20692 48356 21532
rect 48300 9268 48356 20636
rect 48412 14756 48468 25452
rect 48524 23380 48580 27020
rect 48748 25732 48804 29596
rect 48636 24500 48692 24510
rect 48636 23716 48692 24444
rect 48636 23650 48692 23660
rect 48524 23314 48580 23324
rect 48636 22372 48692 22382
rect 48524 22260 48580 22270
rect 48524 18004 48580 22204
rect 48636 21476 48692 22316
rect 48636 21410 48692 21420
rect 48636 20580 48692 20590
rect 48636 18228 48692 20524
rect 48748 20468 48804 25676
rect 48860 28756 48916 31724
rect 48860 24724 48916 28700
rect 48860 24658 48916 24668
rect 48748 20402 48804 20412
rect 48860 20580 48916 20590
rect 48636 18162 48692 18172
rect 48524 17948 48692 18004
rect 48524 15316 48580 15326
rect 48524 14980 48580 15260
rect 48524 14914 48580 14924
rect 48412 14690 48468 14700
rect 48636 14420 48692 17948
rect 48636 14354 48692 14364
rect 48748 16436 48804 16446
rect 48748 12404 48804 16380
rect 48748 12338 48804 12348
rect 48860 10052 48916 20524
rect 48972 19348 49028 34748
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 49980 33012 50036 33022
rect 49644 32116 49700 32126
rect 49644 29092 49700 32060
rect 49980 31668 50036 32956
rect 50528 32956 50848 34468
rect 50988 37828 51044 37838
rect 50988 33348 51044 37772
rect 50988 33282 51044 33292
rect 51100 37716 51156 37726
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 49980 31602 50036 31612
rect 50204 32564 50260 32574
rect 49980 30660 50036 30670
rect 49980 29204 50036 30604
rect 49644 29026 49700 29036
rect 49868 29092 49924 29102
rect 49644 28532 49700 28542
rect 49420 28196 49476 28206
rect 49308 27748 49364 27758
rect 49084 26628 49140 26638
rect 49084 26068 49140 26572
rect 49084 26002 49140 26012
rect 49308 24052 49364 27692
rect 49308 23828 49364 23996
rect 49308 23762 49364 23772
rect 49420 24164 49476 28140
rect 49532 26740 49588 26750
rect 49532 25396 49588 26684
rect 49532 25330 49588 25340
rect 49532 24164 49588 24174
rect 49420 24108 49532 24164
rect 48972 19282 49028 19292
rect 49084 23492 49140 23502
rect 49084 17332 49140 23436
rect 49308 23044 49364 23054
rect 49308 22260 49364 22988
rect 49308 22194 49364 22204
rect 49308 21588 49364 21598
rect 49308 18788 49364 21532
rect 49420 20132 49476 24108
rect 49532 24098 49588 24108
rect 49644 23492 49700 28476
rect 49532 23436 49700 23492
rect 49532 23268 49588 23436
rect 49532 23212 49700 23268
rect 49532 23044 49588 23054
rect 49532 21364 49588 22988
rect 49644 22932 49700 23212
rect 49644 22866 49700 22876
rect 49756 22596 49812 22606
rect 49756 22148 49812 22540
rect 49756 22082 49812 22092
rect 49644 21364 49700 21374
rect 49532 21308 49644 21364
rect 49644 21298 49700 21308
rect 49420 20066 49476 20076
rect 49756 21028 49812 21038
rect 49308 18722 49364 18732
rect 49532 19796 49588 19806
rect 49532 18452 49588 19740
rect 49532 18386 49588 18396
rect 49644 19460 49700 19470
rect 49644 17668 49700 19404
rect 49756 18788 49812 20972
rect 49756 18722 49812 18732
rect 49644 17602 49700 17612
rect 49084 17266 49140 17276
rect 49644 16100 49700 16110
rect 49532 14308 49588 14318
rect 49532 12628 49588 14252
rect 49644 14196 49700 16044
rect 49644 12852 49700 14140
rect 49644 12786 49700 12796
rect 49756 15764 49812 15774
rect 49756 15204 49812 15708
rect 49532 11844 49588 12572
rect 49756 12628 49812 15148
rect 49868 14644 49924 29036
rect 49980 20580 50036 29148
rect 50204 27524 50260 32508
rect 50528 31388 50848 32900
rect 50316 31332 50372 31342
rect 50316 30446 50372 31276
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50316 30436 50428 30446
rect 50316 30380 50372 30436
rect 50372 30360 50428 30380
rect 50204 27458 50260 27468
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50204 26852 50260 26862
rect 50204 23716 50260 26796
rect 50528 26684 50848 28196
rect 51100 26908 51156 37660
rect 51212 37156 51268 37166
rect 51212 33572 51268 37100
rect 51996 35364 52052 38892
rect 51996 35298 52052 35308
rect 51212 33236 51268 33516
rect 51212 33170 51268 33180
rect 52108 32004 52164 32014
rect 51212 31780 51268 31790
rect 51212 31556 51268 31724
rect 51212 31490 51268 31500
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50204 23650 50260 23660
rect 50316 26404 50372 26414
rect 50204 23492 50260 23502
rect 50092 23436 50204 23492
rect 50092 23044 50148 23436
rect 50204 23426 50260 23436
rect 50092 22978 50148 22988
rect 50204 23156 50260 23166
rect 49980 20514 50036 20524
rect 50092 22148 50148 22158
rect 50092 18004 50148 22092
rect 50204 21588 50260 23100
rect 50204 21522 50260 21532
rect 50316 20356 50372 26348
rect 50092 17938 50148 17948
rect 50204 20020 50260 20030
rect 49868 14578 49924 14588
rect 49980 17108 50036 17118
rect 49756 12562 49812 12572
rect 49532 11778 49588 11788
rect 48860 9986 48916 9996
rect 48300 9202 48356 9212
rect 49980 8260 50036 17052
rect 50204 13412 50260 19964
rect 50204 13346 50260 13356
rect 50316 16996 50372 20300
rect 50316 12292 50372 16940
rect 50316 12226 50372 12236
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50988 26852 51156 26908
rect 51436 31332 51492 31342
rect 51436 29204 51492 31276
rect 50988 15204 51044 26852
rect 51100 26292 51156 26302
rect 51100 21924 51156 26236
rect 51324 25956 51380 25966
rect 51100 21858 51156 21868
rect 51212 24948 51268 24958
rect 51212 22148 51268 24892
rect 50988 15138 51044 15148
rect 51100 20916 51156 20926
rect 51100 18340 51156 20860
rect 51212 20244 51268 22092
rect 51212 20178 51268 20188
rect 51324 24276 51380 25900
rect 51324 23716 51380 24220
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 51100 15092 51156 18284
rect 51324 16436 51380 23660
rect 51436 22596 51492 29148
rect 51548 26964 51604 26974
rect 51548 26740 51604 26908
rect 51548 26674 51604 26684
rect 52108 25620 52164 31948
rect 52332 27188 52388 41468
rect 52444 40180 52500 42028
rect 52556 40628 52612 43260
rect 53340 43428 53396 43438
rect 52556 40562 52612 40572
rect 53116 40628 53172 40638
rect 52444 40114 52500 40124
rect 53116 31220 53172 40572
rect 53228 40404 53284 40414
rect 53228 35588 53284 40348
rect 53228 35522 53284 35532
rect 53340 36484 53396 43372
rect 53788 41076 53844 41086
rect 53564 39172 53620 39182
rect 53564 38668 53620 39116
rect 53788 38668 53844 41020
rect 53900 39956 53956 48188
rect 55804 46564 55860 46574
rect 55580 44996 55636 45006
rect 55468 44884 55524 44894
rect 54236 44548 54292 44558
rect 53900 39890 53956 39900
rect 54012 42196 54068 42206
rect 53564 38612 53732 38668
rect 53788 38612 53956 38668
rect 53564 38388 53620 38398
rect 53340 36260 53396 36428
rect 53340 34804 53396 36204
rect 53340 34738 53396 34748
rect 53452 38164 53508 38174
rect 53452 32788 53508 38108
rect 53564 33236 53620 38332
rect 53564 33170 53620 33180
rect 53508 32732 53620 32788
rect 53452 32722 53508 32732
rect 53116 31154 53172 31164
rect 53452 31444 53508 31454
rect 52332 27122 52388 27132
rect 52668 28420 52724 28430
rect 52668 27412 52724 28364
rect 52108 25554 52164 25564
rect 52220 26852 52276 26862
rect 52220 26068 52276 26796
rect 51436 22530 51492 22540
rect 51884 24612 51940 24622
rect 51436 22372 51492 22382
rect 51436 21364 51492 22316
rect 51436 21298 51492 21308
rect 51660 22036 51716 22046
rect 51660 20020 51716 21980
rect 51884 20804 51940 24556
rect 51884 20738 51940 20748
rect 51996 22036 52052 22046
rect 51660 19954 51716 19964
rect 51884 20244 51940 20254
rect 51324 16370 51380 16380
rect 51548 19796 51604 19806
rect 51100 13972 51156 15036
rect 51100 13906 51156 13916
rect 51436 16324 51492 16334
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50316 11732 50372 11742
rect 50316 8932 50372 11676
rect 50316 8866 50372 8876
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 49980 8194 50036 8204
rect 47964 7634 48020 7644
rect 50528 7868 50848 9380
rect 51100 13300 51156 13310
rect 51100 12964 51156 13244
rect 51100 9044 51156 12908
rect 51100 8978 51156 8988
rect 51436 8260 51492 16268
rect 51548 10164 51604 19740
rect 51548 10098 51604 10108
rect 51884 16548 51940 20188
rect 51996 19796 52052 21980
rect 51996 19730 52052 19740
rect 52108 18788 52164 18798
rect 52108 18452 52164 18732
rect 52108 18386 52164 18396
rect 52220 18228 52276 26012
rect 52444 24164 52500 24174
rect 52444 23268 52500 24108
rect 52444 23202 52500 23212
rect 52220 18162 52276 18172
rect 52332 22932 52388 22942
rect 52108 18004 52164 18014
rect 52108 17780 52164 17948
rect 52108 17714 52164 17724
rect 52332 17780 52388 22876
rect 52556 22372 52612 22382
rect 52444 18900 52500 18910
rect 52444 18004 52500 18844
rect 52444 17938 52500 17948
rect 52332 17714 52388 17724
rect 51884 15540 51940 16492
rect 51884 9268 51940 15484
rect 51996 15764 52052 15774
rect 51996 13076 52052 15708
rect 51996 13010 52052 13020
rect 52108 13860 52164 13870
rect 52108 11620 52164 13804
rect 52556 12628 52612 22316
rect 52668 16548 52724 27356
rect 53116 24724 53172 24734
rect 53116 19460 53172 24668
rect 53228 23044 53284 23054
rect 53228 21700 53284 22988
rect 53228 21634 53284 21644
rect 53340 21476 53396 21486
rect 53116 19394 53172 19404
rect 53228 21252 53284 21262
rect 52668 15316 52724 16492
rect 52668 15250 52724 15260
rect 52892 18788 52948 18798
rect 52556 12562 52612 12572
rect 52108 11554 52164 11564
rect 51884 9202 51940 9212
rect 52892 8372 52948 18732
rect 53228 13860 53284 21196
rect 53340 14644 53396 21420
rect 53452 15652 53508 31388
rect 53564 27300 53620 32732
rect 53676 31668 53732 38612
rect 53788 37716 53844 37726
rect 53788 36932 53844 37660
rect 53788 36866 53844 36876
rect 53676 31444 53732 31612
rect 53676 31378 53732 31388
rect 53788 35924 53844 35934
rect 53564 27234 53620 27244
rect 53676 25508 53732 25518
rect 53676 21476 53732 25452
rect 53676 21410 53732 21420
rect 53452 15586 53508 15596
rect 53564 18228 53620 18238
rect 53564 17108 53620 18172
rect 53340 14578 53396 14588
rect 53228 13794 53284 13804
rect 53564 11508 53620 17052
rect 53676 15988 53732 15998
rect 53676 14532 53732 15932
rect 53676 14466 53732 14476
rect 53564 11442 53620 11452
rect 52892 8306 52948 8316
rect 51436 8194 51492 8204
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 47740 5460 47796 6524
rect 47740 5394 47796 5404
rect 50528 6300 50848 7812
rect 53788 7812 53844 35868
rect 53900 34580 53956 38612
rect 54012 35924 54068 42140
rect 54236 39732 54292 44492
rect 54236 39666 54292 39676
rect 54684 44212 54740 44222
rect 54684 38276 54740 44156
rect 54684 38210 54740 38220
rect 55468 44100 55524 44828
rect 54012 35858 54068 35868
rect 55468 36484 55524 44044
rect 53900 34514 53956 34524
rect 54012 32116 54068 32126
rect 53900 20804 53956 20814
rect 53900 13636 53956 20748
rect 54012 19460 54068 32060
rect 55356 31220 55412 31230
rect 54348 28308 54404 28318
rect 54236 27636 54292 27646
rect 54236 26964 54292 27580
rect 54348 27524 54404 28252
rect 54348 27188 54404 27468
rect 54348 27122 54404 27132
rect 54236 26898 54292 26908
rect 54908 26964 54964 26974
rect 54796 26292 54852 26302
rect 54684 21476 54740 21486
rect 54012 19394 54068 19404
rect 54124 21140 54180 21150
rect 54124 17892 54180 21084
rect 54124 17826 54180 17836
rect 54460 18788 54516 18798
rect 54460 17108 54516 18732
rect 54460 15988 54516 17052
rect 54460 15922 54516 15932
rect 53900 13570 53956 13580
rect 54684 9828 54740 21420
rect 54796 11172 54852 26236
rect 54908 19572 54964 26908
rect 55356 25844 55412 31164
rect 55468 26908 55524 36428
rect 55580 30100 55636 44940
rect 55804 38612 55860 46508
rect 57708 46564 57764 46574
rect 57708 46116 57764 46508
rect 56700 43428 56756 43438
rect 55804 38546 55860 38556
rect 56140 41860 56196 41870
rect 55580 29764 55636 30044
rect 55580 29698 55636 29708
rect 56028 35364 56084 35374
rect 56028 28980 56084 35308
rect 56140 34132 56196 41804
rect 56700 38668 56756 43372
rect 57708 39620 57764 46060
rect 57708 39554 57764 39564
rect 56140 34066 56196 34076
rect 56588 38612 56756 38668
rect 56588 34132 56644 38612
rect 56476 31780 56532 31790
rect 56476 30100 56532 31724
rect 56588 30660 56644 34076
rect 56588 30594 56644 30604
rect 56588 30100 56644 30110
rect 56476 30044 56588 30100
rect 55468 26852 55860 26908
rect 55356 25778 55412 25788
rect 55244 23380 55300 23390
rect 54908 17444 54964 19516
rect 54908 12180 54964 17388
rect 54908 11620 54964 12124
rect 55020 22372 55076 22382
rect 55020 11844 55076 22316
rect 55244 21700 55300 23324
rect 55244 21634 55300 21644
rect 55468 22596 55524 22606
rect 55468 21252 55524 22540
rect 55804 22484 55860 26852
rect 56028 23268 56084 28924
rect 56252 28308 56308 28318
rect 56252 26068 56308 28252
rect 56252 26002 56308 26012
rect 56028 23202 56084 23212
rect 56476 25508 56532 25518
rect 55804 22418 55860 22428
rect 55468 21186 55524 21196
rect 56364 21700 56420 21710
rect 55132 19348 55188 19358
rect 55132 19012 55188 19292
rect 55132 12404 55188 18956
rect 55468 19012 55524 19022
rect 55468 15652 55524 18956
rect 55468 15586 55524 15596
rect 55132 12338 55188 12348
rect 56028 14308 56084 14318
rect 55020 11778 55076 11788
rect 54908 11554 54964 11564
rect 54796 11106 54852 11116
rect 54684 9762 54740 9772
rect 53788 7746 53844 7756
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 56028 6132 56084 14252
rect 56364 13188 56420 21644
rect 56476 19012 56532 25452
rect 56476 18946 56532 18956
rect 56364 13122 56420 13132
rect 56476 18676 56532 18686
rect 56028 6066 56084 6076
rect 56476 10500 56532 18620
rect 56588 15540 56644 30044
rect 57484 25060 57540 25070
rect 56588 15474 56644 15484
rect 56924 23492 56980 23502
rect 56924 22932 56980 23436
rect 57484 23492 57540 25004
rect 57484 23426 57540 23436
rect 56924 22260 56980 22876
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 56476 2996 56532 10444
rect 56924 10052 56980 22204
rect 57372 22036 57428 22046
rect 57260 19124 57316 19134
rect 57260 17444 57316 19068
rect 57260 17378 57316 17388
rect 57372 16324 57428 21980
rect 57372 16258 57428 16268
rect 57708 20804 57764 20814
rect 57708 15316 57764 20748
rect 57708 15250 57764 15260
rect 56924 8820 56980 9996
rect 56924 8754 56980 8764
rect 56476 2930 56532 2940
rect 49644 2884 49700 2894
rect 49196 2772 49252 2782
rect 49644 2772 49700 2828
rect 49252 2716 49700 2772
rect 49196 2706 49252 2716
rect 39900 1586 39956 1596
rect 26572 1474 26628 1484
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1444__I dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 52080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1446__I
timestamp 1669390400
transform 1 0 54880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1448__I
timestamp 1669390400
transform 1 0 57904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__I
timestamp 1669390400
transform 1 0 57344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1450__I
timestamp 1669390400
transform 1 0 48496 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1452__I
timestamp 1669390400
transform 1 0 57120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__I
timestamp 1669390400
transform 1 0 57792 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A1
timestamp 1669390400
transform -1 0 53536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1456__A2
timestamp 1669390400
transform -1 0 54320 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A1
timestamp 1669390400
transform 1 0 55328 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A2
timestamp 1669390400
transform 1 0 55776 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__A4
timestamp 1669390400
transform 1 0 56224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1458__I
timestamp 1669390400
transform -1 0 42560 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1459__I
timestamp 1669390400
transform -1 0 38752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1460__I
timestamp 1669390400
transform -1 0 22512 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__I
timestamp 1669390400
transform -1 0 13664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__I
timestamp 1669390400
transform 1 0 21504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1464__I
timestamp 1669390400
transform 1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1465__I
timestamp 1669390400
transform 1 0 25648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1467__I
timestamp 1669390400
transform -1 0 23072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__I
timestamp 1669390400
transform 1 0 24864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1471__I
timestamp 1669390400
transform 1 0 19936 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__A2
timestamp 1669390400
transform 1 0 29456 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__A1
timestamp 1669390400
transform 1 0 22400 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1474__A2
timestamp 1669390400
transform 1 0 23744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1475__I
timestamp 1669390400
transform -1 0 4256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1476__I
timestamp 1669390400
transform 1 0 29904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__I
timestamp 1669390400
transform 1 0 29008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1478__A1
timestamp 1669390400
transform 1 0 19264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1479__I
timestamp 1669390400
transform -1 0 22288 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1480__I
timestamp 1669390400
transform 1 0 3472 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A1
timestamp 1669390400
transform -1 0 5152 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1484__A2
timestamp 1669390400
transform 1 0 4032 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1486__I
timestamp 1669390400
transform 1 0 5264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1487__I
timestamp 1669390400
transform 1 0 29232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A1
timestamp 1669390400
transform 1 0 27888 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__B
timestamp 1669390400
transform 1 0 22960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A1
timestamp 1669390400
transform 1 0 20384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A2
timestamp 1669390400
transform 1 0 15344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1490__A3
timestamp 1669390400
transform 1 0 19488 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1492__I
timestamp 1669390400
transform -1 0 3808 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1494__I
timestamp 1669390400
transform 1 0 30800 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1495__I
timestamp 1669390400
transform 1 0 24080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1496__I
timestamp 1669390400
transform 1 0 4928 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1498__I
timestamp 1669390400
transform 1 0 30352 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A1
timestamp 1669390400
transform 1 0 11312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__A2
timestamp 1669390400
transform -1 0 2016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1500__B
timestamp 1669390400
transform -1 0 8288 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1501__A2
timestamp 1669390400
transform -1 0 21616 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1503__I
timestamp 1669390400
transform 1 0 20272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__I
timestamp 1669390400
transform 1 0 22512 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__B
timestamp 1669390400
transform 1 0 24528 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1506__C
timestamp 1669390400
transform 1 0 22064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1507__A2
timestamp 1669390400
transform -1 0 21840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A1
timestamp 1669390400
transform 1 0 25536 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1508__A2
timestamp 1669390400
transform -1 0 25984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1510__A1
timestamp 1669390400
transform -1 0 21392 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__I
timestamp 1669390400
transform 1 0 49616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1515__I
timestamp 1669390400
transform 1 0 40096 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1516__I
timestamp 1669390400
transform 1 0 34384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1517__I
timestamp 1669390400
transform 1 0 31920 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1520__I
timestamp 1669390400
transform 1 0 28112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A2
timestamp 1669390400
transform 1 0 32928 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1522__A1
timestamp 1669390400
transform 1 0 31696 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1523__A1
timestamp 1669390400
transform -1 0 29568 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A1
timestamp 1669390400
transform -1 0 32480 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1524__A2
timestamp 1669390400
transform -1 0 31360 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__I
timestamp 1669390400
transform 1 0 17696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__I
timestamp 1669390400
transform 1 0 20832 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1530__A1
timestamp 1669390400
transform -1 0 28336 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1531__A2
timestamp 1669390400
transform 1 0 27664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1533__A1
timestamp 1669390400
transform 1 0 26992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__A2
timestamp 1669390400
transform 1 0 30464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__I
timestamp 1669390400
transform -1 0 16912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1541__I
timestamp 1669390400
transform -1 0 8848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__I
timestamp 1669390400
transform -1 0 6944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1545__I
timestamp 1669390400
transform 1 0 3920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1546__I
timestamp 1669390400
transform -1 0 14336 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1548__I
timestamp 1669390400
transform 1 0 4480 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1549__A1
timestamp 1669390400
transform 1 0 4480 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A1
timestamp 1669390400
transform 1 0 6272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__A2
timestamp 1669390400
transform -1 0 8288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1552__I
timestamp 1669390400
transform 1 0 27216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A1
timestamp 1669390400
transform -1 0 19376 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__A2
timestamp 1669390400
transform -1 0 16240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A1
timestamp 1669390400
transform -1 0 4592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__A3
timestamp 1669390400
transform 1 0 4816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__B1
timestamp 1669390400
transform -1 0 2912 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1556__B2
timestamp 1669390400
transform -1 0 2240 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A1
timestamp 1669390400
transform -1 0 16912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1557__A2
timestamp 1669390400
transform -1 0 18928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A1
timestamp 1669390400
transform -1 0 30576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1559__A2
timestamp 1669390400
transform -1 0 29904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1560__I
timestamp 1669390400
transform -1 0 7952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A1
timestamp 1669390400
transform -1 0 15344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1561__A2
timestamp 1669390400
transform 1 0 13776 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A1
timestamp 1669390400
transform 1 0 15904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1562__A2
timestamp 1669390400
transform 1 0 12880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1563__I
timestamp 1669390400
transform -1 0 2688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1565__I
timestamp 1669390400
transform -1 0 2016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__A1
timestamp 1669390400
transform -1 0 2912 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1566__B
timestamp 1669390400
transform 1 0 3584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1568__I
timestamp 1669390400
transform 1 0 26096 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1570__I
timestamp 1669390400
transform 1 0 14560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A1
timestamp 1669390400
transform -1 0 3472 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1571__A2
timestamp 1669390400
transform -1 0 4704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1573__I
timestamp 1669390400
transform 1 0 4592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A1
timestamp 1669390400
transform -1 0 11200 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1574__A2
timestamp 1669390400
transform -1 0 10192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A1
timestamp 1669390400
transform 1 0 5824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__A2
timestamp 1669390400
transform -1 0 4144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1576__C
timestamp 1669390400
transform -1 0 4704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1577__I
timestamp 1669390400
transform 1 0 30800 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1579__I
timestamp 1669390400
transform 1 0 28560 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A1
timestamp 1669390400
transform 1 0 7840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1580__A2
timestamp 1669390400
transform -1 0 5152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__I
timestamp 1669390400
transform -1 0 3808 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A1
timestamp 1669390400
transform 1 0 10864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__A2
timestamp 1669390400
transform -1 0 8176 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1582__B
timestamp 1669390400
transform -1 0 10192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1583__A2
timestamp 1669390400
transform -1 0 11536 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1586__I
timestamp 1669390400
transform -1 0 8848 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1587__I
timestamp 1669390400
transform -1 0 2240 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1588__I
timestamp 1669390400
transform -1 0 4704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1589__I
timestamp 1669390400
transform -1 0 27328 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__I
timestamp 1669390400
transform -1 0 5600 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1593__A1
timestamp 1669390400
transform 1 0 2912 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1593__A2
timestamp 1669390400
transform -1 0 3584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__I
timestamp 1669390400
transform -1 0 2016 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__A1
timestamp 1669390400
transform 1 0 21280 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1597__B
timestamp 1669390400
transform 1 0 22400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__A1
timestamp 1669390400
transform -1 0 3808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__A2
timestamp 1669390400
transform -1 0 2240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__B1
timestamp 1669390400
transform -1 0 8736 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__B2
timestamp 1669390400
transform -1 0 4256 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1598__C
timestamp 1669390400
transform -1 0 2016 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A1
timestamp 1669390400
transform -1 0 2464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1599__A2
timestamp 1669390400
transform 1 0 3136 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A1
timestamp 1669390400
transform 1 0 8960 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1601__A2
timestamp 1669390400
transform 1 0 4928 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1602__A1
timestamp 1669390400
transform -1 0 6496 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__I
timestamp 1669390400
transform 1 0 7168 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A1
timestamp 1669390400
transform -1 0 5152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__A2
timestamp 1669390400
transform -1 0 5936 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1605__B
timestamp 1669390400
transform 1 0 10304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A2
timestamp 1669390400
transform 1 0 8960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A3
timestamp 1669390400
transform -1 0 15456 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1607__I
timestamp 1669390400
transform -1 0 3584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__I
timestamp 1669390400
transform -1 0 5600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A1
timestamp 1669390400
transform -1 0 2464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A3
timestamp 1669390400
transform -1 0 4368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A1
timestamp 1669390400
transform -1 0 2912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1611__A2
timestamp 1669390400
transform -1 0 2016 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1614__I
timestamp 1669390400
transform -1 0 3024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1616__I
timestamp 1669390400
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A1
timestamp 1669390400
transform -1 0 3808 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1617__A2
timestamp 1669390400
transform -1 0 10640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__I0
timestamp 1669390400
transform -1 0 3920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__I1
timestamp 1669390400
transform -1 0 2912 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1618__S
timestamp 1669390400
transform -1 0 3360 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__B1
timestamp 1669390400
transform -1 0 4256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1619__C2
timestamp 1669390400
transform 1 0 2464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1620__A1
timestamp 1669390400
transform 1 0 25984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1621__A1
timestamp 1669390400
transform 1 0 26992 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1622__I
timestamp 1669390400
transform 1 0 27664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__A1
timestamp 1669390400
transform -1 0 19824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1623__B
timestamp 1669390400
transform 1 0 20384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A1
timestamp 1669390400
transform 1 0 8512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A2
timestamp 1669390400
transform -1 0 9744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A3
timestamp 1669390400
transform -1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1624__A4
timestamp 1669390400
transform -1 0 1904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1625__A2
timestamp 1669390400
transform -1 0 6048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1626__A1
timestamp 1669390400
transform -1 0 7392 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A1
timestamp 1669390400
transform 1 0 27664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1627__A2
timestamp 1669390400
transform -1 0 27440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1628__A1
timestamp 1669390400
transform 1 0 23632 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A1
timestamp 1669390400
transform 1 0 28336 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__A2
timestamp 1669390400
transform 1 0 30128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1630__B
timestamp 1669390400
transform -1 0 25760 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A1
timestamp 1669390400
transform 1 0 22288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A2
timestamp 1669390400
transform -1 0 21840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__B
timestamp 1669390400
transform 1 0 20720 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A2
timestamp 1669390400
transform 1 0 29904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A1
timestamp 1669390400
transform 1 0 16464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1634__A2
timestamp 1669390400
transform -1 0 20048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__A2
timestamp 1669390400
transform 1 0 24752 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__B1
timestamp 1669390400
transform -1 0 25312 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__B2
timestamp 1669390400
transform 1 0 22960 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A1
timestamp 1669390400
transform -1 0 4480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1636__A2
timestamp 1669390400
transform -1 0 4928 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__A1
timestamp 1669390400
transform -1 0 4704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1638__A2
timestamp 1669390400
transform -1 0 4144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1639__I
timestamp 1669390400
transform 1 0 11760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A1
timestamp 1669390400
transform -1 0 4256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1640__A2
timestamp 1669390400
transform -1 0 4704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1642__A1
timestamp 1669390400
transform -1 0 7392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1643__I
timestamp 1669390400
transform 1 0 8960 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1644__I
timestamp 1669390400
transform 1 0 28112 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1645__I
timestamp 1669390400
transform 1 0 29904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A1
timestamp 1669390400
transform -1 0 2352 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1646__A2
timestamp 1669390400
transform -1 0 4704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1647__I
timestamp 1669390400
transform -1 0 9856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1649__I
timestamp 1669390400
transform 1 0 12992 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1650__I
timestamp 1669390400
transform -1 0 3360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1651__I
timestamp 1669390400
transform 1 0 12432 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1652__A1
timestamp 1669390400
transform -1 0 5824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A1
timestamp 1669390400
transform -1 0 3472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__A2
timestamp 1669390400
transform -1 0 1904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__B
timestamp 1669390400
transform -1 0 2800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1654__A3
timestamp 1669390400
transform 1 0 4480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A1
timestamp 1669390400
transform -1 0 2016 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1655__A2
timestamp 1669390400
transform 1 0 2240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A1
timestamp 1669390400
transform -1 0 4368 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__A2
timestamp 1669390400
transform -1 0 3808 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A1
timestamp 1669390400
transform -1 0 11088 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__A2
timestamp 1669390400
transform 1 0 9520 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__B1
timestamp 1669390400
transform -1 0 8400 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1658__B2
timestamp 1669390400
transform 1 0 7728 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1661__I
timestamp 1669390400
transform -1 0 22960 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__I
timestamp 1669390400
transform 1 0 18928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__I
timestamp 1669390400
transform 1 0 7616 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__I
timestamp 1669390400
transform 1 0 7168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__I
timestamp 1669390400
transform -1 0 5152 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__A1
timestamp 1669390400
transform 1 0 8176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__B
timestamp 1669390400
transform -1 0 10080 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__I
timestamp 1669390400
transform 1 0 5712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A1
timestamp 1669390400
transform -1 0 3808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__A2
timestamp 1669390400
transform -1 0 4256 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A1
timestamp 1669390400
transform 1 0 4032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__A2
timestamp 1669390400
transform 1 0 5264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__I
timestamp 1669390400
transform 1 0 5264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A1
timestamp 1669390400
transform -1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__A2
timestamp 1669390400
transform -1 0 8736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__I
timestamp 1669390400
transform 1 0 23856 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A1
timestamp 1669390400
transform -1 0 22736 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__A2
timestamp 1669390400
transform 1 0 20832 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__B
timestamp 1669390400
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__A2
timestamp 1669390400
transform 1 0 23408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__B
timestamp 1669390400
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__I
timestamp 1669390400
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__A2
timestamp 1669390400
transform -1 0 22848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__B
timestamp 1669390400
transform 1 0 29904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__I
timestamp 1669390400
transform -1 0 19376 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__I
timestamp 1669390400
transform 1 0 3696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A1
timestamp 1669390400
transform 1 0 5712 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A2
timestamp 1669390400
transform 1 0 7616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__A3
timestamp 1669390400
transform 1 0 3136 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A1
timestamp 1669390400
transform -1 0 3248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__A2
timestamp 1669390400
transform -1 0 3696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__A2
timestamp 1669390400
transform 1 0 3920 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__B1
timestamp 1669390400
transform -1 0 5152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__A2
timestamp 1669390400
transform -1 0 6160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__B
timestamp 1669390400
transform -1 0 6608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__I
timestamp 1669390400
transform 1 0 9072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A1
timestamp 1669390400
transform -1 0 3360 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__A2
timestamp 1669390400
transform -1 0 2128 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A1
timestamp 1669390400
transform -1 0 3808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__A2
timestamp 1669390400
transform -1 0 1904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__B
timestamp 1669390400
transform -1 0 4704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__A2
timestamp 1669390400
transform 1 0 8064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__B
timestamp 1669390400
transform -1 0 6944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__A1
timestamp 1669390400
transform -1 0 6384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__B
timestamp 1669390400
transform -1 0 7392 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A1
timestamp 1669390400
transform 1 0 25536 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__A2
timestamp 1669390400
transform -1 0 25872 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A1
timestamp 1669390400
transform -1 0 10304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__A3
timestamp 1669390400
transform 1 0 9632 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__B1
timestamp 1669390400
transform -1 0 2240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__B2
timestamp 1669390400
transform -1 0 2016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1701__A3
timestamp 1669390400
transform 1 0 5376 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1702__A1
timestamp 1669390400
transform -1 0 7392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1704__I
timestamp 1669390400
transform 1 0 19600 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1706__I
timestamp 1669390400
transform -1 0 19264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A1
timestamp 1669390400
transform -1 0 15904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__A2
timestamp 1669390400
transform 1 0 17248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__B
timestamp 1669390400
transform 1 0 16800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__A2
timestamp 1669390400
transform -1 0 2912 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__B1
timestamp 1669390400
transform -1 0 2240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1708__B2
timestamp 1669390400
transform -1 0 3696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A1
timestamp 1669390400
transform 1 0 31248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__A2
timestamp 1669390400
transform 1 0 28560 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__A2
timestamp 1669390400
transform -1 0 2352 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__A1
timestamp 1669390400
transform -1 0 1904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__C
timestamp 1669390400
transform 1 0 3360 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__I
timestamp 1669390400
transform 1 0 18816 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A1
timestamp 1669390400
transform 1 0 10752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1713__A2
timestamp 1669390400
transform -1 0 2016 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A1
timestamp 1669390400
transform -1 0 4256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__A2
timestamp 1669390400
transform 1 0 6496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1716__I
timestamp 1669390400
transform 1 0 21840 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__A1
timestamp 1669390400
transform 1 0 28224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1717__A2
timestamp 1669390400
transform 1 0 24640 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1718__I
timestamp 1669390400
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A1
timestamp 1669390400
transform 1 0 26432 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__A2
timestamp 1669390400
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1719__B
timestamp 1669390400
transform 1 0 30352 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__A1
timestamp 1669390400
transform -1 0 24304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__A2
timestamp 1669390400
transform 1 0 21840 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__A2
timestamp 1669390400
transform -1 0 10080 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__A1
timestamp 1669390400
transform 1 0 11648 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A1
timestamp 1669390400
transform -1 0 7728 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__A2
timestamp 1669390400
transform 1 0 9520 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__I
timestamp 1669390400
transform 1 0 14560 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__A2
timestamp 1669390400
transform 1 0 10192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__A1
timestamp 1669390400
transform 1 0 12880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__A2
timestamp 1669390400
transform -1 0 5040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__A1
timestamp 1669390400
transform -1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__A2
timestamp 1669390400
transform 1 0 12208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A1
timestamp 1669390400
transform -1 0 2016 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__A2
timestamp 1669390400
transform -1 0 5152 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__I
timestamp 1669390400
transform -1 0 14112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__I0
timestamp 1669390400
transform 1 0 15680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__S0
timestamp 1669390400
transform 1 0 4928 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__I
timestamp 1669390400
transform 1 0 31248 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__I
timestamp 1669390400
transform -1 0 3360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A1
timestamp 1669390400
transform -1 0 9072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__A2
timestamp 1669390400
transform -1 0 10640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__B
timestamp 1669390400
transform -1 0 5488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__C
timestamp 1669390400
transform 1 0 8400 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__A2
timestamp 1669390400
transform 1 0 13104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A1
timestamp 1669390400
transform -1 0 8288 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__A3
timestamp 1669390400
transform -1 0 7840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__I
timestamp 1669390400
transform -1 0 10976 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__I
timestamp 1669390400
transform -1 0 18928 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__A1
timestamp 1669390400
transform 1 0 10752 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__B
timestamp 1669390400
transform -1 0 11424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__I
timestamp 1669390400
transform -1 0 6832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__I
timestamp 1669390400
transform -1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__A1
timestamp 1669390400
transform -1 0 8176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A1
timestamp 1669390400
transform 1 0 6720 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__A3
timestamp 1669390400
transform -1 0 8848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__A1
timestamp 1669390400
transform -1 0 7056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__A2
timestamp 1669390400
transform 1 0 6048 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A1
timestamp 1669390400
transform -1 0 3472 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__A2
timestamp 1669390400
transform -1 0 4592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__B1
timestamp 1669390400
transform -1 0 4256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__B2
timestamp 1669390400
transform -1 0 2576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__A1
timestamp 1669390400
transform 1 0 11200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__A2
timestamp 1669390400
transform -1 0 11648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__A1
timestamp 1669390400
transform 1 0 25536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__A3
timestamp 1669390400
transform 1 0 26544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__A1
timestamp 1669390400
transform 1 0 31360 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__A2
timestamp 1669390400
transform 1 0 27328 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__A2
timestamp 1669390400
transform -1 0 14896 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__B1
timestamp 1669390400
transform 1 0 14112 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__B2
timestamp 1669390400
transform 1 0 13664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__C
timestamp 1669390400
transform 1 0 14560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__A1
timestamp 1669390400
transform 1 0 4480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A1
timestamp 1669390400
transform -1 0 2464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__A2
timestamp 1669390400
transform -1 0 2912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A1
timestamp 1669390400
transform -1 0 10752 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A2
timestamp 1669390400
transform -1 0 12432 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__A3
timestamp 1669390400
transform -1 0 10528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A1
timestamp 1669390400
transform -1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A2
timestamp 1669390400
transform -1 0 10976 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__A3
timestamp 1669390400
transform 1 0 11648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__A1
timestamp 1669390400
transform 1 0 8960 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__A2
timestamp 1669390400
transform -1 0 5152 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A1
timestamp 1669390400
transform -1 0 2912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__A2
timestamp 1669390400
transform 1 0 3136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__B
timestamp 1669390400
transform 1 0 4032 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__I
timestamp 1669390400
transform 1 0 4032 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A1
timestamp 1669390400
transform -1 0 9856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__A2
timestamp 1669390400
transform -1 0 2464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__A1
timestamp 1669390400
transform 1 0 2912 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A1
timestamp 1669390400
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A2
timestamp 1669390400
transform -1 0 15232 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__A3
timestamp 1669390400
transform -1 0 8176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__I
timestamp 1669390400
transform 1 0 17920 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__I
timestamp 1669390400
transform 1 0 15680 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A1
timestamp 1669390400
transform 1 0 8960 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A2
timestamp 1669390400
transform -1 0 16800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__A3
timestamp 1669390400
transform -1 0 10192 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__A1
timestamp 1669390400
transform -1 0 2464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__A2
timestamp 1669390400
transform -1 0 3248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__I
timestamp 1669390400
transform 1 0 23968 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A1
timestamp 1669390400
transform -1 0 22960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A2
timestamp 1669390400
transform 1 0 24528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__A3
timestamp 1669390400
transform -1 0 17248 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__A1
timestamp 1669390400
transform -1 0 2912 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__B1
timestamp 1669390400
transform -1 0 2352 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__B2
timestamp 1669390400
transform -1 0 2240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__A1
timestamp 1669390400
transform -1 0 2464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__B1
timestamp 1669390400
transform 1 0 11984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__A1
timestamp 1669390400
transform 1 0 24080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__I
timestamp 1669390400
transform 1 0 21504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A1
timestamp 1669390400
transform 1 0 14112 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1785__A2
timestamp 1669390400
transform -1 0 15232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__I
timestamp 1669390400
transform 1 0 24640 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A1
timestamp 1669390400
transform 1 0 11760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__A2
timestamp 1669390400
transform 1 0 11312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__B
timestamp 1669390400
transform 1 0 20832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__C
timestamp 1669390400
transform -1 0 21952 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A1
timestamp 1669390400
transform -1 0 17136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__A2
timestamp 1669390400
transform 1 0 16128 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__B
timestamp 1669390400
transform 1 0 12768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__A1
timestamp 1669390400
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__B
timestamp 1669390400
transform 1 0 16912 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A1
timestamp 1669390400
transform 1 0 30128 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__A2
timestamp 1669390400
transform 1 0 31136 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A1
timestamp 1669390400
transform -1 0 2464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__A3
timestamp 1669390400
transform 1 0 5824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__B
timestamp 1669390400
transform -1 0 13440 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__C
timestamp 1669390400
transform 1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__A2
timestamp 1669390400
transform -1 0 16352 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__B1
timestamp 1669390400
transform -1 0 16128 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__C
timestamp 1669390400
transform 1 0 10416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__A1
timestamp 1669390400
transform -1 0 11088 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__A2
timestamp 1669390400
transform -1 0 12208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__B1
timestamp 1669390400
transform -1 0 12656 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__B2
timestamp 1669390400
transform -1 0 12208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A1
timestamp 1669390400
transform 1 0 18816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__A2
timestamp 1669390400
transform -1 0 21056 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__B
timestamp 1669390400
transform 1 0 21056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A1
timestamp 1669390400
transform 1 0 31248 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__A2
timestamp 1669390400
transform -1 0 15680 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__B
timestamp 1669390400
transform -1 0 21392 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1800__A2
timestamp 1669390400
transform 1 0 17920 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A1
timestamp 1669390400
transform 1 0 21392 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A2
timestamp 1669390400
transform 1 0 22400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1801__A3
timestamp 1669390400
transform 1 0 23632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__A1
timestamp 1669390400
transform 1 0 30800 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1802__B2
timestamp 1669390400
transform 1 0 25536 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A2
timestamp 1669390400
transform -1 0 8512 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__A3
timestamp 1669390400
transform -1 0 16016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1805__I
timestamp 1669390400
transform -1 0 15904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1806__A1
timestamp 1669390400
transform 1 0 24752 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1807__I
timestamp 1669390400
transform -1 0 17808 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__A1
timestamp 1669390400
transform -1 0 10304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__A2
timestamp 1669390400
transform 1 0 12656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1808__C
timestamp 1669390400
transform 1 0 6496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A1
timestamp 1669390400
transform 1 0 16016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A3
timestamp 1669390400
transform -1 0 16352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1809__A4
timestamp 1669390400
transform 1 0 12432 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__A1
timestamp 1669390400
transform -1 0 4144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1810__B2
timestamp 1669390400
transform 1 0 5600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__A1
timestamp 1669390400
transform -1 0 4256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1811__A4
timestamp 1669390400
transform -1 0 3696 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A1
timestamp 1669390400
transform 1 0 11984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1813__A2
timestamp 1669390400
transform -1 0 4032 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A1
timestamp 1669390400
transform 1 0 8064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1814__A2
timestamp 1669390400
transform 1 0 12768 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A1
timestamp 1669390400
transform -1 0 1904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__A2
timestamp 1669390400
transform -1 0 5152 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1815__B
timestamp 1669390400
transform -1 0 2800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__A1
timestamp 1669390400
transform -1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1816__A3
timestamp 1669390400
transform -1 0 6384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A1
timestamp 1669390400
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1817__A2
timestamp 1669390400
transform 1 0 14672 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__A1
timestamp 1669390400
transform -1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__B
timestamp 1669390400
transform 1 0 15008 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1818__C
timestamp 1669390400
transform -1 0 16128 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A1
timestamp 1669390400
transform 1 0 4032 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1819__A2
timestamp 1669390400
transform -1 0 6608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1821__B
timestamp 1669390400
transform -1 0 15680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A1
timestamp 1669390400
transform -1 0 13888 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__A2
timestamp 1669390400
transform 1 0 8064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1822__B
timestamp 1669390400
transform -1 0 8736 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1824__A2
timestamp 1669390400
transform -1 0 14560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A1
timestamp 1669390400
transform 1 0 6272 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1825__A4
timestamp 1669390400
transform -1 0 7392 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__A1
timestamp 1669390400
transform -1 0 3808 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1826__B
timestamp 1669390400
transform 1 0 5824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1831__I
timestamp 1669390400
transform 1 0 3584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A1
timestamp 1669390400
transform 1 0 6160 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1832__A4
timestamp 1669390400
transform 1 0 6272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A1
timestamp 1669390400
transform 1 0 4928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1833__A3
timestamp 1669390400
transform 1 0 5376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__A2
timestamp 1669390400
transform -1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1834__B
timestamp 1669390400
transform 1 0 4032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1835__B
timestamp 1669390400
transform 1 0 4928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A1
timestamp 1669390400
transform -1 0 3920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__A2
timestamp 1669390400
transform -1 0 7840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1837__B
timestamp 1669390400
transform -1 0 7840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A1
timestamp 1669390400
transform -1 0 7392 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1838__A2
timestamp 1669390400
transform -1 0 8736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__B
timestamp 1669390400
transform -1 0 14784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1839__C
timestamp 1669390400
transform -1 0 17808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__A2
timestamp 1669390400
transform -1 0 15456 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1840__B
timestamp 1669390400
transform -1 0 15456 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A1
timestamp 1669390400
transform 1 0 16912 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1841__A2
timestamp 1669390400
transform -1 0 18480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A1
timestamp 1669390400
transform 1 0 21504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__A2
timestamp 1669390400
transform -1 0 15904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__B1
timestamp 1669390400
transform -1 0 22176 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1843__C
timestamp 1669390400
transform 1 0 22736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__A1
timestamp 1669390400
transform 1 0 10080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1844__C
timestamp 1669390400
transform -1 0 11200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__A2
timestamp 1669390400
transform 1 0 6496 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1845__A3
timestamp 1669390400
transform 1 0 6048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1846__A1
timestamp 1669390400
transform -1 0 5152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__A2
timestamp 1669390400
transform -1 0 5824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1847__B
timestamp 1669390400
transform -1 0 3808 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A1
timestamp 1669390400
transform -1 0 3920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A2
timestamp 1669390400
transform 1 0 4592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1848__A4
timestamp 1669390400
transform -1 0 7840 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__A1
timestamp 1669390400
transform 1 0 21504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1849__A2
timestamp 1669390400
transform 1 0 20272 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1850__A1
timestamp 1669390400
transform 1 0 16016 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1851__A1
timestamp 1669390400
transform 1 0 21616 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A1
timestamp 1669390400
transform -1 0 19152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__A2
timestamp 1669390400
transform -1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1852__B
timestamp 1669390400
transform 1 0 18368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A1
timestamp 1669390400
transform -1 0 18368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1853__A2
timestamp 1669390400
transform -1 0 17920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1854__A2
timestamp 1669390400
transform -1 0 19600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A1
timestamp 1669390400
transform -1 0 17136 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__A2
timestamp 1669390400
transform -1 0 15792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1855__B1
timestamp 1669390400
transform -1 0 18816 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A1
timestamp 1669390400
transform -1 0 16800 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1856__A2
timestamp 1669390400
transform 1 0 18144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1857__A1
timestamp 1669390400
transform -1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A1
timestamp 1669390400
transform -1 0 15456 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1858__A2
timestamp 1669390400
transform -1 0 15680 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__A2
timestamp 1669390400
transform -1 0 11760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__B1
timestamp 1669390400
transform -1 0 13104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__B2
timestamp 1669390400
transform 1 0 12432 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1859__C
timestamp 1669390400
transform -1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A1
timestamp 1669390400
transform -1 0 10640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1860__A2
timestamp 1669390400
transform 1 0 9072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A1
timestamp 1669390400
transform 1 0 9968 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1861__A2
timestamp 1669390400
transform -1 0 9968 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1862__A1
timestamp 1669390400
transform -1 0 12096 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1863__A3
timestamp 1669390400
transform 1 0 14672 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A1
timestamp 1669390400
transform -1 0 3360 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A2
timestamp 1669390400
transform 1 0 3584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1866__A3
timestamp 1669390400
transform 1 0 5936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1867__B
timestamp 1669390400
transform -1 0 9296 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A1
timestamp 1669390400
transform -1 0 17136 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__A2
timestamp 1669390400
transform 1 0 13552 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__B1
timestamp 1669390400
transform -1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1868__B2
timestamp 1669390400
transform 1 0 19488 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A1
timestamp 1669390400
transform 1 0 11872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1869__A2
timestamp 1669390400
transform 1 0 12880 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1870__I
timestamp 1669390400
transform 1 0 8064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A1
timestamp 1669390400
transform 1 0 20720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__A2
timestamp 1669390400
transform 1 0 18592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__B1
timestamp 1669390400
transform -1 0 17360 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1872__C
timestamp 1669390400
transform 1 0 17920 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1873__A1
timestamp 1669390400
transform 1 0 15792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1874__I
timestamp 1669390400
transform 1 0 4816 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1875__I
timestamp 1669390400
transform 1 0 20048 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A1
timestamp 1669390400
transform 1 0 19040 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__A2
timestamp 1669390400
transform 1 0 22288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1876__C
timestamp 1669390400
transform -1 0 26096 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1877__A1
timestamp 1669390400
transform 1 0 19488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1878__A2
timestamp 1669390400
transform 1 0 16464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1879__A2
timestamp 1669390400
transform -1 0 12096 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1882__I
timestamp 1669390400
transform -1 0 2240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__A1
timestamp 1669390400
transform -1 0 12544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1883__A4
timestamp 1669390400
transform -1 0 12992 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1885__I
timestamp 1669390400
transform 1 0 13104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__A2
timestamp 1669390400
transform 1 0 6160 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__A3
timestamp 1669390400
transform 1 0 6608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1886__A4
timestamp 1669390400
transform 1 0 7056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A1
timestamp 1669390400
transform -1 0 5152 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__A2
timestamp 1669390400
transform -1 0 2912 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1887__B
timestamp 1669390400
transform -1 0 5824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A1
timestamp 1669390400
transform 1 0 7840 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1888__A2
timestamp 1669390400
transform 1 0 9408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1890__B
timestamp 1669390400
transform -1 0 13888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__A1
timestamp 1669390400
transform 1 0 3584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__B1
timestamp 1669390400
transform 1 0 11648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__B2
timestamp 1669390400
transform -1 0 12880 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1891__C
timestamp 1669390400
transform -1 0 2688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1892__B
timestamp 1669390400
transform 1 0 2912 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__A1
timestamp 1669390400
transform 1 0 7504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1893__A2
timestamp 1669390400
transform 1 0 9072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A2
timestamp 1669390400
transform 1 0 9632 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A3
timestamp 1669390400
transform 1 0 9184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1895__A4
timestamp 1669390400
transform -1 0 8624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A1
timestamp 1669390400
transform 1 0 6944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1896__A2
timestamp 1669390400
transform -1 0 7168 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1897__B
timestamp 1669390400
transform 1 0 7280 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1898__A2
timestamp 1669390400
transform -1 0 12544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A1
timestamp 1669390400
transform -1 0 7392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1899__A2
timestamp 1669390400
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A1
timestamp 1669390400
transform 1 0 31248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__A2
timestamp 1669390400
transform 1 0 28112 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1900__B
timestamp 1669390400
transform 1 0 30800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A1
timestamp 1669390400
transform 1 0 2464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A2
timestamp 1669390400
transform -1 0 2912 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1901__A3
timestamp 1669390400
transform -1 0 3360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A1
timestamp 1669390400
transform 1 0 16016 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1902__A2
timestamp 1669390400
transform -1 0 17136 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1903__A2
timestamp 1669390400
transform -1 0 4704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1904__I
timestamp 1669390400
transform 1 0 15120 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A1
timestamp 1669390400
transform -1 0 15680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1905__A2
timestamp 1669390400
transform 1 0 6048 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__A1
timestamp 1669390400
transform 1 0 12208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1906__A2
timestamp 1669390400
transform -1 0 11984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__A1
timestamp 1669390400
transform 1 0 17360 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1907__C
timestamp 1669390400
transform -1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__A1
timestamp 1669390400
transform -1 0 14000 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1908__A2
timestamp 1669390400
transform -1 0 10752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A1
timestamp 1669390400
transform 1 0 16016 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A2
timestamp 1669390400
transform 1 0 15008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1909__A3
timestamp 1669390400
transform 1 0 12880 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1910__A1
timestamp 1669390400
transform 1 0 15568 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1912__A2
timestamp 1669390400
transform -1 0 7840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__A2
timestamp 1669390400
transform -1 0 2688 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1913__B
timestamp 1669390400
transform -1 0 4256 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A1
timestamp 1669390400
transform -1 0 4368 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A2
timestamp 1669390400
transform -1 0 3696 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1914__A4
timestamp 1669390400
transform 1 0 8512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__A1
timestamp 1669390400
transform -1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1915__B
timestamp 1669390400
transform -1 0 9856 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1916__A1
timestamp 1669390400
transform -1 0 2016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A1
timestamp 1669390400
transform 1 0 13216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__A2
timestamp 1669390400
transform 1 0 12768 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1917__B
timestamp 1669390400
transform -1 0 15232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A1
timestamp 1669390400
transform -1 0 11536 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A2
timestamp 1669390400
transform -1 0 13552 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1918__A3
timestamp 1669390400
transform -1 0 12992 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A1
timestamp 1669390400
transform 1 0 15008 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1919__A2
timestamp 1669390400
transform 1 0 11984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A1
timestamp 1669390400
transform 1 0 11088 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1920__A2
timestamp 1669390400
transform -1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A1
timestamp 1669390400
transform 1 0 11088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1921__A2
timestamp 1669390400
transform -1 0 11760 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A1
timestamp 1669390400
transform -1 0 18928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A2
timestamp 1669390400
transform -1 0 17808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__A3
timestamp 1669390400
transform -1 0 8960 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1923__B
timestamp 1669390400
transform 1 0 5936 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__A1
timestamp 1669390400
transform 1 0 16464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1924__B2
timestamp 1669390400
transform 1 0 12880 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1925__I
timestamp 1669390400
transform 1 0 30800 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A1
timestamp 1669390400
transform 1 0 16576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A2
timestamp 1669390400
transform 1 0 16912 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1926__A3
timestamp 1669390400
transform 1 0 16128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A1
timestamp 1669390400
transform 1 0 18592 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A2
timestamp 1669390400
transform 1 0 16464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1928__A3
timestamp 1669390400
transform 1 0 17696 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1929__A1
timestamp 1669390400
transform -1 0 19376 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1930__A1
timestamp 1669390400
transform 1 0 17920 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1931__A2
timestamp 1669390400
transform -1 0 17360 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1933__A2
timestamp 1669390400
transform -1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1942__I
timestamp 1669390400
transform 1 0 26320 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A1
timestamp 1669390400
transform -1 0 12656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1944__A2
timestamp 1669390400
transform 1 0 11536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1945__A2
timestamp 1669390400
transform 1 0 14896 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A1
timestamp 1669390400
transform -1 0 8288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A2
timestamp 1669390400
transform -1 0 3360 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__A3
timestamp 1669390400
transform -1 0 2016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1946__B
timestamp 1669390400
transform -1 0 6832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A1
timestamp 1669390400
transform -1 0 2240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1947__A2
timestamp 1669390400
transform -1 0 2688 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A1
timestamp 1669390400
transform 1 0 31136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1948__A2
timestamp 1669390400
transform 1 0 27776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1949__A1
timestamp 1669390400
transform 1 0 26432 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A1
timestamp 1669390400
transform 1 0 28224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1950__A2
timestamp 1669390400
transform 1 0 26768 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A1
timestamp 1669390400
transform 1 0 4368 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1951__A2
timestamp 1669390400
transform -1 0 5040 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__A2
timestamp 1669390400
transform -1 0 4032 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1952__B
timestamp 1669390400
transform -1 0 2352 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A1
timestamp 1669390400
transform 1 0 9632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1956__A2
timestamp 1669390400
transform 1 0 10864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1958__A1
timestamp 1669390400
transform -1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__A2
timestamp 1669390400
transform 1 0 6720 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1959__B
timestamp 1669390400
transform 1 0 4480 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A1
timestamp 1669390400
transform -1 0 16352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1960__A3
timestamp 1669390400
transform 1 0 16912 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1961__A2
timestamp 1669390400
transform -1 0 16352 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1963__A1
timestamp 1669390400
transform 1 0 24752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A1
timestamp 1669390400
transform 1 0 3584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A2
timestamp 1669390400
transform -1 0 13328 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1964__A3
timestamp 1669390400
transform -1 0 15904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__A2
timestamp 1669390400
transform 1 0 15232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1965__B
timestamp 1669390400
transform -1 0 8960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__A2
timestamp 1669390400
transform 1 0 11648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1966__B
timestamp 1669390400
transform 1 0 16464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__A1
timestamp 1669390400
transform -1 0 19936 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__A2
timestamp 1669390400
transform 1 0 22960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__B2
timestamp 1669390400
transform 1 0 22512 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1967__C
timestamp 1669390400
transform -1 0 19936 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1968__A1
timestamp 1669390400
transform -1 0 5152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A1
timestamp 1669390400
transform 1 0 16128 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1969__A2
timestamp 1669390400
transform -1 0 18368 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1970__A2
timestamp 1669390400
transform -1 0 17360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A1
timestamp 1669390400
transform -1 0 19264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A2
timestamp 1669390400
transform 1 0 18816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1971__A3
timestamp 1669390400
transform 1 0 19264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1973__A1
timestamp 1669390400
transform -1 0 16912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1974__A1
timestamp 1669390400
transform -1 0 18816 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A1
timestamp 1669390400
transform 1 0 11760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1975__A2
timestamp 1669390400
transform -1 0 13328 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A1
timestamp 1669390400
transform 1 0 11536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__A2
timestamp 1669390400
transform 1 0 13552 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1976__B
timestamp 1669390400
transform 1 0 11984 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1978__I
timestamp 1669390400
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1979__I
timestamp 1669390400
transform 1 0 12320 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__A1
timestamp 1669390400
transform -1 0 14896 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1980__A2
timestamp 1669390400
transform 1 0 12208 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__A1
timestamp 1669390400
transform -1 0 17024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1981__A2
timestamp 1669390400
transform 1 0 16016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1982__I
timestamp 1669390400
transform 1 0 23856 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A1
timestamp 1669390400
transform 1 0 11424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1983__A2
timestamp 1669390400
transform 1 0 14448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1984__A2
timestamp 1669390400
transform -1 0 4704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__A1
timestamp 1669390400
transform -1 0 3360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1985__B
timestamp 1669390400
transform 1 0 2240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1986__A1
timestamp 1669390400
transform 1 0 2464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__A1
timestamp 1669390400
transform -1 0 18480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1987__B
timestamp 1669390400
transform 1 0 16016 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1988__I
timestamp 1669390400
transform 1 0 20944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1989__A2
timestamp 1669390400
transform -1 0 19936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1992__A3
timestamp 1669390400
transform 1 0 15120 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A1
timestamp 1669390400
transform 1 0 14000 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1997__A2
timestamp 1669390400
transform 1 0 14672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1998__A3
timestamp 1669390400
transform 1 0 14896 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__A1
timestamp 1669390400
transform -1 0 19264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2000__A2
timestamp 1669390400
transform 1 0 22512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2001__A2
timestamp 1669390400
transform -1 0 20720 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A2
timestamp 1669390400
transform 1 0 26880 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A3
timestamp 1669390400
transform 1 0 30800 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2002__A4
timestamp 1669390400
transform 1 0 27328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A1
timestamp 1669390400
transform 1 0 24864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2003__A3
timestamp 1669390400
transform 1 0 25648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2005__C
timestamp 1669390400
transform 1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A1
timestamp 1669390400
transform 1 0 29456 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2006__A2
timestamp 1669390400
transform 1 0 27216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A1
timestamp 1669390400
transform 1 0 19152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2008__A2
timestamp 1669390400
transform 1 0 17584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2009__A1
timestamp 1669390400
transform -1 0 18704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A1
timestamp 1669390400
transform 1 0 16912 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2010__A2
timestamp 1669390400
transform -1 0 14448 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2011__A1
timestamp 1669390400
transform -1 0 15344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A1
timestamp 1669390400
transform -1 0 2464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2012__A3
timestamp 1669390400
transform -1 0 4704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A1
timestamp 1669390400
transform -1 0 2800 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2013__A3
timestamp 1669390400
transform -1 0 3360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A1
timestamp 1669390400
transform -1 0 3808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2014__A3
timestamp 1669390400
transform -1 0 4256 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2015__C
timestamp 1669390400
transform -1 0 4704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2017__S
timestamp 1669390400
transform 1 0 18032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A1
timestamp 1669390400
transform 1 0 14672 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2018__A2
timestamp 1669390400
transform 1 0 16240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A1
timestamp 1669390400
transform 1 0 14224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2019__A2
timestamp 1669390400
transform -1 0 15344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2020__A1
timestamp 1669390400
transform 1 0 13552 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2021__B
timestamp 1669390400
transform 1 0 21840 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A1
timestamp 1669390400
transform 1 0 19600 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__A2
timestamp 1669390400
transform -1 0 19040 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2022__B
timestamp 1669390400
transform -1 0 21728 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A1
timestamp 1669390400
transform -1 0 12656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__A2
timestamp 1669390400
transform -1 0 9856 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__B1
timestamp 1669390400
transform 1 0 9296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2024__B2
timestamp 1669390400
transform 1 0 11760 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__A1
timestamp 1669390400
transform -1 0 17136 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2025__A2
timestamp 1669390400
transform -1 0 15232 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2029__B
timestamp 1669390400
transform -1 0 12880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2035__I
timestamp 1669390400
transform -1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__A1
timestamp 1669390400
transform 1 0 18032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2036__A2
timestamp 1669390400
transform 1 0 17248 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__A2
timestamp 1669390400
transform 1 0 14112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__B
timestamp 1669390400
transform -1 0 13888 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2038__C
timestamp 1669390400
transform -1 0 12656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2039__A2
timestamp 1669390400
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__A1
timestamp 1669390400
transform 1 0 4928 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2040__B
timestamp 1669390400
transform -1 0 5936 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A1
timestamp 1669390400
transform -1 0 22736 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__A2
timestamp 1669390400
transform -1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2042__B2
timestamp 1669390400
transform -1 0 21056 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__A1
timestamp 1669390400
transform -1 0 15792 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2043__B
timestamp 1669390400
transform -1 0 17808 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2044__A3
timestamp 1669390400
transform -1 0 17808 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A1
timestamp 1669390400
transform 1 0 19152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__A2
timestamp 1669390400
transform -1 0 18704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2045__B
timestamp 1669390400
transform 1 0 19824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2046__A2
timestamp 1669390400
transform -1 0 21728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A1
timestamp 1669390400
transform 1 0 30576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2047__A2
timestamp 1669390400
transform 1 0 29456 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__A1
timestamp 1669390400
transform -1 0 17920 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2048__A2
timestamp 1669390400
transform 1 0 20832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A1
timestamp 1669390400
transform 1 0 15568 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__A2
timestamp 1669390400
transform 1 0 23968 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2049__C
timestamp 1669390400
transform 1 0 16912 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A1
timestamp 1669390400
transform 1 0 19264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2050__A2
timestamp 1669390400
transform 1 0 20832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2051__A1
timestamp 1669390400
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2051__C
timestamp 1669390400
transform -1 0 14000 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2053__B2
timestamp 1669390400
transform -1 0 18816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2055__I
timestamp 1669390400
transform -1 0 21504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A1
timestamp 1669390400
transform 1 0 22400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2056__A2
timestamp 1669390400
transform -1 0 21952 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2057__A1
timestamp 1669390400
transform 1 0 20832 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A1
timestamp 1669390400
transform 1 0 18480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2058__A3
timestamp 1669390400
transform 1 0 20832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A1
timestamp 1669390400
transform 1 0 25648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2059__A2
timestamp 1669390400
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2060__A1
timestamp 1669390400
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2061__A2
timestamp 1669390400
transform 1 0 26992 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2062__A1
timestamp 1669390400
transform 1 0 24416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A1
timestamp 1669390400
transform 1 0 23296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2063__A2
timestamp 1669390400
transform 1 0 25760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2069__I
timestamp 1669390400
transform 1 0 57904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2070__I
timestamp 1669390400
transform 1 0 20832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2071__A1
timestamp 1669390400
transform 1 0 21392 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2072__I
timestamp 1669390400
transform 1 0 19152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__A1
timestamp 1669390400
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2073__B
timestamp 1669390400
transform 1 0 29456 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__A1
timestamp 1669390400
transform -1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__A2
timestamp 1669390400
transform 1 0 18144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2074__B
timestamp 1669390400
transform -1 0 11648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2075__A2
timestamp 1669390400
transform 1 0 18032 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__A2
timestamp 1669390400
transform 1 0 8512 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2076__C
timestamp 1669390400
transform 1 0 11536 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__A1
timestamp 1669390400
transform 1 0 15120 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2077__C
timestamp 1669390400
transform -1 0 16128 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__A1
timestamp 1669390400
transform -1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__A2
timestamp 1669390400
transform 1 0 18368 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2078__A3
timestamp 1669390400
transform -1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__I0
timestamp 1669390400
transform -1 0 20272 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2079__S
timestamp 1669390400
transform -1 0 19152 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2080__A1
timestamp 1669390400
transform -1 0 18928 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2082__I
timestamp 1669390400
transform -1 0 25760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2083__A1
timestamp 1669390400
transform -1 0 22736 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2084__A1
timestamp 1669390400
transform -1 0 23296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2085__I
timestamp 1669390400
transform 1 0 28672 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2086__A1
timestamp 1669390400
transform 1 0 30800 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2087__A1
timestamp 1669390400
transform 1 0 29456 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__A1
timestamp 1669390400
transform 1 0 28112 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2088__A2
timestamp 1669390400
transform 1 0 22064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__A1
timestamp 1669390400
transform -1 0 23184 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2089__A2
timestamp 1669390400
transform 1 0 21616 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__B
timestamp 1669390400
transform 1 0 23744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2090__C
timestamp 1669390400
transform 1 0 25984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__A2
timestamp 1669390400
transform -1 0 25088 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2091__C
timestamp 1669390400
transform 1 0 22624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__A1
timestamp 1669390400
transform 1 0 16352 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__A2
timestamp 1669390400
transform 1 0 18704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__B2
timestamp 1669390400
transform -1 0 30128 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2095__C
timestamp 1669390400
transform -1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2099__A2
timestamp 1669390400
transform 1 0 23632 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2110__A2
timestamp 1669390400
transform 1 0 22288 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__A1
timestamp 1669390400
transform 1 0 25536 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__A2
timestamp 1669390400
transform 1 0 31696 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__B
timestamp 1669390400
transform 1 0 25760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2113__C
timestamp 1669390400
transform 1 0 26992 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__A1
timestamp 1669390400
transform 1 0 24416 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2114__A2
timestamp 1669390400
transform 1 0 25312 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__A1
timestamp 1669390400
transform -1 0 18256 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__A2
timestamp 1669390400
transform -1 0 21056 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2115__B2
timestamp 1669390400
transform 1 0 18816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2116__A2
timestamp 1669390400
transform 1 0 22624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A1
timestamp 1669390400
transform 1 0 22176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2117__A2
timestamp 1669390400
transform 1 0 23184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2118__A1
timestamp 1669390400
transform 1 0 17696 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2119__A1
timestamp 1669390400
transform 1 0 21280 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2120__A1
timestamp 1669390400
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2120__A2
timestamp 1669390400
transform 1 0 29456 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__A2
timestamp 1669390400
transform 1 0 26768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2121__B
timestamp 1669390400
transform 1 0 29904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__A1
timestamp 1669390400
transform 1 0 28000 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2123__A2
timestamp 1669390400
transform 1 0 26320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__A2
timestamp 1669390400
transform 1 0 28224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2124__C
timestamp 1669390400
transform 1 0 25312 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A1
timestamp 1669390400
transform 1 0 26656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2126__A2
timestamp 1669390400
transform 1 0 26208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2127__A1
timestamp 1669390400
transform 1 0 23632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2128__A1
timestamp 1669390400
transform 1 0 25312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2129__A3
timestamp 1669390400
transform 1 0 27776 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2134__I
timestamp 1669390400
transform -1 0 57568 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2135__A1
timestamp 1669390400
transform -1 0 2464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2135__A2
timestamp 1669390400
transform -1 0 2912 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2135__B
timestamp 1669390400
transform -1 0 2016 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__A1
timestamp 1669390400
transform 1 0 3808 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__A2
timestamp 1669390400
transform -1 0 5936 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2136__B2
timestamp 1669390400
transform -1 0 10976 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__A2
timestamp 1669390400
transform 1 0 18032 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2137__B
timestamp 1669390400
transform -1 0 17808 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2138__A2
timestamp 1669390400
transform 1 0 17584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__A1
timestamp 1669390400
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2139__A2
timestamp 1669390400
transform 1 0 28672 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__A1
timestamp 1669390400
transform 1 0 23632 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2140__A2
timestamp 1669390400
transform -1 0 24864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__A2
timestamp 1669390400
transform 1 0 27776 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2141__C
timestamp 1669390400
transform 1 0 23184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A1
timestamp 1669390400
transform -1 0 20048 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2142__A2
timestamp 1669390400
transform -1 0 21952 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2143__B2
timestamp 1669390400
transform -1 0 22736 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2144__A2
timestamp 1669390400
transform 1 0 23184 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2147__A2
timestamp 1669390400
transform 1 0 26656 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2148__A2
timestamp 1669390400
transform 1 0 27440 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A1
timestamp 1669390400
transform 1 0 20832 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2156__A2
timestamp 1669390400
transform 1 0 22400 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2157__A2
timestamp 1669390400
transform 1 0 22848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2159__A1
timestamp 1669390400
transform 1 0 20832 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__A1
timestamp 1669390400
transform -1 0 25984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__A2
timestamp 1669390400
transform -1 0 26432 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2160__B
timestamp 1669390400
transform 1 0 28000 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2161__A1
timestamp 1669390400
transform 1 0 27664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2162__A2
timestamp 1669390400
transform -1 0 20496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A1
timestamp 1669390400
transform 1 0 20832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__A2
timestamp 1669390400
transform 1 0 22960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2163__C
timestamp 1669390400
transform 1 0 22736 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2165__A1
timestamp 1669390400
transform 1 0 24080 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2166__A1
timestamp 1669390400
transform 1 0 23184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2168__A1
timestamp 1669390400
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2170__A2
timestamp 1669390400
transform -1 0 26880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2173__I
timestamp 1669390400
transform -1 0 3360 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2178__A1
timestamp 1669390400
transform 1 0 21168 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2180__A1
timestamp 1669390400
transform 1 0 19936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2181__B
timestamp 1669390400
transform -1 0 26208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2184__I
timestamp 1669390400
transform 1 0 51184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2185__A2
timestamp 1669390400
transform 1 0 51184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__A1
timestamp 1669390400
transform 1 0 53984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2190__B
timestamp 1669390400
transform 1 0 55328 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A1
timestamp 1669390400
transform 1 0 47264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2191__A2
timestamp 1669390400
transform -1 0 44912 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2192__A1
timestamp 1669390400
transform 1 0 46704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2193__I
timestamp 1669390400
transform 1 0 49952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2195__I
timestamp 1669390400
transform 1 0 52640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2196__I
timestamp 1669390400
transform 1 0 48720 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2198__I
timestamp 1669390400
transform -1 0 52192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2200__A1
timestamp 1669390400
transform 1 0 49392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2202__I
timestamp 1669390400
transform 1 0 48496 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A1
timestamp 1669390400
transform 1 0 44688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A2
timestamp 1669390400
transform -1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2203__A3
timestamp 1669390400
transform 1 0 44688 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2204__A1
timestamp 1669390400
transform -1 0 52864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2204__A2
timestamp 1669390400
transform 1 0 53312 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A1
timestamp 1669390400
transform -1 0 42784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2207__A2
timestamp 1669390400
transform 1 0 43008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A1
timestamp 1669390400
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A2
timestamp 1669390400
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2208__A3
timestamp 1669390400
transform 1 0 49168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2210__I
timestamp 1669390400
transform 1 0 58016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2211__B
timestamp 1669390400
transform -1 0 44240 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A1
timestamp 1669390400
transform 1 0 50736 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2214__A2
timestamp 1669390400
transform 1 0 51184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2216__I
timestamp 1669390400
transform -1 0 58016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__A1
timestamp 1669390400
transform -1 0 44128 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2219__A2
timestamp 1669390400
transform -1 0 43680 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2220__I
timestamp 1669390400
transform 1 0 57568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2223__I
timestamp 1669390400
transform 1 0 36288 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2224__A1
timestamp 1669390400
transform 1 0 47264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2225__A1
timestamp 1669390400
transform -1 0 47040 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2228__I
timestamp 1669390400
transform 1 0 54544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2233__A1
timestamp 1669390400
transform 1 0 50288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2233__A2
timestamp 1669390400
transform 1 0 51184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2234__A1
timestamp 1669390400
transform -1 0 47936 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__A1
timestamp 1669390400
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__B1
timestamp 1669390400
transform 1 0 44688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2235__B2
timestamp 1669390400
transform 1 0 48160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A1
timestamp 1669390400
transform 1 0 51296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2236__A2
timestamp 1669390400
transform 1 0 57792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2237__I
timestamp 1669390400
transform 1 0 51296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__A1
timestamp 1669390400
transform 1 0 35952 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__A2
timestamp 1669390400
transform -1 0 36288 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2238__B2
timestamp 1669390400
transform 1 0 36512 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2239__A1
timestamp 1669390400
transform 1 0 36512 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__A1
timestamp 1669390400
transform 1 0 39648 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2241__A2
timestamp 1669390400
transform -1 0 39424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__A1
timestamp 1669390400
transform 1 0 46256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__A2
timestamp 1669390400
transform 1 0 46480 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2244__B
timestamp 1669390400
transform 1 0 47600 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2247__I
timestamp 1669390400
transform 1 0 50288 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__A1
timestamp 1669390400
transform 1 0 47712 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__A2
timestamp 1669390400
transform -1 0 46816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2248__B
timestamp 1669390400
transform 1 0 47040 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2249__I
timestamp 1669390400
transform 1 0 58016 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2250__I
timestamp 1669390400
transform 1 0 53872 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A1
timestamp 1669390400
transform 1 0 50624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2253__A2
timestamp 1669390400
transform 1 0 51072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2254__A1
timestamp 1669390400
transform -1 0 53872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2255__I
timestamp 1669390400
transform 1 0 55552 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__A2
timestamp 1669390400
transform 1 0 50288 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__B2
timestamp 1669390400
transform 1 0 49616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2257__C
timestamp 1669390400
transform 1 0 47376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2258__I
timestamp 1669390400
transform 1 0 54432 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2259__I
timestamp 1669390400
transform -1 0 44016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2260__I
timestamp 1669390400
transform 1 0 43344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2261__I
timestamp 1669390400
transform 1 0 44240 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__A1
timestamp 1669390400
transform -1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2262__A2
timestamp 1669390400
transform 1 0 44688 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__A2
timestamp 1669390400
transform 1 0 45472 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2263__B
timestamp 1669390400
transform 1 0 44352 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A1
timestamp 1669390400
transform -1 0 46368 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__A2
timestamp 1669390400
transform 1 0 49392 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2264__C
timestamp 1669390400
transform -1 0 47712 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2265__I
timestamp 1669390400
transform 1 0 56560 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2266__I
timestamp 1669390400
transform 1 0 53312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2267__I
timestamp 1669390400
transform 1 0 57568 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2268__A3
timestamp 1669390400
transform -1 0 57568 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2269__A2
timestamp 1669390400
transform 1 0 54208 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2270__A1
timestamp 1669390400
transform -1 0 57456 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2270__A2
timestamp 1669390400
transform 1 0 57792 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2271__I
timestamp 1669390400
transform -1 0 44912 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2273__I
timestamp 1669390400
transform 1 0 46368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2274__A2
timestamp 1669390400
transform 1 0 47152 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2277__I
timestamp 1669390400
transform -1 0 38416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2278__I
timestamp 1669390400
transform 1 0 57344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__A1
timestamp 1669390400
transform 1 0 50176 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__A2
timestamp 1669390400
transform 1 0 41888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2280__B
timestamp 1669390400
transform 1 0 45584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2281__B1
timestamp 1669390400
transform -1 0 46480 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A1
timestamp 1669390400
transform 1 0 46816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A2
timestamp 1669390400
transform 1 0 47264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__A3
timestamp 1669390400
transform 1 0 48496 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2282__B1
timestamp 1669390400
transform 1 0 47712 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2283__I
timestamp 1669390400
transform 1 0 48608 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2287__A2
timestamp 1669390400
transform -1 0 55216 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2288__A2
timestamp 1669390400
transform 1 0 55104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A1
timestamp 1669390400
transform 1 0 52080 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2290__A2
timestamp 1669390400
transform 1 0 52528 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A1
timestamp 1669390400
transform 1 0 57792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__A2
timestamp 1669390400
transform 1 0 55664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__B1
timestamp 1669390400
transform 1 0 56112 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2291__B2
timestamp 1669390400
transform 1 0 56672 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2294__A2
timestamp 1669390400
transform 1 0 56224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__A1
timestamp 1669390400
transform -1 0 54768 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__A2
timestamp 1669390400
transform 1 0 55888 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2296__B
timestamp 1669390400
transform -1 0 55664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A1
timestamp 1669390400
transform -1 0 58016 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2298__A2
timestamp 1669390400
transform -1 0 57344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__A1
timestamp 1669390400
transform 1 0 56560 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2299__A2
timestamp 1669390400
transform -1 0 57344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__A3
timestamp 1669390400
transform -1 0 57232 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2301__B2
timestamp 1669390400
transform -1 0 56672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__A1
timestamp 1669390400
transform 1 0 53312 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__A2
timestamp 1669390400
transform -1 0 53312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2302__B
timestamp 1669390400
transform 1 0 52640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2303__I
timestamp 1669390400
transform -1 0 54320 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2305__A1
timestamp 1669390400
transform -1 0 38304 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2305__A2
timestamp 1669390400
transform -1 0 38752 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2306__A1
timestamp 1669390400
transform 1 0 34832 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2307__A1
timestamp 1669390400
transform 1 0 34384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2308__I
timestamp 1669390400
transform -1 0 3360 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2310__I
timestamp 1669390400
transform 1 0 38304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2311__A2
timestamp 1669390400
transform 1 0 57568 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2314__A1
timestamp 1669390400
transform 1 0 49840 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2314__A2
timestamp 1669390400
transform 1 0 51184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A1
timestamp 1669390400
transform -1 0 47264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2315__A2
timestamp 1669390400
transform 1 0 53760 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2316__I
timestamp 1669390400
transform 1 0 42560 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2317__I
timestamp 1669390400
transform 1 0 38528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A2
timestamp 1669390400
transform 1 0 43456 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2318__A3
timestamp 1669390400
transform 1 0 43008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2319__A1
timestamp 1669390400
transform 1 0 49504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2322__I
timestamp 1669390400
transform -1 0 49616 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A1
timestamp 1669390400
transform 1 0 44576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__A2
timestamp 1669390400
transform -1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2323__B
timestamp 1669390400
transform -1 0 44016 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A1
timestamp 1669390400
transform 1 0 43008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__A2
timestamp 1669390400
transform 1 0 41440 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2326__B
timestamp 1669390400
transform 1 0 42560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2327__I
timestamp 1669390400
transform -1 0 48272 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2328__A1
timestamp 1669390400
transform -1 0 52080 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2328__A2
timestamp 1669390400
transform 1 0 54208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2328__A3
timestamp 1669390400
transform -1 0 54880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2329__I
timestamp 1669390400
transform -1 0 48048 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__B
timestamp 1669390400
transform 1 0 43680 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2330__C
timestamp 1669390400
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2331__I
timestamp 1669390400
transform -1 0 52864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2333__A2
timestamp 1669390400
transform -1 0 42560 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2334__A1
timestamp 1669390400
transform 1 0 44576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A1
timestamp 1669390400
transform 1 0 36288 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__A2
timestamp 1669390400
transform 1 0 36736 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__B1
timestamp 1669390400
transform -1 0 41664 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2335__B2
timestamp 1669390400
transform 1 0 41664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2336__I
timestamp 1669390400
transform 1 0 48720 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2338__I
timestamp 1669390400
transform -1 0 42112 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2339__I
timestamp 1669390400
transform 1 0 45360 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2340__I
timestamp 1669390400
transform 1 0 55104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2341__I
timestamp 1669390400
transform 1 0 50624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__A1
timestamp 1669390400
transform 1 0 54992 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__A2
timestamp 1669390400
transform -1 0 52864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__B
timestamp 1669390400
transform -1 0 55664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2344__C
timestamp 1669390400
transform 1 0 55888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A1
timestamp 1669390400
transform 1 0 52080 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2346__A2
timestamp 1669390400
transform -1 0 51856 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__A2
timestamp 1669390400
transform 1 0 49840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2347__B
timestamp 1669390400
transform -1 0 51856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A1
timestamp 1669390400
transform 1 0 51520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__A2
timestamp 1669390400
transform 1 0 53760 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2348__B
timestamp 1669390400
transform 1 0 51632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A1
timestamp 1669390400
transform 1 0 57568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2350__A2
timestamp 1669390400
transform 1 0 57792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A1
timestamp 1669390400
transform 1 0 56672 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__A2
timestamp 1669390400
transform 1 0 56224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2351__B
timestamp 1669390400
transform 1 0 58016 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2352__I
timestamp 1669390400
transform 1 0 57568 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2353__B
timestamp 1669390400
transform 1 0 58016 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__A2
timestamp 1669390400
transform 1 0 57344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2354__B
timestamp 1669390400
transform 1 0 57792 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2355__A1
timestamp 1669390400
transform 1 0 56560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2356__I
timestamp 1669390400
transform -1 0 55216 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2357__A1
timestamp 1669390400
transform 1 0 54544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2358__A1
timestamp 1669390400
transform -1 0 42784 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2358__A2
timestamp 1669390400
transform -1 0 46256 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A1
timestamp 1669390400
transform 1 0 49952 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2360__A2
timestamp 1669390400
transform 1 0 54320 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2362__I
timestamp 1669390400
transform 1 0 46928 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2363__A1
timestamp 1669390400
transform 1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2363__A2
timestamp 1669390400
transform 1 0 51856 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2364__I
timestamp 1669390400
transform 1 0 53312 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__A1
timestamp 1669390400
transform 1 0 45360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__A2
timestamp 1669390400
transform 1 0 45808 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2365__A3
timestamp 1669390400
transform 1 0 45808 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2367__A1
timestamp 1669390400
transform 1 0 48272 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2367__A2
timestamp 1669390400
transform 1 0 54656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2369__I
timestamp 1669390400
transform 1 0 42224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__B2
timestamp 1669390400
transform 1 0 43568 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2371__C
timestamp 1669390400
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2372__I
timestamp 1669390400
transform 1 0 57680 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2373__I
timestamp 1669390400
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2375__I
timestamp 1669390400
transform 1 0 39760 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2376__A1
timestamp 1669390400
transform -1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2376__A2
timestamp 1669390400
transform -1 0 55776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A1
timestamp 1669390400
transform 1 0 46704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__A2
timestamp 1669390400
transform 1 0 48720 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2379__B
timestamp 1669390400
transform 1 0 46256 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__A2
timestamp 1669390400
transform 1 0 40992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2380__B
timestamp 1669390400
transform 1 0 44016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__A2
timestamp 1669390400
transform 1 0 43232 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2381__A3
timestamp 1669390400
transform 1 0 42784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__A1
timestamp 1669390400
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__B
timestamp 1669390400
transform 1 0 44016 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2382__C
timestamp 1669390400
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A1
timestamp 1669390400
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2384__A2
timestamp 1669390400
transform 1 0 47824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2385__A1
timestamp 1669390400
transform 1 0 54208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2388__I
timestamp 1669390400
transform -1 0 54320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2389__A1
timestamp 1669390400
transform 1 0 50848 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2389__A2
timestamp 1669390400
transform 1 0 53760 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2389__B
timestamp 1669390400
transform -1 0 52864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__A1
timestamp 1669390400
transform -1 0 54992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__A2
timestamp 1669390400
transform 1 0 53760 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2390__B
timestamp 1669390400
transform 1 0 55216 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A1
timestamp 1669390400
transform 1 0 44576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2391__A2
timestamp 1669390400
transform -1 0 48272 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__A1
timestamp 1669390400
transform 1 0 46256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2392__A3
timestamp 1669390400
transform -1 0 45584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__A2
timestamp 1669390400
transform -1 0 42224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2393__A3
timestamp 1669390400
transform 1 0 42448 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2394__A2
timestamp 1669390400
transform 1 0 45360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2394__B
timestamp 1669390400
transform 1 0 45584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A1
timestamp 1669390400
transform 1 0 45472 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2395__A2
timestamp 1669390400
transform 1 0 45136 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__A2
timestamp 1669390400
transform -1 0 45808 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__B1
timestamp 1669390400
transform 1 0 46144 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2396__B2
timestamp 1669390400
transform 1 0 44576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2397__A1
timestamp 1669390400
transform -1 0 45136 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A1
timestamp 1669390400
transform 1 0 46144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__A2
timestamp 1669390400
transform 1 0 46592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__B
timestamp 1669390400
transform -1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2400__C
timestamp 1669390400
transform 1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2401__A1
timestamp 1669390400
transform 1 0 47936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2402__A2
timestamp 1669390400
transform 1 0 50400 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2402__B
timestamp 1669390400
transform 1 0 49392 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__A1
timestamp 1669390400
transform 1 0 47152 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2403__B
timestamp 1669390400
transform -1 0 48272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2404__A1
timestamp 1669390400
transform 1 0 51968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__A1
timestamp 1669390400
transform 1 0 50736 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__A2
timestamp 1669390400
transform -1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2407__B
timestamp 1669390400
transform 1 0 54320 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A1
timestamp 1669390400
transform -1 0 50512 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A2
timestamp 1669390400
transform -1 0 49504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2408__A3
timestamp 1669390400
transform 1 0 50624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2409__A1
timestamp 1669390400
transform -1 0 50400 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2411__A2
timestamp 1669390400
transform 1 0 32592 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2412__A1
timestamp 1669390400
transform -1 0 35616 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2413__A2
timestamp 1669390400
transform 1 0 38304 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A1
timestamp 1669390400
transform 1 0 41440 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2416__A3
timestamp 1669390400
transform -1 0 44016 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2419__B
timestamp 1669390400
transform -1 0 52192 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__A1
timestamp 1669390400
transform -1 0 49952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__A2
timestamp 1669390400
transform -1 0 47152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2420__B2
timestamp 1669390400
transform 1 0 50288 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__A1
timestamp 1669390400
transform 1 0 51856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__A2
timestamp 1669390400
transform 1 0 52304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2421__B
timestamp 1669390400
transform -1 0 51184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A1
timestamp 1669390400
transform 1 0 49392 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2422__A2
timestamp 1669390400
transform 1 0 48720 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A1
timestamp 1669390400
transform 1 0 52416 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__A2
timestamp 1669390400
transform 1 0 52080 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__B1
timestamp 1669390400
transform -1 0 32592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2423__B2
timestamp 1669390400
transform 1 0 52976 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__A1
timestamp 1669390400
transform 1 0 55776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2425__B
timestamp 1669390400
transform 1 0 56672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A1
timestamp 1669390400
transform -1 0 56672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2426__A3
timestamp 1669390400
transform 1 0 56448 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2427__A1
timestamp 1669390400
transform -1 0 52416 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2427__A2
timestamp 1669390400
transform 1 0 54208 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2427__A3
timestamp 1669390400
transform -1 0 54096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2427__A4
timestamp 1669390400
transform 1 0 53312 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A1
timestamp 1669390400
transform -1 0 55440 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2428__A2
timestamp 1669390400
transform 1 0 54768 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2429__A1
timestamp 1669390400
transform 1 0 51632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2430__I
timestamp 1669390400
transform -1 0 50848 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2433__A1
timestamp 1669390400
transform 1 0 57344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2433__A2
timestamp 1669390400
transform 1 0 54320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__A2
timestamp 1669390400
transform 1 0 55664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2435__B
timestamp 1669390400
transform 1 0 53648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__A1
timestamp 1669390400
transform 1 0 55552 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2436__A2
timestamp 1669390400
transform -1 0 53536 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A1
timestamp 1669390400
transform 1 0 49840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2439__A2
timestamp 1669390400
transform -1 0 49616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A1
timestamp 1669390400
transform 1 0 56224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A2
timestamp 1669390400
transform -1 0 53872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__A3
timestamp 1669390400
transform 1 0 54432 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2441__B
timestamp 1669390400
transform 1 0 56560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A1
timestamp 1669390400
transform -1 0 53312 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A2
timestamp 1669390400
transform 1 0 54768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A3
timestamp 1669390400
transform 1 0 55664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2442__A4
timestamp 1669390400
transform 1 0 55216 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A1
timestamp 1669390400
transform 1 0 56560 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2443__A3
timestamp 1669390400
transform -1 0 54208 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A1
timestamp 1669390400
transform -1 0 57120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__A2
timestamp 1669390400
transform 1 0 57792 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2444__B
timestamp 1669390400
transform 1 0 57344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__A1
timestamp 1669390400
transform 1 0 56336 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2445__B2
timestamp 1669390400
transform -1 0 56336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2446__I
timestamp 1669390400
transform -1 0 51408 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2447__A1
timestamp 1669390400
transform 1 0 33600 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2448__A1
timestamp 1669390400
transform -1 0 40432 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2448__A2
timestamp 1669390400
transform -1 0 40880 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2449__A2
timestamp 1669390400
transform -1 0 47936 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A1
timestamp 1669390400
transform 1 0 50960 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2450__A2
timestamp 1669390400
transform 1 0 48720 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2451__A2
timestamp 1669390400
transform -1 0 46480 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__A1
timestamp 1669390400
transform 1 0 36848 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2454__B
timestamp 1669390400
transform 1 0 36064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2455__A1
timestamp 1669390400
transform -1 0 34496 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2456__A1
timestamp 1669390400
transform 1 0 51632 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2456__A2
timestamp 1669390400
transform -1 0 50960 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2456__B
timestamp 1669390400
transform 1 0 51632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__A1
timestamp 1669390400
transform -1 0 51632 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__B
timestamp 1669390400
transform 1 0 57792 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2457__C
timestamp 1669390400
transform 1 0 55552 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2458__A1
timestamp 1669390400
transform 1 0 54656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2458__A2
timestamp 1669390400
transform -1 0 54432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A1
timestamp 1669390400
transform -1 0 52416 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__A2
timestamp 1669390400
transform 1 0 51744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__B
timestamp 1669390400
transform -1 0 54432 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2459__C
timestamp 1669390400
transform 1 0 50400 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2460__A1
timestamp 1669390400
transform -1 0 40992 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2460__A2
timestamp 1669390400
transform 1 0 40208 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2461__A1
timestamp 1669390400
transform 1 0 56560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2461__A2
timestamp 1669390400
transform 1 0 47712 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2461__C
timestamp 1669390400
transform 1 0 57904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2463__A2
timestamp 1669390400
transform -1 0 35280 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2464__A4
timestamp 1669390400
transform 1 0 45360 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__A1
timestamp 1669390400
transform -1 0 42560 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2465__B
timestamp 1669390400
transform -1 0 44464 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2470__I
timestamp 1669390400
transform 1 0 3136 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__A1
timestamp 1669390400
transform 1 0 41328 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2473__A3
timestamp 1669390400
transform 1 0 40880 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__A1
timestamp 1669390400
transform -1 0 51744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2475__B2
timestamp 1669390400
transform -1 0 50848 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2476__A1
timestamp 1669390400
transform 1 0 51072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2477__A1
timestamp 1669390400
transform -1 0 49952 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2478__A1
timestamp 1669390400
transform 1 0 47264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2478__A2
timestamp 1669390400
transform 1 0 47040 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A1
timestamp 1669390400
transform -1 0 47936 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2479__A2
timestamp 1669390400
transform -1 0 31920 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2480__A1
timestamp 1669390400
transform 1 0 49056 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2480__A2
timestamp 1669390400
transform 1 0 49504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A1
timestamp 1669390400
transform 1 0 47600 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__A2
timestamp 1669390400
transform 1 0 56560 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2481__B
timestamp 1669390400
transform 1 0 54208 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A1
timestamp 1669390400
transform 1 0 53312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2483__A2
timestamp 1669390400
transform -1 0 51408 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A1
timestamp 1669390400
transform 1 0 52528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2484__A2
timestamp 1669390400
transform -1 0 53648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2485__I
timestamp 1669390400
transform 1 0 54656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A1
timestamp 1669390400
transform 1 0 57568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__A2
timestamp 1669390400
transform -1 0 53648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__B
timestamp 1669390400
transform 1 0 56672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2486__C
timestamp 1669390400
transform 1 0 58016 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__A1
timestamp 1669390400
transform 1 0 56672 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2487__C
timestamp 1669390400
transform 1 0 57120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A1
timestamp 1669390400
transform 1 0 51296 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A2
timestamp 1669390400
transform 1 0 52192 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2488__A3
timestamp 1669390400
transform 1 0 54768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2489__A3
timestamp 1669390400
transform 1 0 57456 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2490__A1
timestamp 1669390400
transform 1 0 57008 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2492__A1
timestamp 1669390400
transform 1 0 43904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2492__A2
timestamp 1669390400
transform -1 0 43680 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A1
timestamp 1669390400
transform 1 0 44016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2493__A2
timestamp 1669390400
transform -1 0 41328 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2494__A1
timestamp 1669390400
transform -1 0 53760 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2494__A2
timestamp 1669390400
transform 1 0 57344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__A1
timestamp 1669390400
transform -1 0 55888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2495__B
timestamp 1669390400
transform 1 0 57792 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2496__B
timestamp 1669390400
transform 1 0 57792 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2497__I
timestamp 1669390400
transform -1 0 52864 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A1
timestamp 1669390400
transform 1 0 53200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2498__A2
timestamp 1669390400
transform 1 0 57680 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__A2
timestamp 1669390400
transform -1 0 52752 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2499__B
timestamp 1669390400
transform 1 0 53312 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2500__A2
timestamp 1669390400
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__A1
timestamp 1669390400
transform 1 0 57792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__A2
timestamp 1669390400
transform 1 0 53312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2501__B
timestamp 1669390400
transform 1 0 54656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2502__A1
timestamp 1669390400
transform 1 0 54656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2503__I
timestamp 1669390400
transform -1 0 53984 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A1
timestamp 1669390400
transform -1 0 45696 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2504__A2
timestamp 1669390400
transform 1 0 48832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A1
timestamp 1669390400
transform -1 0 50960 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2508__A2
timestamp 1669390400
transform -1 0 48720 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2509__B
timestamp 1669390400
transform 1 0 48608 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__A2
timestamp 1669390400
transform 1 0 41888 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__B1
timestamp 1669390400
transform 1 0 41216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2510__B2
timestamp 1669390400
transform 1 0 42336 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A2
timestamp 1669390400
transform 1 0 41440 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A3
timestamp 1669390400
transform 1 0 44128 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2511__A4
timestamp 1669390400
transform -1 0 43008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__A1
timestamp 1669390400
transform 1 0 43344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__A2
timestamp 1669390400
transform 1 0 39648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2512__B
timestamp 1669390400
transform 1 0 41440 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__A2
timestamp 1669390400
transform 1 0 41888 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2513__B
timestamp 1669390400
transform 1 0 42336 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__A1
timestamp 1669390400
transform -1 0 52976 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__A2
timestamp 1669390400
transform -1 0 51632 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__B2
timestamp 1669390400
transform 1 0 53760 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2514__C
timestamp 1669390400
transform 1 0 53200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2515__B
timestamp 1669390400
transform 1 0 48160 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A1
timestamp 1669390400
transform 1 0 50848 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2516__A2
timestamp 1669390400
transform 1 0 50736 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__A1
timestamp 1669390400
transform -1 0 41664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2517__A2
timestamp 1669390400
transform 1 0 42672 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__A1
timestamp 1669390400
transform -1 0 42672 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__A2
timestamp 1669390400
transform 1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__B1
timestamp 1669390400
transform 1 0 43456 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2518__C
timestamp 1669390400
transform 1 0 47264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2519__A1
timestamp 1669390400
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2520__A2
timestamp 1669390400
transform 1 0 32816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2521__A1
timestamp 1669390400
transform -1 0 34832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2522__A4
timestamp 1669390400
transform -1 0 38976 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2523__A1
timestamp 1669390400
transform 1 0 41664 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2523__B
timestamp 1669390400
transform -1 0 39424 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__A1
timestamp 1669390400
transform 1 0 45024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__A2
timestamp 1669390400
transform -1 0 41664 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__A3
timestamp 1669390400
transform -1 0 42112 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2529__A4
timestamp 1669390400
transform 1 0 44576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2531__A3
timestamp 1669390400
transform 1 0 51296 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__A1
timestamp 1669390400
transform -1 0 52528 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2532__B
timestamp 1669390400
transform -1 0 54880 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2533__A2
timestamp 1669390400
transform -1 0 51296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__A2
timestamp 1669390400
transform -1 0 49504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2535__B
timestamp 1669390400
transform 1 0 50624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A2
timestamp 1669390400
transform 1 0 56560 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2536__A3
timestamp 1669390400
transform -1 0 53312 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A1
timestamp 1669390400
transform 1 0 52640 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A2
timestamp 1669390400
transform -1 0 53424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2537__A3
timestamp 1669390400
transform 1 0 50624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2538__A1
timestamp 1669390400
transform -1 0 50400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A1
timestamp 1669390400
transform 1 0 50176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__A2
timestamp 1669390400
transform -1 0 50960 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2539__B
timestamp 1669390400
transform 1 0 50736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__A2
timestamp 1669390400
transform 1 0 56560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2540__B
timestamp 1669390400
transform 1 0 55104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__A1
timestamp 1669390400
transform 1 0 57904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2541__B
timestamp 1669390400
transform -1 0 51296 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A1
timestamp 1669390400
transform 1 0 45920 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2543__A2
timestamp 1669390400
transform 1 0 48384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2544__I
timestamp 1669390400
transform -1 0 42336 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__A1
timestamp 1669390400
transform 1 0 46816 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2545__A2
timestamp 1669390400
transform -1 0 49616 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__A1
timestamp 1669390400
transform -1 0 50512 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2546__B
timestamp 1669390400
transform -1 0 50064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__A1
timestamp 1669390400
transform 1 0 58016 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__A2
timestamp 1669390400
transform 1 0 52304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2547__A3
timestamp 1669390400
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A1
timestamp 1669390400
transform -1 0 49616 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2548__A2
timestamp 1669390400
transform 1 0 53312 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__A2
timestamp 1669390400
transform -1 0 47824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2549__B
timestamp 1669390400
transform 1 0 52416 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2550__A2
timestamp 1669390400
transform 1 0 57344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__A1
timestamp 1669390400
transform -1 0 58016 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2551__A3
timestamp 1669390400
transform 1 0 57344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2552__A1
timestamp 1669390400
transform 1 0 51408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__A1
timestamp 1669390400
transform 1 0 51184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__A2
timestamp 1669390400
transform 1 0 54656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2553__B
timestamp 1669390400
transform 1 0 54208 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2554__S
timestamp 1669390400
transform -1 0 50512 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A1
timestamp 1669390400
transform 1 0 55216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A2
timestamp 1669390400
transform 1 0 55664 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2555__A3
timestamp 1669390400
transform 1 0 54208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2558__A2
timestamp 1669390400
transform -1 0 42336 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2559__I
timestamp 1669390400
transform 1 0 44912 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2560__I
timestamp 1669390400
transform 1 0 41440 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__A1
timestamp 1669390400
transform 1 0 46144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__A2
timestamp 1669390400
transform -1 0 32592 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2561__B
timestamp 1669390400
transform 1 0 43456 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A1
timestamp 1669390400
transform -1 0 46144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2562__A3
timestamp 1669390400
transform -1 0 47488 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__A1
timestamp 1669390400
transform 1 0 48272 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2563__A2
timestamp 1669390400
transform -1 0 46032 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2564__A2
timestamp 1669390400
transform 1 0 48272 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__A2
timestamp 1669390400
transform 1 0 53312 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2565__B
timestamp 1669390400
transform 1 0 51520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2566__I
timestamp 1669390400
transform -1 0 46592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2567__A1
timestamp 1669390400
transform 1 0 51856 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2568__A2
timestamp 1669390400
transform 1 0 46704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__A1
timestamp 1669390400
transform 1 0 46592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2570__A2
timestamp 1669390400
transform -1 0 45584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2571__C
timestamp 1669390400
transform 1 0 47040 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__A1
timestamp 1669390400
transform 1 0 51072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2572__A2
timestamp 1669390400
transform 1 0 51968 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__A1
timestamp 1669390400
transform 1 0 46144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2573__A2
timestamp 1669390400
transform -1 0 45584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2577__B
timestamp 1669390400
transform -1 0 44912 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2579__A1
timestamp 1669390400
transform 1 0 53760 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__A1
timestamp 1669390400
transform 1 0 49728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2580__C
timestamp 1669390400
transform 1 0 51744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2581__A1
timestamp 1669390400
transform -1 0 49616 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A1
timestamp 1669390400
transform 1 0 52192 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2582__A3
timestamp 1669390400
transform 1 0 51184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2584__A1
timestamp 1669390400
transform 1 0 44352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__A1
timestamp 1669390400
transform -1 0 46144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__A2
timestamp 1669390400
transform -1 0 45248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2585__B
timestamp 1669390400
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__A1
timestamp 1669390400
transform 1 0 45360 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2586__A2
timestamp 1669390400
transform 1 0 48720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__A2
timestamp 1669390400
transform -1 0 39872 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2587__A3
timestamp 1669390400
transform 1 0 40432 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2588__I
timestamp 1669390400
transform 1 0 38304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A1
timestamp 1669390400
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A2
timestamp 1669390400
transform 1 0 47152 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2589__A3
timestamp 1669390400
transform 1 0 41664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A1
timestamp 1669390400
transform -1 0 36512 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__A2
timestamp 1669390400
transform -1 0 33040 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2590__B
timestamp 1669390400
transform 1 0 36624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__A1
timestamp 1669390400
transform -1 0 32592 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__A2
timestamp 1669390400
transform 1 0 38640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2591__A3
timestamp 1669390400
transform 1 0 37072 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__A1
timestamp 1669390400
transform 1 0 37520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2592__A2
timestamp 1669390400
transform 1 0 37408 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2593__I
timestamp 1669390400
transform 1 0 43344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2594__A1
timestamp 1669390400
transform -1 0 38304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__A1
timestamp 1669390400
transform 1 0 39536 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2595__B
timestamp 1669390400
transform -1 0 39312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2596__I
timestamp 1669390400
transform 1 0 34384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__A1
timestamp 1669390400
transform -1 0 38528 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2597__C
timestamp 1669390400
transform 1 0 37968 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__A2
timestamp 1669390400
transform 1 0 34944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2599__A3
timestamp 1669390400
transform 1 0 35168 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2600__A1
timestamp 1669390400
transform -1 0 34944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2601__A3
timestamp 1669390400
transform 1 0 34720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__A1
timestamp 1669390400
transform -1 0 35728 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2607__A2
timestamp 1669390400
transform 1 0 35952 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2609__I
timestamp 1669390400
transform 1 0 34608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__A1
timestamp 1669390400
transform 1 0 45472 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2610__B
timestamp 1669390400
transform 1 0 45024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A1
timestamp 1669390400
transform -1 0 37520 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A2
timestamp 1669390400
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__A3
timestamp 1669390400
transform 1 0 35616 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2611__B
timestamp 1669390400
transform -1 0 37072 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2612__I
timestamp 1669390400
transform 1 0 42896 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2613__I
timestamp 1669390400
transform -1 0 43008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__A1
timestamp 1669390400
transform 1 0 41440 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__A2
timestamp 1669390400
transform 1 0 46144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2614__B
timestamp 1669390400
transform 1 0 46592 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2616__I
timestamp 1669390400
transform 1 0 42336 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2617__A2
timestamp 1669390400
transform 1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__A1
timestamp 1669390400
transform 1 0 41216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__A2
timestamp 1669390400
transform 1 0 42784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2618__A3
timestamp 1669390400
transform 1 0 39984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__A1
timestamp 1669390400
transform 1 0 40320 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2619__A2
timestamp 1669390400
transform 1 0 40768 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2620__A1
timestamp 1669390400
transform 1 0 41888 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A1
timestamp 1669390400
transform -1 0 41664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2621__A3
timestamp 1669390400
transform -1 0 40768 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__A1
timestamp 1669390400
transform 1 0 41888 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__A2
timestamp 1669390400
transform -1 0 41664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2622__A3
timestamp 1669390400
transform 1 0 43232 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__A1
timestamp 1669390400
transform -1 0 51968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__A2
timestamp 1669390400
transform -1 0 51632 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2624__A3
timestamp 1669390400
transform -1 0 52192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__A1
timestamp 1669390400
transform 1 0 56112 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__A2
timestamp 1669390400
transform 1 0 56000 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2625__A3
timestamp 1669390400
transform 1 0 53200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__A3
timestamp 1669390400
transform -1 0 53872 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2626__B
timestamp 1669390400
transform 1 0 56448 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2627__A1
timestamp 1669390400
transform 1 0 50848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__A1
timestamp 1669390400
transform 1 0 48608 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2629__A2
timestamp 1669390400
transform -1 0 48384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2630__C
timestamp 1669390400
transform 1 0 47936 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2631__A1
timestamp 1669390400
transform -1 0 49392 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2632__I
timestamp 1669390400
transform 1 0 50736 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2633__B
timestamp 1669390400
transform 1 0 50736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__A1
timestamp 1669390400
transform -1 0 48832 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2634__A2
timestamp 1669390400
transform -1 0 48496 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2636__B
timestamp 1669390400
transform 1 0 46480 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A1
timestamp 1669390400
transform 1 0 32032 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2637__A2
timestamp 1669390400
transform 1 0 32480 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A1
timestamp 1669390400
transform 1 0 39760 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__A2
timestamp 1669390400
transform 1 0 40768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__B1
timestamp 1669390400
transform 1 0 39312 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__B2
timestamp 1669390400
transform 1 0 38864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2638__C
timestamp 1669390400
transform -1 0 41328 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__A1
timestamp 1669390400
transform 1 0 37408 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2639__A2
timestamp 1669390400
transform 1 0 37408 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__A2
timestamp 1669390400
transform 1 0 39088 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2640__B
timestamp 1669390400
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__A1
timestamp 1669390400
transform 1 0 38752 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2641__B
timestamp 1669390400
transform 1 0 38752 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2642__A1
timestamp 1669390400
transform 1 0 36400 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A2
timestamp 1669390400
transform -1 0 38976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A3
timestamp 1669390400
transform 1 0 39200 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2644__A4
timestamp 1669390400
transform 1 0 41216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2646__A1
timestamp 1669390400
transform -1 0 30800 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2647__A3
timestamp 1669390400
transform 1 0 31808 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__A1
timestamp 1669390400
transform 1 0 38304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__A2
timestamp 1669390400
transform 1 0 37408 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__A3
timestamp 1669390400
transform 1 0 37856 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2648__A4
timestamp 1669390400
transform 1 0 35168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__A1
timestamp 1669390400
transform 1 0 37408 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__A2
timestamp 1669390400
transform 1 0 37856 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__A3
timestamp 1669390400
transform 1 0 38304 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2649__B
timestamp 1669390400
transform -1 0 36624 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2653__I
timestamp 1669390400
transform 1 0 57904 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2654__A1
timestamp 1669390400
transform -1 0 48048 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__A2
timestamp 1669390400
transform -1 0 29680 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2655__B
timestamp 1669390400
transform -1 0 31472 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2656__I
timestamp 1669390400
transform 1 0 39536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2658__A1
timestamp 1669390400
transform -1 0 52976 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2658__A4
timestamp 1669390400
transform 1 0 51520 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2659__I
timestamp 1669390400
transform 1 0 33488 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__A1
timestamp 1669390400
transform -1 0 35840 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__A2
timestamp 1669390400
transform 1 0 35840 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2660__A3
timestamp 1669390400
transform 1 0 35168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A1
timestamp 1669390400
transform 1 0 38976 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2661__A2
timestamp 1669390400
transform 1 0 38528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A1
timestamp 1669390400
transform 1 0 38528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2662__A3
timestamp 1669390400
transform 1 0 42000 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2663__I
timestamp 1669390400
transform 1 0 39648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__A1
timestamp 1669390400
transform 1 0 39424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__A2
timestamp 1669390400
transform 1 0 38864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__B1
timestamp 1669390400
transform -1 0 38192 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2664__B2
timestamp 1669390400
transform 1 0 38976 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__A1
timestamp 1669390400
transform 1 0 41440 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2665__A2
timestamp 1669390400
transform 1 0 46032 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2666__I
timestamp 1669390400
transform 1 0 34272 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2667__C
timestamp 1669390400
transform 1 0 37408 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__A1
timestamp 1669390400
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2668__A2
timestamp 1669390400
transform 1 0 38416 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__A1
timestamp 1669390400
transform 1 0 41440 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2669__A2
timestamp 1669390400
transform -1 0 42336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2670__I
timestamp 1669390400
transform 1 0 40208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__A1
timestamp 1669390400
transform -1 0 37632 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2671__A2
timestamp 1669390400
transform 1 0 39984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__A1
timestamp 1669390400
transform -1 0 52080 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2672__A4
timestamp 1669390400
transform 1 0 52528 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2673__A3
timestamp 1669390400
transform -1 0 39984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2674__I
timestamp 1669390400
transform -1 0 34384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__A2
timestamp 1669390400
transform 1 0 41888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2675__A3
timestamp 1669390400
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__A1
timestamp 1669390400
transform 1 0 43456 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__A2
timestamp 1669390400
transform -1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__A3
timestamp 1669390400
transform 1 0 43008 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2676__A4
timestamp 1669390400
transform 1 0 43680 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__A1
timestamp 1669390400
transform -1 0 42336 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__A2
timestamp 1669390400
transform -1 0 44688 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2678__A3
timestamp 1669390400
transform 1 0 42560 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2679__B
timestamp 1669390400
transform -1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__B1
timestamp 1669390400
transform -1 0 44240 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2680__B2
timestamp 1669390400
transform -1 0 42896 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__A2
timestamp 1669390400
transform 1 0 43568 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2681__A4
timestamp 1669390400
transform -1 0 43344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2682__A1
timestamp 1669390400
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__A1
timestamp 1669390400
transform -1 0 47152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2683__A2
timestamp 1669390400
transform 1 0 46480 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2684__C
timestamp 1669390400
transform 1 0 48496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__A1
timestamp 1669390400
transform 1 0 50176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2685__A2
timestamp 1669390400
transform 1 0 48496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2687__A1
timestamp 1669390400
transform 1 0 48048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2688__A1
timestamp 1669390400
transform 1 0 39536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2689__A2
timestamp 1669390400
transform -1 0 41776 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__A1
timestamp 1669390400
transform 1 0 41216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2690__A3
timestamp 1669390400
transform 1 0 43680 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2691__A1
timestamp 1669390400
transform 1 0 48384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2693__A1
timestamp 1669390400
transform 1 0 41664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2694__A1
timestamp 1669390400
transform 1 0 31696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2695__I
timestamp 1669390400
transform 1 0 36624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2696__I
timestamp 1669390400
transform -1 0 36960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__A1
timestamp 1669390400
transform -1 0 40208 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__A2
timestamp 1669390400
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2697__B
timestamp 1669390400
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__B
timestamp 1669390400
transform 1 0 38416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2698__C
timestamp 1669390400
transform 1 0 39312 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2699__A2
timestamp 1669390400
transform 1 0 35280 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2700__I
timestamp 1669390400
transform -1 0 32816 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__A1
timestamp 1669390400
transform 1 0 34944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__A2
timestamp 1669390400
transform -1 0 31472 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2701__B2
timestamp 1669390400
transform 1 0 31920 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2703__A2
timestamp 1669390400
transform 1 0 33040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A1
timestamp 1669390400
transform -1 0 34832 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2705__A3
timestamp 1669390400
transform 1 0 35056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A1
timestamp 1669390400
transform -1 0 33152 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2706__A2
timestamp 1669390400
transform -1 0 33600 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2707__I
timestamp 1669390400
transform 1 0 31696 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__A1
timestamp 1669390400
transform 1 0 34832 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2710__A2
timestamp 1669390400
transform 1 0 35168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__A1
timestamp 1669390400
transform 1 0 34272 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2711__A2
timestamp 1669390400
transform 1 0 34720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2712__A1
timestamp 1669390400
transform 1 0 35952 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2716__I
timestamp 1669390400
transform -1 0 39200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2717__A2
timestamp 1669390400
transform 1 0 32144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2718__I
timestamp 1669390400
transform 1 0 45808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__A1
timestamp 1669390400
transform -1 0 46480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__A2
timestamp 1669390400
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__B1
timestamp 1669390400
transform 1 0 48496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2719__B2
timestamp 1669390400
transform 1 0 47376 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2720__A1
timestamp 1669390400
transform 1 0 50400 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2720__A2
timestamp 1669390400
transform 1 0 50848 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2721__A1
timestamp 1669390400
transform -1 0 43456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__A2
timestamp 1669390400
transform 1 0 44352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2722__A3
timestamp 1669390400
transform 1 0 52080 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__A1
timestamp 1669390400
transform 1 0 51632 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__A2
timestamp 1669390400
transform -1 0 46816 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2724__A3
timestamp 1669390400
transform 1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__A1
timestamp 1669390400
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2726__B2
timestamp 1669390400
transform -1 0 50848 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2727__A2
timestamp 1669390400
transform -1 0 44576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2728__A2
timestamp 1669390400
transform 1 0 45136 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2729__A1
timestamp 1669390400
transform 1 0 36064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__A1
timestamp 1669390400
transform 1 0 38304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2730__A2
timestamp 1669390400
transform 1 0 41776 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2731__I
timestamp 1669390400
transform 1 0 36736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__A1
timestamp 1669390400
transform 1 0 38528 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2732__A2
timestamp 1669390400
transform -1 0 35056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__A1
timestamp 1669390400
transform 1 0 35504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__A2
timestamp 1669390400
transform 1 0 35056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2733__B
timestamp 1669390400
transform 1 0 33936 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2734__B
timestamp 1669390400
transform 1 0 37856 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2735__A1
timestamp 1669390400
transform 1 0 38080 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A1
timestamp 1669390400
transform -1 0 38976 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A2
timestamp 1669390400
transform 1 0 40656 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__A3
timestamp 1669390400
transform -1 0 37744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2736__B
timestamp 1669390400
transform 1 0 41104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2737__A2
timestamp 1669390400
transform 1 0 38304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2739__I
timestamp 1669390400
transform 1 0 35504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__A1
timestamp 1669390400
transform -1 0 33040 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2740__A2
timestamp 1669390400
transform 1 0 37856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__A1
timestamp 1669390400
transform 1 0 33936 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__A2
timestamp 1669390400
transform 1 0 33488 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2741__C
timestamp 1669390400
transform 1 0 32480 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A1
timestamp 1669390400
transform 1 0 34832 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A2
timestamp 1669390400
transform -1 0 32368 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A3
timestamp 1669390400
transform 1 0 36176 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2743__A4
timestamp 1669390400
transform -1 0 34384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2744__A1
timestamp 1669390400
transform 1 0 33488 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__A1
timestamp 1669390400
transform 1 0 32256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2746__A3
timestamp 1669390400
transform 1 0 33488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2747__A1
timestamp 1669390400
transform 1 0 33936 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2747__B
timestamp 1669390400
transform -1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2754__I
timestamp 1669390400
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2757__A1
timestamp 1669390400
transform -1 0 41664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2757__A2
timestamp 1669390400
transform 1 0 41888 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2757__B
timestamp 1669390400
transform -1 0 41776 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2758__A2
timestamp 1669390400
transform -1 0 43120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2758__A3
timestamp 1669390400
transform 1 0 39872 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2759__A1
timestamp 1669390400
transform 1 0 37968 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2759__C
timestamp 1669390400
transform -1 0 35952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A1
timestamp 1669390400
transform 1 0 42896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2760__A2
timestamp 1669390400
transform 1 0 43344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2761__A1
timestamp 1669390400
transform -1 0 37744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2762__A1
timestamp 1669390400
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2762__A2
timestamp 1669390400
transform 1 0 36176 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A1
timestamp 1669390400
transform 1 0 37856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2763__A2
timestamp 1669390400
transform 1 0 39088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2764__A1
timestamp 1669390400
transform 1 0 41888 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2764__A2
timestamp 1669390400
transform 1 0 47488 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__A1
timestamp 1669390400
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__B
timestamp 1669390400
transform -1 0 40656 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2765__C
timestamp 1669390400
transform 1 0 37408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2766__A1
timestamp 1669390400
transform 1 0 45360 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2766__A2
timestamp 1669390400
transform 1 0 42224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2767__A2
timestamp 1669390400
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2767__B
timestamp 1669390400
transform 1 0 37408 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2768__A2
timestamp 1669390400
transform -1 0 39984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2770__B
timestamp 1669390400
transform -1 0 41776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2773__A1
timestamp 1669390400
transform 1 0 36960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2773__A2
timestamp 1669390400
transform -1 0 38416 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2774__A1
timestamp 1669390400
transform -1 0 33264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2774__A2
timestamp 1669390400
transform 1 0 33488 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2775__A1
timestamp 1669390400
transform -1 0 34944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2776__I
timestamp 1669390400
transform 1 0 37968 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2777__A1
timestamp 1669390400
transform 1 0 37072 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2777__A2
timestamp 1669390400
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2777__B
timestamp 1669390400
transform 1 0 37520 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2778__A1
timestamp 1669390400
transform 1 0 32704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2780__A1
timestamp 1669390400
transform -1 0 28224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2781__B1
timestamp 1669390400
transform 1 0 39984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2781__B2
timestamp 1669390400
transform -1 0 35504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2783__A2
timestamp 1669390400
transform 1 0 32256 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2785__A2
timestamp 1669390400
transform -1 0 30128 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2791__I
timestamp 1669390400
transform 1 0 3136 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2793__A2
timestamp 1669390400
transform 1 0 30576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2794__A1
timestamp 1669390400
transform 1 0 49392 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2795__A2
timestamp 1669390400
transform -1 0 40992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2795__A3
timestamp 1669390400
transform 1 0 40880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__A1
timestamp 1669390400
transform -1 0 38528 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__A2
timestamp 1669390400
transform 1 0 38528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__B1
timestamp 1669390400
transform 1 0 38864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2796__B2
timestamp 1669390400
transform 1 0 40320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2797__A1
timestamp 1669390400
transform 1 0 36848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2797__A2
timestamp 1669390400
transform 1 0 37296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__A1
timestamp 1669390400
transform -1 0 38080 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__A2
timestamp 1669390400
transform -1 0 33712 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2798__B
timestamp 1669390400
transform 1 0 34720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2799__A1
timestamp 1669390400
transform -1 0 35168 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2799__A2
timestamp 1669390400
transform 1 0 35392 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2801__I
timestamp 1669390400
transform 1 0 34720 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2803__B
timestamp 1669390400
transform 1 0 36400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2804__A2
timestamp 1669390400
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2805__A1
timestamp 1669390400
transform 1 0 38304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2805__A3
timestamp 1669390400
transform 1 0 38752 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2806__A1
timestamp 1669390400
transform 1 0 35504 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2809__A1
timestamp 1669390400
transform 1 0 31584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2811__A1
timestamp 1669390400
transform 1 0 31696 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2812__A2
timestamp 1669390400
transform -1 0 32480 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2819__I
timestamp 1669390400
transform 1 0 41440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2820__A1
timestamp 1669390400
transform 1 0 50176 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2820__A2
timestamp 1669390400
transform 1 0 50736 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2821__A2
timestamp 1669390400
transform 1 0 38192 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2821__B
timestamp 1669390400
transform 1 0 39536 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2821__C
timestamp 1669390400
transform 1 0 38976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__A1
timestamp 1669390400
transform 1 0 40992 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__B1
timestamp 1669390400
transform -1 0 38080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2822__B2
timestamp 1669390400
transform 1 0 40544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2823__A2
timestamp 1669390400
transform 1 0 54208 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2824__A1
timestamp 1669390400
transform 1 0 55664 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2825__A1
timestamp 1669390400
transform -1 0 35728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2825__A2
timestamp 1669390400
transform 1 0 36960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2827__A1
timestamp 1669390400
transform 1 0 37072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2828__A1
timestamp 1669390400
transform 1 0 40432 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2829__A2
timestamp 1669390400
transform 1 0 57792 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2831__I
timestamp 1669390400
transform 1 0 56112 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2833__A2
timestamp 1669390400
transform 1 0 32704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2835__A2
timestamp 1669390400
transform -1 0 55440 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2841__A2
timestamp 1669390400
transform 1 0 57344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2842__I
timestamp 1669390400
transform -1 0 38192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2843__A1
timestamp 1669390400
transform -1 0 55328 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2843__A3
timestamp 1669390400
transform -1 0 54432 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2845__A1
timestamp 1669390400
transform -1 0 39424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2845__A2
timestamp 1669390400
transform -1 0 40320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2845__B1
timestamp 1669390400
transform 1 0 39648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2845__B2
timestamp 1669390400
transform 1 0 41440 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2846__A2
timestamp 1669390400
transform 1 0 49728 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2847__A1
timestamp 1669390400
transform 1 0 49280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2847__A2
timestamp 1669390400
transform -1 0 48160 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2848__A1
timestamp 1669390400
transform 1 0 50288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2849__A1
timestamp 1669390400
transform 1 0 51184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2849__A2
timestamp 1669390400
transform 1 0 50288 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2850__A1
timestamp 1669390400
transform -1 0 53536 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2850__A2
timestamp 1669390400
transform -1 0 52416 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2852__A2
timestamp 1669390400
transform 1 0 56560 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2853__A2
timestamp 1669390400
transform -1 0 57344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2855__I
timestamp 1669390400
transform -1 0 37744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2857__A1
timestamp 1669390400
transform 1 0 58016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2864__A1
timestamp 1669390400
transform 1 0 56560 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2865__B2
timestamp 1669390400
transform 1 0 57344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2868__A2
timestamp 1669390400
transform -1 0 36960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2869__A1
timestamp 1669390400
transform -1 0 37856 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2869__A2
timestamp 1669390400
transform 1 0 39424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__I0
timestamp 1669390400
transform 1 0 32816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__I1
timestamp 1669390400
transform 1 0 35280 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2870__S
timestamp 1669390400
transform 1 0 35728 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2872__A1
timestamp 1669390400
transform -1 0 33488 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2872__A2
timestamp 1669390400
transform -1 0 33040 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2872__A3
timestamp 1669390400
transform -1 0 33936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2874__A1
timestamp 1669390400
transform 1 0 34608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2875__A1
timestamp 1669390400
transform 1 0 32816 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2876__I
timestamp 1669390400
transform -1 0 37632 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2877__A1
timestamp 1669390400
transform -1 0 37408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2880__A2
timestamp 1669390400
transform -1 0 42336 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2881__A1
timestamp 1669390400
transform -1 0 43232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2881__A2
timestamp 1669390400
transform -1 0 39200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2881__B1
timestamp 1669390400
transform -1 0 43120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2882__A1
timestamp 1669390400
transform 1 0 36736 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2882__A2
timestamp 1669390400
transform 1 0 34832 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2885__A1
timestamp 1669390400
transform -1 0 39312 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2885__C
timestamp 1669390400
transform 1 0 38640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2886__A1
timestamp 1669390400
transform -1 0 35392 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__A1
timestamp 1669390400
transform 1 0 35056 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2888__B
timestamp 1669390400
transform -1 0 35840 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2889__A2
timestamp 1669390400
transform 1 0 36288 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2889__B2
timestamp 1669390400
transform 1 0 34608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2890__I
timestamp 1669390400
transform 1 0 34048 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2891__A1
timestamp 1669390400
transform -1 0 34496 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2891__A2
timestamp 1669390400
transform -1 0 34048 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2891__A4
timestamp 1669390400
transform 1 0 37632 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__A1
timestamp 1669390400
transform 1 0 33936 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__A3
timestamp 1669390400
transform 1 0 34608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2893__A4
timestamp 1669390400
transform 1 0 34720 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2894__A1
timestamp 1669390400
transform 1 0 34496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2894__B
timestamp 1669390400
transform -1 0 35504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2897__A1
timestamp 1669390400
transform 1 0 34272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2898__A1
timestamp 1669390400
transform 1 0 31696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2899__A1
timestamp 1669390400
transform 1 0 31696 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2899__A2
timestamp 1669390400
transform 1 0 31248 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2899__B1
timestamp 1669390400
transform -1 0 29680 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__A1
timestamp 1669390400
transform 1 0 27776 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__A2
timestamp 1669390400
transform 1 0 29904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__B1
timestamp 1669390400
transform 1 0 30912 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2900__B2
timestamp 1669390400
transform 1 0 30352 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2901__A1
timestamp 1669390400
transform 1 0 28784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2901__A2
timestamp 1669390400
transform 1 0 29232 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2901__B1
timestamp 1669390400
transform 1 0 31248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2901__B2
timestamp 1669390400
transform -1 0 29680 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2903__A1
timestamp 1669390400
transform 1 0 30688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2904__A1
timestamp 1669390400
transform -1 0 31808 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2905__A1
timestamp 1669390400
transform 1 0 31808 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2906__A1
timestamp 1669390400
transform -1 0 29008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2906__B2
timestamp 1669390400
transform 1 0 30464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2907__A1
timestamp 1669390400
transform -1 0 5152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2908__A1
timestamp 1669390400
transform 1 0 6384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2909__A1
timestamp 1669390400
transform 1 0 35168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2910__I1
timestamp 1669390400
transform 1 0 35616 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2912__A1
timestamp 1669390400
transform 1 0 38304 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2912__A2
timestamp 1669390400
transform 1 0 39088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2913__A1
timestamp 1669390400
transform -1 0 35168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2914__CLK
timestamp 1669390400
transform -1 0 46816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2914__D
timestamp 1669390400
transform -1 0 40992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2914__RN
timestamp 1669390400
transform 1 0 46144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2915__CLK
timestamp 1669390400
transform -1 0 36960 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2916__CLK
timestamp 1669390400
transform 1 0 37632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2916__D
timestamp 1669390400
transform -1 0 38080 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2917__CLK
timestamp 1669390400
transform 1 0 57008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2917__D
timestamp 1669390400
transform 1 0 57456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2918__CLK
timestamp 1669390400
transform -1 0 56784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2918__D
timestamp 1669390400
transform -1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2918__RN
timestamp 1669390400
transform 1 0 58016 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2919__CLK
timestamp 1669390400
transform -1 0 51184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2919__D
timestamp 1669390400
transform -1 0 39648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2920__CLK
timestamp 1669390400
transform 1 0 54096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2920__D
timestamp 1669390400
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2921__CLK
timestamp 1669390400
transform -1 0 49392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2921__D
timestamp 1669390400
transform -1 0 45920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2922__CLK
timestamp 1669390400
transform 1 0 54992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2922__D
timestamp 1669390400
transform 1 0 56672 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2923__CLK
timestamp 1669390400
transform -1 0 36960 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2923__D
timestamp 1669390400
transform -1 0 36512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2924__CLK
timestamp 1669390400
transform 1 0 40768 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2924__D
timestamp 1669390400
transform -1 0 41440 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2925__CLK
timestamp 1669390400
transform -1 0 36960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2925__D
timestamp 1669390400
transform 1 0 36288 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2926__CLK
timestamp 1669390400
transform 1 0 37744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2926__D
timestamp 1669390400
transform 1 0 38304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2927__CLK
timestamp 1669390400
transform 1 0 37632 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2927__D
timestamp 1669390400
transform -1 0 38304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2928__CLK
timestamp 1669390400
transform -1 0 48944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2928__D
timestamp 1669390400
transform -1 0 44800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2929__CLK
timestamp 1669390400
transform 1 0 7728 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2929__RN
timestamp 1669390400
transform 1 0 5712 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2930__CLK
timestamp 1669390400
transform -1 0 8288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2930__D
timestamp 1669390400
transform -1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2930__RN
timestamp 1669390400
transform 1 0 9632 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2931__CLK
timestamp 1669390400
transform 1 0 50624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2931__D
timestamp 1669390400
transform -1 0 49056 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2931__RN
timestamp 1669390400
transform 1 0 51184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2933__CLK
timestamp 1669390400
transform 1 0 50288 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2933__D
timestamp 1669390400
transform 1 0 55552 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2933__RN
timestamp 1669390400
transform -1 0 50064 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2934__CLK
timestamp 1669390400
transform 1 0 37520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2935__CLK
timestamp 1669390400
transform 1 0 25536 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2935__D
timestamp 1669390400
transform -1 0 26208 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2937__CLK
timestamp 1669390400
transform 1 0 23184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2937__D
timestamp 1669390400
transform 1 0 28336 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2938__CLK
timestamp 1669390400
transform 1 0 38192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2938__RN
timestamp 1669390400
transform -1 0 33712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__CLK
timestamp 1669390400
transform 1 0 34496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__D
timestamp 1669390400
transform 1 0 40768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__2939__RN
timestamp 1669390400
transform 1 0 35392 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_CLK_I
timestamp 1669390400
transform 1 0 52416 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout42_I
timestamp 1669390400
transform -1 0 40208 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout43_I
timestamp 1669390400
transform -1 0 38864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout44_I
timestamp 1669390400
transform 1 0 30688 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout45_I
timestamp 1669390400
transform 1 0 30240 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout46_I
timestamp 1669390400
transform 1 0 28672 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout47_I
timestamp 1669390400
transform 1 0 53088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout48_I
timestamp 1669390400
transform 1 0 10528 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout49_I
timestamp 1669390400
transform 1 0 22064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout50_I
timestamp 1669390400
transform -1 0 11200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout51_I
timestamp 1669390400
transform 1 0 51408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout52_I
timestamp 1669390400
transform -1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout53_I
timestamp 1669390400
transform -1 0 48160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout54_I
timestamp 1669390400
transform 1 0 56560 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout55_I
timestamp 1669390400
transform -1 0 49840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout56_I
timestamp 1669390400
transform 1 0 38416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout57_I
timestamp 1669390400
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout58_I
timestamp 1669390400
transform 1 0 47488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_fanout59_I
timestamp 1669390400
transform -1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1669390400
transform -1 0 1904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1669390400
transform -1 0 31472 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1669390400
transform -1 0 4704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output8_I
timestamp 1669390400
transform -1 0 4816 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1669390400
transform -1 0 20272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output16_I
timestamp 1669390400
transform 1 0 2912 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1669390400
transform -1 0 36512 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output18_I
timestamp 1669390400
transform -1 0 54320 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output19_I
timestamp 1669390400
transform 1 0 3472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output20_I
timestamp 1669390400
transform 1 0 55440 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output21_I
timestamp 1669390400
transform -1 0 14000 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output24_I
timestamp 1669390400
transform 1 0 54544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output28_I
timestamp 1669390400
transform -1 0 42560 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output29_I
timestamp 1669390400
transform -1 0 56560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output30_I
timestamp 1669390400
transform -1 0 19376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output31_I
timestamp 1669390400
transform -1 0 25424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output32_I
timestamp 1669390400
transform 1 0 55104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output33_I
timestamp 1669390400
transform -1 0 31136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output34_I
timestamp 1669390400
transform 1 0 54320 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output35_I
timestamp 1669390400
transform 1 0 56560 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output36_I
timestamp 1669390400
transform -1 0 21504 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output37_I
timestamp 1669390400
transform -1 0 27664 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output38_I
timestamp 1669390400
transform 1 0 41664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output39_I
timestamp 1669390400
transform -1 0 2464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output40_I
timestamp 1669390400
transform 1 0 3472 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output41_I
timestamp 1669390400
transform 1 0 54880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 4144 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27
timestamp 1669390400
transform 1 0 4368 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30
timestamp 1669390400
transform 1 0 4704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34
timestamp 1669390400
transform 1 0 5152 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1669390400
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54
timestamp 1669390400
transform 1 0 7392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58
timestamp 1669390400
transform 1 0 7840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_62
timestamp 1669390400
transform 1 0 8288 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_72
timestamp 1669390400
transform 1 0 9408 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_76
timestamp 1669390400
transform 1 0 9856 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_80
timestamp 1669390400
transform 1 0 10304 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_84
timestamp 1669390400
transform 1 0 10752 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_88
timestamp 1669390400
transform 1 0 11200 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_104
timestamp 1669390400
transform 1 0 12992 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_107
timestamp 1669390400
transform 1 0 13328 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_110
timestamp 1669390400
transform 1 0 13664 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_116
timestamp 1669390400
transform 1 0 14336 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_120
timestamp 1669390400
transform 1 0 14784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_124
timestamp 1669390400
transform 1 0 15232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_128
timestamp 1669390400
transform 1 0 15680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_130
timestamp 1669390400
transform 1 0 15904 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_133
timestamp 1669390400
transform 1 0 16240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1669390400
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_142
timestamp 1669390400
transform 1 0 17248 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_157
timestamp 1669390400
transform 1 0 18928 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_161
timestamp 1669390400
transform 1 0 19376 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_165
timestamp 1669390400
transform 1 0 19824 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_169
timestamp 1669390400
transform 1 0 20272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_173
timestamp 1669390400
transform 1 0 20720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_177 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 21168 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_207
timestamp 1669390400
transform 1 0 24528 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1669390400
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_212
timestamp 1669390400
transform 1 0 25088 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_215
timestamp 1669390400
transform 1 0 25424 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_231
timestamp 1669390400
transform 1 0 27216 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_239
timestamp 1669390400
transform 1 0 28112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_243
timestamp 1669390400
transform 1 0 28560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1669390400
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_262
timestamp 1669390400
transform 1 0 30688 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_266
timestamp 1669390400
transform 1 0 31136 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_274
timestamp 1669390400
transform 1 0 32032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_278
timestamp 1669390400
transform 1 0 32480 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_282
timestamp 1669390400
transform 1 0 32928 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_290
timestamp 1669390400
transform 1 0 33824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_294
timestamp 1669390400
transform 1 0 34272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_309
timestamp 1669390400
transform 1 0 35952 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_313
timestamp 1669390400
transform 1 0 36400 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_317
timestamp 1669390400
transform 1 0 36848 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_321
timestamp 1669390400
transform 1 0 37296 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_325
timestamp 1669390400
transform 1 0 37744 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_329
timestamp 1669390400
transform 1 0 38192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_333
timestamp 1669390400
transform 1 0 38640 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1669390400
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_352
timestamp 1669390400
transform 1 0 40768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_358
timestamp 1669390400
transform 1 0 41440 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_362
timestamp 1669390400
transform 1 0 41888 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_364
timestamp 1669390400
transform 1 0 42112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_381
timestamp 1669390400
transform 1 0 44016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_387
timestamp 1669390400
transform 1 0 44688 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_394
timestamp 1669390400
transform 1 0 45472 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_398
timestamp 1669390400
transform 1 0 45920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_402
timestamp 1669390400
transform 1 0 46368 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_406
timestamp 1669390400
transform 1 0 46816 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_410
timestamp 1669390400
transform 1 0 47264 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_414
timestamp 1669390400
transform 1 0 47712 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_418
timestamp 1669390400
transform 1 0 48160 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_422
timestamp 1669390400
transform 1 0 48608 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_425
timestamp 1669390400
transform 1 0 48944 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_429
timestamp 1669390400
transform 1 0 49392 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_433
timestamp 1669390400
transform 1 0 49840 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_441
timestamp 1669390400
transform 1 0 50736 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_445
timestamp 1669390400
transform 1 0 51184 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_449
timestamp 1669390400
transform 1 0 51632 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_453
timestamp 1669390400
transform 1 0 52080 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_457
timestamp 1669390400
transform 1 0 52528 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_472
timestamp 1669390400
transform 1 0 54208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_474
timestamp 1669390400
transform 1 0 54432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_489
timestamp 1669390400
transform 1 0 56112 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_492
timestamp 1669390400
transform 1 0 56448 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_495
timestamp 1669390400
transform 1 0 56784 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_499
timestamp 1669390400
transform 1 0 57232 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_503
timestamp 1669390400
transform 1 0 57680 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_507
timestamp 1669390400
transform 1 0 58128 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_2
timestamp 1669390400
transform 1 0 1568 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_6
timestamp 1669390400
transform 1 0 2016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_14
timestamp 1669390400
transform 1 0 2912 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_18
timestamp 1669390400
transform 1 0 3360 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_22
timestamp 1669390400
transform 1 0 3808 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_26
timestamp 1669390400
transform 1 0 4256 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_30
timestamp 1669390400
transform 1 0 4704 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_34
timestamp 1669390400
transform 1 0 5152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_38
timestamp 1669390400
transform 1 0 5600 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_42
timestamp 1669390400
transform 1 0 6048 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_46
timestamp 1669390400
transform 1 0 6496 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_50
timestamp 1669390400
transform 1 0 6944 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_54
timestamp 1669390400
transform 1 0 7392 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_58
timestamp 1669390400
transform 1 0 7840 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_62
timestamp 1669390400
transform 1 0 8288 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_66
timestamp 1669390400
transform 1 0 8736 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_70
timestamp 1669390400
transform 1 0 9184 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_73
timestamp 1669390400
transform 1 0 9520 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_75
timestamp 1669390400
transform 1 0 9744 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_78
timestamp 1669390400
transform 1 0 10080 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_82
timestamp 1669390400
transform 1 0 10528 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_86
timestamp 1669390400
transform 1 0 10976 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_90
timestamp 1669390400
transform 1 0 11424 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_94
timestamp 1669390400
transform 1 0 11872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_96
timestamp 1669390400
transform 1 0 12096 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_99
timestamp 1669390400
transform 1 0 12432 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_103
timestamp 1669390400
transform 1 0 12880 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_106
timestamp 1669390400
transform 1 0 13216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_112
timestamp 1669390400
transform 1 0 13888 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_116
timestamp 1669390400
transform 1 0 14336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_120
timestamp 1669390400
transform 1 0 14784 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_126
timestamp 1669390400
transform 1 0 15456 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_130
timestamp 1669390400
transform 1 0 15904 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_134
timestamp 1669390400
transform 1 0 16352 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_137
timestamp 1669390400
transform 1 0 16688 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1669390400
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_144
timestamp 1669390400
transform 1 0 17472 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_147
timestamp 1669390400
transform 1 0 17808 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_153
timestamp 1669390400
transform 1 0 18480 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_157
timestamp 1669390400
transform 1 0 18928 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_161
timestamp 1669390400
transform 1 0 19376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_165
timestamp 1669390400
transform 1 0 19824 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_168
timestamp 1669390400
transform 1 0 20160 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_172
timestamp 1669390400
transform 1 0 20608 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_176
timestamp 1669390400
transform 1 0 21056 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_180
timestamp 1669390400
transform 1 0 21504 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_184
timestamp 1669390400
transform 1 0 21952 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_186
timestamp 1669390400
transform 1 0 22176 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_189
timestamp 1669390400
transform 1 0 22512 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_205
timestamp 1669390400
transform 1 0 24304 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1669390400
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1669390400
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_286
timestamp 1669390400
transform 1 0 33376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_290
timestamp 1669390400
transform 1 0 33824 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_292
timestamp 1669390400
transform 1 0 34048 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_343
timestamp 1669390400
transform 1 0 39760 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_347
timestamp 1669390400
transform 1 0 40208 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_350
timestamp 1669390400
transform 1 0 40544 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1669390400
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_357
timestamp 1669390400
transform 1 0 41328 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_411
timestamp 1669390400
transform 1 0 47376 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_419
timestamp 1669390400
transform 1 0 48272 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_425
timestamp 1669390400
transform 1 0 48944 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_428
timestamp 1669390400
transform 1 0 49280 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_463
timestamp 1669390400
transform 1 0 53200 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_469
timestamp 1669390400
transform 1 0 53872 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_473
timestamp 1669390400
transform 1 0 54320 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_491
timestamp 1669390400
transform 1 0 56336 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_495
timestamp 1669390400
transform 1 0 56784 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_499
timestamp 1669390400
transform 1 0 57232 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_506
timestamp 1669390400
transform 1 0 58016 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_508
timestamp 1669390400
transform 1 0 58240 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_2
timestamp 1669390400
transform 1 0 1568 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_8
timestamp 1669390400
transform 1 0 2240 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_12
timestamp 1669390400
transform 1 0 2688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_16
timestamp 1669390400
transform 1 0 3136 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_19
timestamp 1669390400
transform 1 0 3472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_23
timestamp 1669390400
transform 1 0 3920 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_27
timestamp 1669390400
transform 1 0 4368 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_30
timestamp 1669390400
transform 1 0 4704 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1669390400
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_37
timestamp 1669390400
transform 1 0 5488 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_39
timestamp 1669390400
transform 1 0 5712 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_42
timestamp 1669390400
transform 1 0 6048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_46
timestamp 1669390400
transform 1 0 6496 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_50
timestamp 1669390400
transform 1 0 6944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_54
timestamp 1669390400
transform 1 0 7392 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_56
timestamp 1669390400
transform 1 0 7616 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_59
timestamp 1669390400
transform 1 0 7952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_63
timestamp 1669390400
transform 1 0 8400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_67
timestamp 1669390400
transform 1 0 8848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_71
timestamp 1669390400
transform 1 0 9296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_75
timestamp 1669390400
transform 1 0 9744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_79
timestamp 1669390400
transform 1 0 10192 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_83
timestamp 1669390400
transform 1 0 10640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_85
timestamp 1669390400
transform 1 0 10864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_88
timestamp 1669390400
transform 1 0 11200 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_92
timestamp 1669390400
transform 1 0 11648 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_96
timestamp 1669390400
transform 1 0 12096 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_99
timestamp 1669390400
transform 1 0 12432 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1669390400
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_108
timestamp 1669390400
transform 1 0 13440 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_114
timestamp 1669390400
transform 1 0 14112 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_118
timestamp 1669390400
transform 1 0 14560 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_121
timestamp 1669390400
transform 1 0 14896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_123
timestamp 1669390400
transform 1 0 15120 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_126
timestamp 1669390400
transform 1 0 15456 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_130
timestamp 1669390400
transform 1 0 15904 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_134
timestamp 1669390400
transform 1 0 16352 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_140
timestamp 1669390400
transform 1 0 17024 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_144
timestamp 1669390400
transform 1 0 17472 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_148
timestamp 1669390400
transform 1 0 17920 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_152
timestamp 1669390400
transform 1 0 18368 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_156
timestamp 1669390400
transform 1 0 18816 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_159
timestamp 1669390400
transform 1 0 19152 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_163
timestamp 1669390400
transform 1 0 19600 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_167
timestamp 1669390400
transform 1 0 20048 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_171
timestamp 1669390400
transform 1 0 20496 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_175
timestamp 1669390400
transform 1 0 20944 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_179
timestamp 1669390400
transform 1 0 21392 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_182
timestamp 1669390400
transform 1 0 21728 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_186
timestamp 1669390400
transform 1 0 22176 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_190
timestamp 1669390400
transform 1 0 22624 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_194
timestamp 1669390400
transform 1 0 23072 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_198
timestamp 1669390400
transform 1 0 23520 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_201
timestamp 1669390400
transform 1 0 23856 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_205
timestamp 1669390400
transform 1 0 24304 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_209
timestamp 1669390400
transform 1 0 24752 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_212
timestamp 1669390400
transform 1 0 25088 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_228
timestamp 1669390400
transform 1 0 26880 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_236
timestamp 1669390400
transform 1 0 27776 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_243
timestamp 1669390400
transform 1 0 28560 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1669390400
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_250 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29344 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_282
timestamp 1669390400
transform 1 0 32928 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_286
timestamp 1669390400
transform 1 0 33376 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_288
timestamp 1669390400
transform 1 0 33600 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_295
timestamp 1669390400
transform 1 0 34384 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_299
timestamp 1669390400
transform 1 0 34832 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_307
timestamp 1669390400
transform 1 0 35728 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_311
timestamp 1669390400
transform 1 0 36176 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_314
timestamp 1669390400
transform 1 0 36512 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1669390400
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_321
timestamp 1669390400
transform 1 0 37296 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_356
timestamp 1669390400
transform 1 0 41216 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_358
timestamp 1669390400
transform 1 0 41440 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_384
timestamp 1669390400
transform 1 0 44352 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_388
timestamp 1669390400
transform 1 0 44800 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_392
timestamp 1669390400
transform 1 0 45248 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_427
timestamp 1669390400
transform 1 0 49168 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_431
timestamp 1669390400
transform 1 0 49616 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_434
timestamp 1669390400
transform 1 0 49952 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_438
timestamp 1669390400
transform 1 0 50400 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_442
timestamp 1669390400
transform 1 0 50848 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_446
timestamp 1669390400
transform 1 0 51296 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_450
timestamp 1669390400
transform 1 0 51744 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_454
timestamp 1669390400
transform 1 0 52192 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_458
timestamp 1669390400
transform 1 0 52640 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_460
timestamp 1669390400
transform 1 0 52864 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_463
timestamp 1669390400
transform 1 0 53200 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_466
timestamp 1669390400
transform 1 0 53536 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_470
timestamp 1669390400
transform 1 0 53984 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_473
timestamp 1669390400
transform 1 0 54320 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_477
timestamp 1669390400
transform 1 0 54768 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_481
timestamp 1669390400
transform 1 0 55216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_485
timestamp 1669390400
transform 1 0 55664 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_492
timestamp 1669390400
transform 1 0 56448 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_496
timestamp 1669390400
transform 1 0 56896 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_500
timestamp 1669390400
transform 1 0 57344 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_2_504
timestamp 1669390400
transform 1 0 57792 0 1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_508
timestamp 1669390400
transform 1 0 58240 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_2
timestamp 1669390400
transform 1 0 1568 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_17
timestamp 1669390400
transform 1 0 3248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_21
timestamp 1669390400
transform 1 0 3696 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_25
timestamp 1669390400
transform 1 0 4144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_29
timestamp 1669390400
transform 1 0 4592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_33
timestamp 1669390400
transform 1 0 5040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_37
timestamp 1669390400
transform 1 0 5488 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_41
timestamp 1669390400
transform 1 0 5936 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_45
timestamp 1669390400
transform 1 0 6384 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_49
timestamp 1669390400
transform 1 0 6832 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_51
timestamp 1669390400
transform 1 0 7056 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_54
timestamp 1669390400
transform 1 0 7392 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_58
timestamp 1669390400
transform 1 0 7840 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_62
timestamp 1669390400
transform 1 0 8288 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_66
timestamp 1669390400
transform 1 0 8736 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1669390400
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_73
timestamp 1669390400
transform 1 0 9520 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_82
timestamp 1669390400
transform 1 0 10528 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_86
timestamp 1669390400
transform 1 0 10976 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_88
timestamp 1669390400
transform 1 0 11200 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_91
timestamp 1669390400
transform 1 0 11536 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_99
timestamp 1669390400
transform 1 0 12432 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_107
timestamp 1669390400
transform 1 0 13328 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_109
timestamp 1669390400
transform 1 0 13552 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_112
timestamp 1669390400
transform 1 0 13888 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_116
timestamp 1669390400
transform 1 0 14336 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_120
timestamp 1669390400
transform 1 0 14784 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_124
timestamp 1669390400
transform 1 0 15232 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_130
timestamp 1669390400
transform 1 0 15904 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_134
timestamp 1669390400
transform 1 0 16352 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_138
timestamp 1669390400
transform 1 0 16800 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1669390400
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_144
timestamp 1669390400
transform 1 0 17472 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_150
timestamp 1669390400
transform 1 0 18144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_154
timestamp 1669390400
transform 1 0 18592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_158
timestamp 1669390400
transform 1 0 19040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_166
timestamp 1669390400
transform 1 0 19936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_170
timestamp 1669390400
transform 1 0 20384 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_173
timestamp 1669390400
transform 1 0 20720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_175
timestamp 1669390400
transform 1 0 20944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_178
timestamp 1669390400
transform 1 0 21280 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_180
timestamp 1669390400
transform 1 0 21504 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_183
timestamp 1669390400
transform 1 0 21840 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_189
timestamp 1669390400
transform 1 0 22512 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_193
timestamp 1669390400
transform 1 0 22960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_195
timestamp 1669390400
transform 1 0 23184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_202
timestamp 1669390400
transform 1 0 23968 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_210
timestamp 1669390400
transform 1 0 24864 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1669390400
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_215
timestamp 1669390400
transform 1 0 25424 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_218
timestamp 1669390400
transform 1 0 25760 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_282
timestamp 1669390400
transform 1 0 32928 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_286
timestamp 1669390400
transform 1 0 33376 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_302
timestamp 1669390400
transform 1 0 35168 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_310
timestamp 1669390400
transform 1 0 36064 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_314
timestamp 1669390400
transform 1 0 36512 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_318
timestamp 1669390400
transform 1 0 36960 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1669390400
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_357
timestamp 1669390400
transform 1 0 41328 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_392
timestamp 1669390400
transform 1 0 45248 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_400
timestamp 1669390400
transform 1 0 46144 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_404
timestamp 1669390400
transform 1 0 46592 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_408
timestamp 1669390400
transform 1 0 47040 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_412
timestamp 1669390400
transform 1 0 47488 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_416
timestamp 1669390400
transform 1 0 47936 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_419
timestamp 1669390400
transform 1 0 48272 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_423
timestamp 1669390400
transform 1 0 48720 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_425
timestamp 1669390400
transform 1 0 48944 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_428
timestamp 1669390400
transform 1 0 49280 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_463
timestamp 1669390400
transform 1 0 53200 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_467
timestamp 1669390400
transform 1 0 53648 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_473
timestamp 1669390400
transform 1 0 54320 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_477
timestamp 1669390400
transform 1 0 54768 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_481
timestamp 1669390400
transform 1 0 55216 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_485
timestamp 1669390400
transform 1 0 55664 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_489
timestamp 1669390400
transform 1 0 56112 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_493
timestamp 1669390400
transform 1 0 56560 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_499
timestamp 1669390400
transform 1 0 57232 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_502
timestamp 1669390400
transform 1 0 57568 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_506
timestamp 1669390400
transform 1 0 58016 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_508
timestamp 1669390400
transform 1 0 58240 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_2
timestamp 1669390400
transform 1 0 1568 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_6
timestamp 1669390400
transform 1 0 2016 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_14
timestamp 1669390400
transform 1 0 2912 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_18
timestamp 1669390400
transform 1 0 3360 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_22
timestamp 1669390400
transform 1 0 3808 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_26
timestamp 1669390400
transform 1 0 4256 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_30
timestamp 1669390400
transform 1 0 4704 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1669390400
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_37
timestamp 1669390400
transform 1 0 5488 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_40
timestamp 1669390400
transform 1 0 5824 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_55
timestamp 1669390400
transform 1 0 7504 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_57
timestamp 1669390400
transform 1 0 7728 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_60
timestamp 1669390400
transform 1 0 8064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_70
timestamp 1669390400
transform 1 0 9184 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_80
timestamp 1669390400
transform 1 0 10304 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_88
timestamp 1669390400
transform 1 0 11200 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_100
timestamp 1669390400
transform 1 0 12544 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_102
timestamp 1669390400
transform 1 0 12768 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1669390400
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_108
timestamp 1669390400
transform 1 0 13440 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_117
timestamp 1669390400
transform 1 0 14448 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_125
timestamp 1669390400
transform 1 0 15344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_127
timestamp 1669390400
transform 1 0 15568 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_130
timestamp 1669390400
transform 1 0 15904 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_132
timestamp 1669390400
transform 1 0 16128 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_151
timestamp 1669390400
transform 1 0 18256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_155
timestamp 1669390400
transform 1 0 18704 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_164
timestamp 1669390400
transform 1 0 19712 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_172
timestamp 1669390400
transform 1 0 20608 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1669390400
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_179
timestamp 1669390400
transform 1 0 21392 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_187
timestamp 1669390400
transform 1 0 22288 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_191
timestamp 1669390400
transform 1 0 22736 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_195
timestamp 1669390400
transform 1 0 23184 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_207
timestamp 1669390400
transform 1 0 24528 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_215
timestamp 1669390400
transform 1 0 25424 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_219
timestamp 1669390400
transform 1 0 25872 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_223
timestamp 1669390400
transform 1 0 26320 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_227
timestamp 1669390400
transform 1 0 26768 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1669390400
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1669390400
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1669390400
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1669390400
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1669390400
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_321
timestamp 1669390400
transform 1 0 37296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_327
timestamp 1669390400
transform 1 0 37968 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_363
timestamp 1669390400
transform 1 0 42000 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_365
timestamp 1669390400
transform 1 0 42224 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_382
timestamp 1669390400
transform 1 0 44128 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_384
timestamp 1669390400
transform 1 0 44352 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_387
timestamp 1669390400
transform 1 0 44688 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1669390400
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_392
timestamp 1669390400
transform 1 0 45248 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_427
timestamp 1669390400
transform 1 0 49168 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_431
timestamp 1669390400
transform 1 0 49616 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_435
timestamp 1669390400
transform 1 0 50064 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_439
timestamp 1669390400
transform 1 0 50512 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_443
timestamp 1669390400
transform 1 0 50960 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_447
timestamp 1669390400
transform 1 0 51408 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_451
timestamp 1669390400
transform 1 0 51856 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_455
timestamp 1669390400
transform 1 0 52304 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_459
timestamp 1669390400
transform 1 0 52752 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_463
timestamp 1669390400
transform 1 0 53200 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_466
timestamp 1669390400
transform 1 0 53536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_472
timestamp 1669390400
transform 1 0 54208 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_476
timestamp 1669390400
transform 1 0 54656 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_480
timestamp 1669390400
transform 1 0 55104 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_484
timestamp 1669390400
transform 1 0 55552 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_488
timestamp 1669390400
transform 1 0 56000 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_492
timestamp 1669390400
transform 1 0 56448 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_496
timestamp 1669390400
transform 1 0 56896 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_500
timestamp 1669390400
transform 1 0 57344 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_504
timestamp 1669390400
transform 1 0 57792 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_508
timestamp 1669390400
transform 1 0 58240 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_2
timestamp 1669390400
transform 1 0 1568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_4
timestamp 1669390400
transform 1 0 1792 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_7
timestamp 1669390400
transform 1 0 2128 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_11
timestamp 1669390400
transform 1 0 2576 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_15
timestamp 1669390400
transform 1 0 3024 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_19
timestamp 1669390400
transform 1 0 3472 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_23
timestamp 1669390400
transform 1 0 3920 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_27
timestamp 1669390400
transform 1 0 4368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_31
timestamp 1669390400
transform 1 0 4816 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_39
timestamp 1669390400
transform 1 0 5712 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_49
timestamp 1669390400
transform 1 0 6832 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_59
timestamp 1669390400
transform 1 0 7952 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_63
timestamp 1669390400
transform 1 0 8400 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_70
timestamp 1669390400
transform 1 0 9184 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_73
timestamp 1669390400
transform 1 0 9520 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_98
timestamp 1669390400
transform 1 0 12320 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_106
timestamp 1669390400
transform 1 0 13216 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_112
timestamp 1669390400
transform 1 0 13888 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_120
timestamp 1669390400
transform 1 0 14784 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_130
timestamp 1669390400
transform 1 0 15904 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_132
timestamp 1669390400
transform 1 0 16128 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1669390400
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_144
timestamp 1669390400
transform 1 0 17472 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_152
timestamp 1669390400
transform 1 0 18368 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_162
timestamp 1669390400
transform 1 0 19488 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_166
timestamp 1669390400
transform 1 0 19936 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_176
timestamp 1669390400
transform 1 0 21056 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_178
timestamp 1669390400
transform 1 0 21280 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_185
timestamp 1669390400
transform 1 0 22064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_199
timestamp 1669390400
transform 1 0 23632 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_203
timestamp 1669390400
transform 1 0 24080 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_205
timestamp 1669390400
transform 1 0 24304 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1669390400
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_215
timestamp 1669390400
transform 1 0 25424 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_218
timestamp 1669390400
transform 1 0 25760 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_226
timestamp 1669390400
transform 1 0 26656 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_230
timestamp 1669390400
transform 1 0 27104 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_262
timestamp 1669390400
transform 1 0 30688 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_278
timestamp 1669390400
transform 1 0 32480 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_282
timestamp 1669390400
transform 1 0 32928 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_286
timestamp 1669390400
transform 1 0 33376 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_318
timestamp 1669390400
transform 1 0 36960 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_328
timestamp 1669390400
transform 1 0 38080 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_332
timestamp 1669390400
transform 1 0 38528 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_338
timestamp 1669390400
transform 1 0 39200 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_342
timestamp 1669390400
transform 1 0 39648 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_346
timestamp 1669390400
transform 1 0 40096 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_350
timestamp 1669390400
transform 1 0 40544 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1669390400
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_357
timestamp 1669390400
transform 1 0 41328 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_408
timestamp 1669390400
transform 1 0 47040 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_412
timestamp 1669390400
transform 1 0 47488 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_416
timestamp 1669390400
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_420
timestamp 1669390400
transform 1 0 48384 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_423
timestamp 1669390400
transform 1 0 48720 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_425
timestamp 1669390400
transform 1 0 48944 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_428
timestamp 1669390400
transform 1 0 49280 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_431
timestamp 1669390400
transform 1 0 49616 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_435
timestamp 1669390400
transform 1 0 50064 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_439
timestamp 1669390400
transform 1 0 50512 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_441
timestamp 1669390400
transform 1 0 50736 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_444
timestamp 1669390400
transform 1 0 51072 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_448
timestamp 1669390400
transform 1 0 51520 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_451
timestamp 1669390400
transform 1 0 51856 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_453
timestamp 1669390400
transform 1 0 52080 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_456
timestamp 1669390400
transform 1 0 52416 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_460
timestamp 1669390400
transform 1 0 52864 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_464
timestamp 1669390400
transform 1 0 53312 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_468
timestamp 1669390400
transform 1 0 53760 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_471
timestamp 1669390400
transform 1 0 54096 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_475
timestamp 1669390400
transform 1 0 54544 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_479
timestamp 1669390400
transform 1 0 54992 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_483
timestamp 1669390400
transform 1 0 55440 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_487
timestamp 1669390400
transform 1 0 55888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_491
timestamp 1669390400
transform 1 0 56336 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_494
timestamp 1669390400
transform 1 0 56672 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_496
timestamp 1669390400
transform 1 0 56896 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_499
timestamp 1669390400
transform 1 0 57232 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_502
timestamp 1669390400
transform 1 0 57568 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_506
timestamp 1669390400
transform 1 0 58016 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_508
timestamp 1669390400
transform 1 0 58240 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_2
timestamp 1669390400
transform 1 0 1568 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_5
timestamp 1669390400
transform 1 0 1904 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_7
timestamp 1669390400
transform 1 0 2128 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_10
timestamp 1669390400
transform 1 0 2464 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_14
timestamp 1669390400
transform 1 0 2912 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_18
timestamp 1669390400
transform 1 0 3360 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_22
timestamp 1669390400
transform 1 0 3808 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_26
timestamp 1669390400
transform 1 0 4256 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_30
timestamp 1669390400
transform 1 0 4704 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1669390400
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_37
timestamp 1669390400
transform 1 0 5488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_51
timestamp 1669390400
transform 1 0 7056 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_59
timestamp 1669390400
transform 1 0 7952 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_61
timestamp 1669390400
transform 1 0 8176 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_98
timestamp 1669390400
transform 1 0 12320 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_100
timestamp 1669390400
transform 1 0 12544 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_103
timestamp 1669390400
transform 1 0 12880 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1669390400
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_108
timestamp 1669390400
transform 1 0 13440 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_115
timestamp 1669390400
transform 1 0 14224 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_117
timestamp 1669390400
transform 1 0 14448 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_124
timestamp 1669390400
transform 1 0 15232 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_130
timestamp 1669390400
transform 1 0 15904 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_134
timestamp 1669390400
transform 1 0 16352 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_138
timestamp 1669390400
transform 1 0 16800 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_155
timestamp 1669390400
transform 1 0 18704 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_157
timestamp 1669390400
transform 1 0 18928 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_164
timestamp 1669390400
transform 1 0 19712 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_174
timestamp 1669390400
transform 1 0 20832 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1669390400
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_179
timestamp 1669390400
transform 1 0 21392 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_183
timestamp 1669390400
transform 1 0 21840 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_191
timestamp 1669390400
transform 1 0 22736 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_199
timestamp 1669390400
transform 1 0 23632 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_203
timestamp 1669390400
transform 1 0 24080 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_207
timestamp 1669390400
transform 1 0 24528 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_210
timestamp 1669390400
transform 1 0 24864 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_218
timestamp 1669390400
transform 1 0 25760 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_222
timestamp 1669390400
transform 1 0 26208 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_229
timestamp 1669390400
transform 1 0 26992 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_233
timestamp 1669390400
transform 1 0 27440 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_6_237
timestamp 1669390400
transform 1 0 27888 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_245
timestamp 1669390400
transform 1 0 28784 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1669390400
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1669390400
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1669390400
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1669390400
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_321
timestamp 1669390400
transform 1 0 37296 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_323
timestamp 1669390400
transform 1 0 37520 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_326
timestamp 1669390400
transform 1 0 37856 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_362
timestamp 1669390400
transform 1 0 41888 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_366
timestamp 1669390400
transform 1 0 42336 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_368
timestamp 1669390400
transform 1 0 42560 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_371
timestamp 1669390400
transform 1 0 42896 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_375
timestamp 1669390400
transform 1 0 43344 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_379
timestamp 1669390400
transform 1 0 43792 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_383
timestamp 1669390400
transform 1 0 44240 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1669390400
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_392
timestamp 1669390400
transform 1 0 45248 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_427
timestamp 1669390400
transform 1 0 49168 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_431
timestamp 1669390400
transform 1 0 49616 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_435
timestamp 1669390400
transform 1 0 50064 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_439
timestamp 1669390400
transform 1 0 50512 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_443
timestamp 1669390400
transform 1 0 50960 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_447
timestamp 1669390400
transform 1 0 51408 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_451
timestamp 1669390400
transform 1 0 51856 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_455
timestamp 1669390400
transform 1 0 52304 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_459
timestamp 1669390400
transform 1 0 52752 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_463
timestamp 1669390400
transform 1 0 53200 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_466
timestamp 1669390400
transform 1 0 53536 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_470
timestamp 1669390400
transform 1 0 53984 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_474
timestamp 1669390400
transform 1 0 54432 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_476
timestamp 1669390400
transform 1 0 54656 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_491
timestamp 1669390400
transform 1 0 56336 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_495
timestamp 1669390400
transform 1 0 56784 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_499
timestamp 1669390400
transform 1 0 57232 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_501
timestamp 1669390400
transform 1 0 57456 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_504
timestamp 1669390400
transform 1 0 57792 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_508
timestamp 1669390400
transform 1 0 58240 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_2
timestamp 1669390400
transform 1 0 1568 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_6
timestamp 1669390400
transform 1 0 2016 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_10
timestamp 1669390400
transform 1 0 2464 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_14
timestamp 1669390400
transform 1 0 2912 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_18
timestamp 1669390400
transform 1 0 3360 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_22
timestamp 1669390400
transform 1 0 3808 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_26
timestamp 1669390400
transform 1 0 4256 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_30
timestamp 1669390400
transform 1 0 4704 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_34
timestamp 1669390400
transform 1 0 5152 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_38
timestamp 1669390400
transform 1 0 5600 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_49
timestamp 1669390400
transform 1 0 6832 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_51
timestamp 1669390400
transform 1 0 7056 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_54
timestamp 1669390400
transform 1 0 7392 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_58
timestamp 1669390400
transform 1 0 7840 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_62
timestamp 1669390400
transform 1 0 8288 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_66
timestamp 1669390400
transform 1 0 8736 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_70
timestamp 1669390400
transform 1 0 9184 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_73
timestamp 1669390400
transform 1 0 9520 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_76
timestamp 1669390400
transform 1 0 9856 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_78
timestamp 1669390400
transform 1 0 10080 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_87
timestamp 1669390400
transform 1 0 11088 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_91
timestamp 1669390400
transform 1 0 11536 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_94
timestamp 1669390400
transform 1 0 11872 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_102
timestamp 1669390400
transform 1 0 12768 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_104
timestamp 1669390400
transform 1 0 12992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_107
timestamp 1669390400
transform 1 0 13328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_115
timestamp 1669390400
transform 1 0 14224 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_117
timestamp 1669390400
transform 1 0 14448 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_126
timestamp 1669390400
transform 1 0 15456 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_133
timestamp 1669390400
transform 1 0 16240 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_137
timestamp 1669390400
transform 1 0 16688 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1669390400
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_144
timestamp 1669390400
transform 1 0 17472 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_160
timestamp 1669390400
transform 1 0 19264 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_168
timestamp 1669390400
transform 1 0 20160 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_172
timestamp 1669390400
transform 1 0 20608 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_175
timestamp 1669390400
transform 1 0 20944 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_179
timestamp 1669390400
transform 1 0 21392 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_187
timestamp 1669390400
transform 1 0 22288 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_191
timestamp 1669390400
transform 1 0 22736 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_195
timestamp 1669390400
transform 1 0 23184 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_199
timestamp 1669390400
transform 1 0 23632 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_201
timestamp 1669390400
transform 1 0 23856 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_204
timestamp 1669390400
transform 1 0 24192 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_206
timestamp 1669390400
transform 1 0 24416 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_209
timestamp 1669390400
transform 1 0 24752 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_215
timestamp 1669390400
transform 1 0 25424 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_225
timestamp 1669390400
transform 1 0 26544 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_235
timestamp 1669390400
transform 1 0 27664 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_239
timestamp 1669390400
transform 1 0 28112 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_243
timestamp 1669390400
transform 1 0 28560 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_275
timestamp 1669390400
transform 1 0 32144 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1669390400
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_286
timestamp 1669390400
transform 1 0 33376 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_302
timestamp 1669390400
transform 1 0 35168 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_310
timestamp 1669390400
transform 1 0 36064 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_314
timestamp 1669390400
transform 1 0 36512 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_318
timestamp 1669390400
transform 1 0 36960 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1669390400
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_357
timestamp 1669390400
transform 1 0 41328 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_395
timestamp 1669390400
transform 1 0 45584 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_397
timestamp 1669390400
transform 1 0 45808 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_400
timestamp 1669390400
transform 1 0 46144 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_404
timestamp 1669390400
transform 1 0 46592 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_408
timestamp 1669390400
transform 1 0 47040 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_412
timestamp 1669390400
transform 1 0 47488 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_416
timestamp 1669390400
transform 1 0 47936 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_420
timestamp 1669390400
transform 1 0 48384 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_424
timestamp 1669390400
transform 1 0 48832 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_428
timestamp 1669390400
transform 1 0 49280 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_431
timestamp 1669390400
transform 1 0 49616 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_433
timestamp 1669390400
transform 1 0 49840 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_436
timestamp 1669390400
transform 1 0 50176 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_440
timestamp 1669390400
transform 1 0 50624 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_442
timestamp 1669390400
transform 1 0 50848 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_445
timestamp 1669390400
transform 1 0 51184 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_449
timestamp 1669390400
transform 1 0 51632 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_453
timestamp 1669390400
transform 1 0 52080 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_457
timestamp 1669390400
transform 1 0 52528 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_461
timestamp 1669390400
transform 1 0 52976 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_465
timestamp 1669390400
transform 1 0 53424 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_469
timestamp 1669390400
transform 1 0 53872 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_471
timestamp 1669390400
transform 1 0 54096 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_474
timestamp 1669390400
transform 1 0 54432 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_478
timestamp 1669390400
transform 1 0 54880 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_482
timestamp 1669390400
transform 1 0 55328 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_486
timestamp 1669390400
transform 1 0 55776 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_490
timestamp 1669390400
transform 1 0 56224 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_496
timestamp 1669390400
transform 1 0 56896 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_499
timestamp 1669390400
transform 1 0 57232 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_506
timestamp 1669390400
transform 1 0 58016 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_508
timestamp 1669390400
transform 1 0 58240 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_2
timestamp 1669390400
transform 1 0 1568 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_6
timestamp 1669390400
transform 1 0 2016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_10
timestamp 1669390400
transform 1 0 2464 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_14
timestamp 1669390400
transform 1 0 2912 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_18
timestamp 1669390400
transform 1 0 3360 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_22
timestamp 1669390400
transform 1 0 3808 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_26
timestamp 1669390400
transform 1 0 4256 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1669390400
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_37
timestamp 1669390400
transform 1 0 5488 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_49
timestamp 1669390400
transform 1 0 6832 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_56
timestamp 1669390400
transform 1 0 7616 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_58
timestamp 1669390400
transform 1 0 7840 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_61
timestamp 1669390400
transform 1 0 8176 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_81
timestamp 1669390400
transform 1 0 10416 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_91
timestamp 1669390400
transform 1 0 11536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_97
timestamp 1669390400
transform 1 0 12208 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1669390400
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_108
timestamp 1669390400
transform 1 0 13440 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_117
timestamp 1669390400
transform 1 0 14448 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_119
timestamp 1669390400
transform 1 0 14672 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_138
timestamp 1669390400
transform 1 0 16800 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_140
timestamp 1669390400
transform 1 0 17024 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_151
timestamp 1669390400
transform 1 0 18256 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_159
timestamp 1669390400
transform 1 0 19152 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_163
timestamp 1669390400
transform 1 0 19600 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_166
timestamp 1669390400
transform 1 0 19936 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1669390400
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_179
timestamp 1669390400
transform 1 0 21392 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_197
timestamp 1669390400
transform 1 0 23408 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_205
timestamp 1669390400
transform 1 0 24304 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_209
timestamp 1669390400
transform 1 0 24752 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_213
timestamp 1669390400
transform 1 0 25200 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_226
timestamp 1669390400
transform 1 0 26656 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_234
timestamp 1669390400
transform 1 0 27552 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_238
timestamp 1669390400
transform 1 0 28000 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_242
timestamp 1669390400
transform 1 0 28448 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_246
timestamp 1669390400
transform 1 0 28896 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_250
timestamp 1669390400
transform 1 0 29344 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_253
timestamp 1669390400
transform 1 0 29680 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_317
timestamp 1669390400
transform 1 0 36848 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_321
timestamp 1669390400
transform 1 0 37296 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_325
timestamp 1669390400
transform 1 0 37744 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_361
timestamp 1669390400
transform 1 0 41776 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_369
timestamp 1669390400
transform 1 0 42672 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_373
timestamp 1669390400
transform 1 0 43120 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_377
timestamp 1669390400
transform 1 0 43568 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_381
timestamp 1669390400
transform 1 0 44016 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_385
timestamp 1669390400
transform 1 0 44464 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1669390400
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_392
timestamp 1669390400
transform 1 0 45248 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_427
timestamp 1669390400
transform 1 0 49168 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_454
timestamp 1669390400
transform 1 0 52192 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_458
timestamp 1669390400
transform 1 0 52640 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_460
timestamp 1669390400
transform 1 0 52864 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_463
timestamp 1669390400
transform 1 0 53200 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_466
timestamp 1669390400
transform 1 0 53536 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_470
timestamp 1669390400
transform 1 0 53984 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_474
timestamp 1669390400
transform 1 0 54432 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_478
timestamp 1669390400
transform 1 0 54880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_482
timestamp 1669390400
transform 1 0 55328 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_486
timestamp 1669390400
transform 1 0 55776 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_492
timestamp 1669390400
transform 1 0 56448 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_496
timestamp 1669390400
transform 1 0 56896 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_500
timestamp 1669390400
transform 1 0 57344 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_504
timestamp 1669390400
transform 1 0 57792 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_508
timestamp 1669390400
transform 1 0 58240 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_2
timestamp 1669390400
transform 1 0 1568 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_10
timestamp 1669390400
transform 1 0 2464 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_18
timestamp 1669390400
transform 1 0 3360 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_20
timestamp 1669390400
transform 1 0 3584 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_23
timestamp 1669390400
transform 1 0 3920 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_27
timestamp 1669390400
transform 1 0 4368 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_31
timestamp 1669390400
transform 1 0 4816 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_39
timestamp 1669390400
transform 1 0 5712 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_41
timestamp 1669390400
transform 1 0 5936 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_51
timestamp 1669390400
transform 1 0 7056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_68
timestamp 1669390400
transform 1 0 8960 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_70
timestamp 1669390400
transform 1 0 9184 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_73
timestamp 1669390400
transform 1 0 9520 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_92
timestamp 1669390400
transform 1 0 11648 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_100
timestamp 1669390400
transform 1 0 12544 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_104
timestamp 1669390400
transform 1 0 12992 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_114
timestamp 1669390400
transform 1 0 14112 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_122
timestamp 1669390400
transform 1 0 15008 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_126
timestamp 1669390400
transform 1 0 15456 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1669390400
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_144
timestamp 1669390400
transform 1 0 17472 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_146
timestamp 1669390400
transform 1 0 17696 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_153
timestamp 1669390400
transform 1 0 18480 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_161
timestamp 1669390400
transform 1 0 19376 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_176
timestamp 1669390400
transform 1 0 21056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_182
timestamp 1669390400
transform 1 0 21728 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_197
timestamp 1669390400
transform 1 0 23408 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_207
timestamp 1669390400
transform 1 0 24528 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_211
timestamp 1669390400
transform 1 0 24976 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_215
timestamp 1669390400
transform 1 0 25424 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_223
timestamp 1669390400
transform 1 0 26320 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_227
timestamp 1669390400
transform 1 0 26768 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_236
timestamp 1669390400
transform 1 0 27776 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_244
timestamp 1669390400
transform 1 0 28672 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_248
timestamp 1669390400
transform 1 0 29120 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_251
timestamp 1669390400
transform 1 0 29456 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_255
timestamp 1669390400
transform 1 0 29904 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_259
timestamp 1669390400
transform 1 0 30352 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_275
timestamp 1669390400
transform 1 0 32144 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1669390400
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_286
timestamp 1669390400
transform 1 0 33376 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_294
timestamp 1669390400
transform 1 0 34272 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_302
timestamp 1669390400
transform 1 0 35168 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_312
timestamp 1669390400
transform 1 0 36288 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_322
timestamp 1669390400
transform 1 0 37408 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_326
timestamp 1669390400
transform 1 0 37856 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_330
timestamp 1669390400
transform 1 0 38304 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_334
timestamp 1669390400
transform 1 0 38752 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_338
timestamp 1669390400
transform 1 0 39200 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_342
timestamp 1669390400
transform 1 0 39648 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_344
timestamp 1669390400
transform 1 0 39872 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_347
timestamp 1669390400
transform 1 0 40208 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_351
timestamp 1669390400
transform 1 0 40656 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_357
timestamp 1669390400
transform 1 0 41328 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_360
timestamp 1669390400
transform 1 0 41664 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_364
timestamp 1669390400
transform 1 0 42112 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_370
timestamp 1669390400
transform 1 0 42784 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_374
timestamp 1669390400
transform 1 0 43232 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_378
timestamp 1669390400
transform 1 0 43680 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_382
timestamp 1669390400
transform 1 0 44128 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_386
timestamp 1669390400
transform 1 0 44576 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_422
timestamp 1669390400
transform 1 0 48608 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_428
timestamp 1669390400
transform 1 0 49280 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_431
timestamp 1669390400
transform 1 0 49616 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_435
timestamp 1669390400
transform 1 0 50064 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_439
timestamp 1669390400
transform 1 0 50512 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_443
timestamp 1669390400
transform 1 0 50960 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_447
timestamp 1669390400
transform 1 0 51408 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_451
timestamp 1669390400
transform 1 0 51856 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_455
timestamp 1669390400
transform 1 0 52304 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_459
timestamp 1669390400
transform 1 0 52752 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_463
timestamp 1669390400
transform 1 0 53200 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_467
timestamp 1669390400
transform 1 0 53648 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_471
timestamp 1669390400
transform 1 0 54096 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_475
timestamp 1669390400
transform 1 0 54544 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_479
timestamp 1669390400
transform 1 0 54992 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_483
timestamp 1669390400
transform 1 0 55440 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_487
timestamp 1669390400
transform 1 0 55888 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_491
timestamp 1669390400
transform 1 0 56336 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_494
timestamp 1669390400
transform 1 0 56672 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_496
timestamp 1669390400
transform 1 0 56896 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_499
timestamp 1669390400
transform 1 0 57232 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_502
timestamp 1669390400
transform 1 0 57568 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_506
timestamp 1669390400
transform 1 0 58016 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_508
timestamp 1669390400
transform 1 0 58240 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_2
timestamp 1669390400
transform 1 0 1568 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_5
timestamp 1669390400
transform 1 0 1904 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_13
timestamp 1669390400
transform 1 0 2800 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_21
timestamp 1669390400
transform 1 0 3696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_25
timestamp 1669390400
transform 1 0 4144 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1669390400
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_37
timestamp 1669390400
transform 1 0 5488 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_41
timestamp 1669390400
transform 1 0 5936 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_86
timestamp 1669390400
transform 1 0 10976 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_95
timestamp 1669390400
transform 1 0 11984 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_103
timestamp 1669390400
transform 1 0 12880 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1669390400
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_108
timestamp 1669390400
transform 1 0 13440 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_124
timestamp 1669390400
transform 1 0 15232 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_128
timestamp 1669390400
transform 1 0 15680 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_131
timestamp 1669390400
transform 1 0 16016 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1669390400
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_179
timestamp 1669390400
transform 1 0 21392 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_182
timestamp 1669390400
transform 1 0 21728 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_184
timestamp 1669390400
transform 1 0 21952 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_187
timestamp 1669390400
transform 1 0 22288 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_197
timestamp 1669390400
transform 1 0 23408 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_205
timestamp 1669390400
transform 1 0 24304 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_213
timestamp 1669390400
transform 1 0 25200 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_224
timestamp 1669390400
transform 1 0 26432 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_226
timestamp 1669390400
transform 1 0 26656 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_235
timestamp 1669390400
transform 1 0 27664 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1669390400
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_250
timestamp 1669390400
transform 1 0 29344 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_257
timestamp 1669390400
transform 1 0 30128 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_261
timestamp 1669390400
transform 1 0 30576 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_265
timestamp 1669390400
transform 1 0 31024 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_281
timestamp 1669390400
transform 1 0 32816 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_295
timestamp 1669390400
transform 1 0 34384 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_299
timestamp 1669390400
transform 1 0 34832 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_305
timestamp 1669390400
transform 1 0 35504 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_309
timestamp 1669390400
transform 1 0 35952 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_311
timestamp 1669390400
transform 1 0 36176 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_314
timestamp 1669390400
transform 1 0 36512 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1669390400
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_321
timestamp 1669390400
transform 1 0 37296 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_323
timestamp 1669390400
transform 1 0 37520 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_326
timestamp 1669390400
transform 1 0 37856 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_362
timestamp 1669390400
transform 1 0 41888 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_366
timestamp 1669390400
transform 1 0 42336 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_370
timestamp 1669390400
transform 1 0 42784 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_374
timestamp 1669390400
transform 1 0 43232 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_378
timestamp 1669390400
transform 1 0 43680 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_382
timestamp 1669390400
transform 1 0 44128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_386
timestamp 1669390400
transform 1 0 44576 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1669390400
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_392
timestamp 1669390400
transform 1 0 45248 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_396
timestamp 1669390400
transform 1 0 45696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_402
timestamp 1669390400
transform 1 0 46368 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_406
timestamp 1669390400
transform 1 0 46816 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_410
timestamp 1669390400
transform 1 0 47264 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_414
timestamp 1669390400
transform 1 0 47712 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_418
timestamp 1669390400
transform 1 0 48160 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_426
timestamp 1669390400
transform 1 0 49056 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_430
timestamp 1669390400
transform 1 0 49504 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_434
timestamp 1669390400
transform 1 0 49952 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_438
timestamp 1669390400
transform 1 0 50400 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_442
timestamp 1669390400
transform 1 0 50848 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_444
timestamp 1669390400
transform 1 0 51072 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_451
timestamp 1669390400
transform 1 0 51856 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_455
timestamp 1669390400
transform 1 0 52304 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_457
timestamp 1669390400
transform 1 0 52528 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_460
timestamp 1669390400
transform 1 0 52864 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_463
timestamp 1669390400
transform 1 0 53200 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_466
timestamp 1669390400
transform 1 0 53536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_476
timestamp 1669390400
transform 1 0 54656 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_480
timestamp 1669390400
transform 1 0 55104 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_484
timestamp 1669390400
transform 1 0 55552 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_488
timestamp 1669390400
transform 1 0 56000 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_492
timestamp 1669390400
transform 1 0 56448 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_496
timestamp 1669390400
transform 1 0 56896 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_500
timestamp 1669390400
transform 1 0 57344 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_10_504
timestamp 1669390400
transform 1 0 57792 0 1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_508
timestamp 1669390400
transform 1 0 58240 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_2
timestamp 1669390400
transform 1 0 1568 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_17
timestamp 1669390400
transform 1 0 3248 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_21
timestamp 1669390400
transform 1 0 3696 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_29
timestamp 1669390400
transform 1 0 4592 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_47
timestamp 1669390400
transform 1 0 6608 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_62
timestamp 1669390400
transform 1 0 8288 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1669390400
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_73
timestamp 1669390400
transform 1 0 9520 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_90
timestamp 1669390400
transform 1 0 11424 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_94
timestamp 1669390400
transform 1 0 11872 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_102
timestamp 1669390400
transform 1 0 12768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_110
timestamp 1669390400
transform 1 0 13664 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_118
timestamp 1669390400
transform 1 0 14560 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_122
timestamp 1669390400
transform 1 0 15008 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_125
timestamp 1669390400
transform 1 0 15344 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_129
timestamp 1669390400
transform 1 0 15792 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_133
timestamp 1669390400
transform 1 0 16240 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1669390400
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_144
timestamp 1669390400
transform 1 0 17472 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_150
timestamp 1669390400
transform 1 0 18144 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_159
timestamp 1669390400
transform 1 0 19152 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_169
timestamp 1669390400
transform 1 0 20272 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_177
timestamp 1669390400
transform 1 0 21168 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_181
timestamp 1669390400
transform 1 0 21616 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_188
timestamp 1669390400
transform 1 0 22400 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_190
timestamp 1669390400
transform 1 0 22624 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_197
timestamp 1669390400
transform 1 0 23408 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_201
timestamp 1669390400
transform 1 0 23856 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_209
timestamp 1669390400
transform 1 0 24752 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_215
timestamp 1669390400
transform 1 0 25424 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_218
timestamp 1669390400
transform 1 0 25760 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_222
timestamp 1669390400
transform 1 0 26208 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_226
timestamp 1669390400
transform 1 0 26656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_230
timestamp 1669390400
transform 1 0 27104 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_237
timestamp 1669390400
transform 1 0 27888 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_241
timestamp 1669390400
transform 1 0 28336 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_248
timestamp 1669390400
transform 1 0 29120 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_256
timestamp 1669390400
transform 1 0 30016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_260
timestamp 1669390400
transform 1 0 30464 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_264
timestamp 1669390400
transform 1 0 30912 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_268
timestamp 1669390400
transform 1 0 31360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_276
timestamp 1669390400
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_280
timestamp 1669390400
transform 1 0 32704 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1669390400
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_286
timestamp 1669390400
transform 1 0 33376 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_303
timestamp 1669390400
transform 1 0 35280 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_320
timestamp 1669390400
transform 1 0 37184 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_324
timestamp 1669390400
transform 1 0 37632 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_328
timestamp 1669390400
transform 1 0 38080 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_331
timestamp 1669390400
transform 1 0 38416 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_335
timestamp 1669390400
transform 1 0 38864 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_339
timestamp 1669390400
transform 1 0 39312 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_343
timestamp 1669390400
transform 1 0 39760 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_346
timestamp 1669390400
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_352
timestamp 1669390400
transform 1 0 40768 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1669390400
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_357
timestamp 1669390400
transform 1 0 41328 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_360
timestamp 1669390400
transform 1 0 41664 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_364
timestamp 1669390400
transform 1 0 42112 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_367
timestamp 1669390400
transform 1 0 42448 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_371
timestamp 1669390400
transform 1 0 42896 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_373
timestamp 1669390400
transform 1 0 43120 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_376
timestamp 1669390400
transform 1 0 43456 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_380
timestamp 1669390400
transform 1 0 43904 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_390
timestamp 1669390400
transform 1 0 45024 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_398
timestamp 1669390400
transform 1 0 45920 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_402
timestamp 1669390400
transform 1 0 46368 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_406
timestamp 1669390400
transform 1 0 46816 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_412
timestamp 1669390400
transform 1 0 47488 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_416
timestamp 1669390400
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_420
timestamp 1669390400
transform 1 0 48384 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_425
timestamp 1669390400
transform 1 0 48944 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_428
timestamp 1669390400
transform 1 0 49280 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_435
timestamp 1669390400
transform 1 0 50064 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_439
timestamp 1669390400
transform 1 0 50512 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_443
timestamp 1669390400
transform 1 0 50960 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_447
timestamp 1669390400
transform 1 0 51408 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_451
timestamp 1669390400
transform 1 0 51856 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_459
timestamp 1669390400
transform 1 0 52752 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_467
timestamp 1669390400
transform 1 0 53648 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_482
timestamp 1669390400
transform 1 0 55328 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_490
timestamp 1669390400
transform 1 0 56224 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_494
timestamp 1669390400
transform 1 0 56672 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_496
timestamp 1669390400
transform 1 0 56896 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_499
timestamp 1669390400
transform 1 0 57232 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_502
timestamp 1669390400
transform 1 0 57568 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_506
timestamp 1669390400
transform 1 0 58016 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_508
timestamp 1669390400
transform 1 0 58240 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_2
timestamp 1669390400
transform 1 0 1568 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_6
timestamp 1669390400
transform 1 0 2016 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_14
timestamp 1669390400
transform 1 0 2912 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_18
timestamp 1669390400
transform 1 0 3360 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_25
timestamp 1669390400
transform 1 0 4144 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_27
timestamp 1669390400
transform 1 0 4368 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_30
timestamp 1669390400
transform 1 0 4704 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1669390400
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_37
timestamp 1669390400
transform 1 0 5488 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_39
timestamp 1669390400
transform 1 0 5712 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_73
timestamp 1669390400
transform 1 0 9520 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_79
timestamp 1669390400
transform 1 0 10192 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1669390400
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_108
timestamp 1669390400
transform 1 0 13440 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_112
timestamp 1669390400
transform 1 0 13888 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_120
timestamp 1669390400
transform 1 0 14784 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_124
timestamp 1669390400
transform 1 0 15232 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_128
timestamp 1669390400
transform 1 0 15680 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_132
timestamp 1669390400
transform 1 0 16128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_142
timestamp 1669390400
transform 1 0 17248 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_150
timestamp 1669390400
transform 1 0 18144 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_161
timestamp 1669390400
transform 1 0 19376 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1669390400
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_179
timestamp 1669390400
transform 1 0 21392 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_182
timestamp 1669390400
transform 1 0 21728 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_190
timestamp 1669390400
transform 1 0 22624 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_192
timestamp 1669390400
transform 1 0 22848 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_195
timestamp 1669390400
transform 1 0 23184 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_197
timestamp 1669390400
transform 1 0 23408 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_204
timestamp 1669390400
transform 1 0 24192 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_210
timestamp 1669390400
transform 1 0 24864 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_218
timestamp 1669390400
transform 1 0 25760 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_228
timestamp 1669390400
transform 1 0 26880 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_234
timestamp 1669390400
transform 1 0 27552 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_238
timestamp 1669390400
transform 1 0 28000 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_244
timestamp 1669390400
transform 1 0 28672 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_250
timestamp 1669390400
transform 1 0 29344 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_253
timestamp 1669390400
transform 1 0 29680 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_257
timestamp 1669390400
transform 1 0 30128 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_261
timestamp 1669390400
transform 1 0 30576 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_265
timestamp 1669390400
transform 1 0 31024 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_12_269
timestamp 1669390400
transform 1 0 31472 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_277
timestamp 1669390400
transform 1 0 32368 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_283
timestamp 1669390400
transform 1 0 33040 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_293
timestamp 1669390400
transform 1 0 34160 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_300
timestamp 1669390400
transform 1 0 34944 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_304
timestamp 1669390400
transform 1 0 35392 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_308
timestamp 1669390400
transform 1 0 35840 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_314
timestamp 1669390400
transform 1 0 36512 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1669390400
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_321
timestamp 1669390400
transform 1 0 37296 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_329
timestamp 1669390400
transform 1 0 38192 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_331
timestamp 1669390400
transform 1 0 38416 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_334
timestamp 1669390400
transform 1 0 38752 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_342
timestamp 1669390400
transform 1 0 39648 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_349
timestamp 1669390400
transform 1 0 40432 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_356
timestamp 1669390400
transform 1 0 41216 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_370
timestamp 1669390400
transform 1 0 42784 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_372
timestamp 1669390400
transform 1 0 43008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_379
timestamp 1669390400
transform 1 0 43792 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_383
timestamp 1669390400
transform 1 0 44240 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_387
timestamp 1669390400
transform 1 0 44688 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1669390400
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_392
timestamp 1669390400
transform 1 0 45248 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_405
timestamp 1669390400
transform 1 0 46704 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_407
timestamp 1669390400
transform 1 0 46928 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_410
timestamp 1669390400
transform 1 0 47264 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_412
timestamp 1669390400
transform 1 0 47488 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_421
timestamp 1669390400
transform 1 0 48496 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_423
timestamp 1669390400
transform 1 0 48720 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_434
timestamp 1669390400
transform 1 0 49952 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_442
timestamp 1669390400
transform 1 0 50848 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_452
timestamp 1669390400
transform 1 0 51968 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_460
timestamp 1669390400
transform 1 0 52864 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_463
timestamp 1669390400
transform 1 0 53200 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_466
timestamp 1669390400
transform 1 0 53536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_476
timestamp 1669390400
transform 1 0 54656 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_483
timestamp 1669390400
transform 1 0 55440 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_487
timestamp 1669390400
transform 1 0 55888 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_491
timestamp 1669390400
transform 1 0 56336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_495
timestamp 1669390400
transform 1 0 56784 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_502
timestamp 1669390400
transform 1 0 57568 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_506
timestamp 1669390400
transform 1 0 58016 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_508
timestamp 1669390400
transform 1 0 58240 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_2
timestamp 1669390400
transform 1 0 1568 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_5
timestamp 1669390400
transform 1 0 1904 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_9
timestamp 1669390400
transform 1 0 2352 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_13
timestamp 1669390400
transform 1 0 2800 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_17
timestamp 1669390400
transform 1 0 3248 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_21
timestamp 1669390400
transform 1 0 3696 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_25
timestamp 1669390400
transform 1 0 4144 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_29
timestamp 1669390400
transform 1 0 4592 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_33
timestamp 1669390400
transform 1 0 5040 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_37
timestamp 1669390400
transform 1 0 5488 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_45
timestamp 1669390400
transform 1 0 6384 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_47
timestamp 1669390400
transform 1 0 6608 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_50
timestamp 1669390400
transform 1 0 6944 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_54
timestamp 1669390400
transform 1 0 7392 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_61
timestamp 1669390400
transform 1 0 8176 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_69
timestamp 1669390400
transform 1 0 9072 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_73
timestamp 1669390400
transform 1 0 9520 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_117
timestamp 1669390400
transform 1 0 14448 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_121
timestamp 1669390400
transform 1 0 14896 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_131
timestamp 1669390400
transform 1 0 16016 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1669390400
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_144
timestamp 1669390400
transform 1 0 17472 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_148
timestamp 1669390400
transform 1 0 17920 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_152
timestamp 1669390400
transform 1 0 18368 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_156
timestamp 1669390400
transform 1 0 18816 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_160
timestamp 1669390400
transform 1 0 19264 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_164
timestamp 1669390400
transform 1 0 19712 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_168
timestamp 1669390400
transform 1 0 20160 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_171
timestamp 1669390400
transform 1 0 20496 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_187
timestamp 1669390400
transform 1 0 22288 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_191
timestamp 1669390400
transform 1 0 22736 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_193
timestamp 1669390400
transform 1 0 22960 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_207
timestamp 1669390400
transform 1 0 24528 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_211
timestamp 1669390400
transform 1 0 24976 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_215
timestamp 1669390400
transform 1 0 25424 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_217
timestamp 1669390400
transform 1 0 25648 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_236
timestamp 1669390400
transform 1 0 27776 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_248
timestamp 1669390400
transform 1 0 29120 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_262
timestamp 1669390400
transform 1 0 30688 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_266
timestamp 1669390400
transform 1 0 31136 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_270
timestamp 1669390400
transform 1 0 31584 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_278
timestamp 1669390400
transform 1 0 32480 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_282
timestamp 1669390400
transform 1 0 32928 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_286
timestamp 1669390400
transform 1 0 33376 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_293
timestamp 1669390400
transform 1 0 34160 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_297
timestamp 1669390400
transform 1 0 34608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_301
timestamp 1669390400
transform 1 0 35056 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_304
timestamp 1669390400
transform 1 0 35392 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_308
timestamp 1669390400
transform 1 0 35840 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_322
timestamp 1669390400
transform 1 0 37408 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_326
timestamp 1669390400
transform 1 0 37856 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_330
timestamp 1669390400
transform 1 0 38304 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_340
timestamp 1669390400
transform 1 0 39424 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1669390400
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_357
timestamp 1669390400
transform 1 0 41328 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_359
timestamp 1669390400
transform 1 0 41552 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_366
timestamp 1669390400
transform 1 0 42336 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_370
timestamp 1669390400
transform 1 0 42784 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_374
timestamp 1669390400
transform 1 0 43232 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_378
timestamp 1669390400
transform 1 0 43680 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_382
timestamp 1669390400
transform 1 0 44128 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_385
timestamp 1669390400
transform 1 0 44464 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_389
timestamp 1669390400
transform 1 0 44912 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_391
timestamp 1669390400
transform 1 0 45136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_398
timestamp 1669390400
transform 1 0 45920 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_402
timestamp 1669390400
transform 1 0 46368 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_405
timestamp 1669390400
transform 1 0 46704 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_409
timestamp 1669390400
transform 1 0 47152 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_417
timestamp 1669390400
transform 1 0 48048 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_425
timestamp 1669390400
transform 1 0 48944 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_428
timestamp 1669390400
transform 1 0 49280 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_441
timestamp 1669390400
transform 1 0 50736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_447
timestamp 1669390400
transform 1 0 51408 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_451
timestamp 1669390400
transform 1 0 51856 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_461
timestamp 1669390400
transform 1 0 52976 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_465
timestamp 1669390400
transform 1 0 53424 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_467
timestamp 1669390400
transform 1 0 53648 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_476
timestamp 1669390400
transform 1 0 54656 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_493
timestamp 1669390400
transform 1 0 56560 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_499
timestamp 1669390400
transform 1 0 57232 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_506
timestamp 1669390400
transform 1 0 58016 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_508
timestamp 1669390400
transform 1 0 58240 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_2
timestamp 1669390400
transform 1 0 1568 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_6
timestamp 1669390400
transform 1 0 2016 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_10
timestamp 1669390400
transform 1 0 2464 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_14
timestamp 1669390400
transform 1 0 2912 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_18
timestamp 1669390400
transform 1 0 3360 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_22
timestamp 1669390400
transform 1 0 3808 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_26
timestamp 1669390400
transform 1 0 4256 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_30
timestamp 1669390400
transform 1 0 4704 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_34
timestamp 1669390400
transform 1 0 5152 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_37
timestamp 1669390400
transform 1 0 5488 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_39
timestamp 1669390400
transform 1 0 5712 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_42
timestamp 1669390400
transform 1 0 6048 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_52
timestamp 1669390400
transform 1 0 7168 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_62
timestamp 1669390400
transform 1 0 8288 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_64
timestamp 1669390400
transform 1 0 8512 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_77
timestamp 1669390400
transform 1 0 9968 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_88
timestamp 1669390400
transform 1 0 11200 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_97
timestamp 1669390400
transform 1 0 12208 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1669390400
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_108
timestamp 1669390400
transform 1 0 13440 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_122
timestamp 1669390400
transform 1 0 15008 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_128
timestamp 1669390400
transform 1 0 15680 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_136
timestamp 1669390400
transform 1 0 16576 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_138
timestamp 1669390400
transform 1 0 16800 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_141
timestamp 1669390400
transform 1 0 17136 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_145
timestamp 1669390400
transform 1 0 17584 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_151
timestamp 1669390400
transform 1 0 18256 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_161
timestamp 1669390400
transform 1 0 19376 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_171
timestamp 1669390400
transform 1 0 20496 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_173
timestamp 1669390400
transform 1 0 20720 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1669390400
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_179
timestamp 1669390400
transform 1 0 21392 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_181
timestamp 1669390400
transform 1 0 21616 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_184
timestamp 1669390400
transform 1 0 21952 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_190
timestamp 1669390400
transform 1 0 22624 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_202
timestamp 1669390400
transform 1 0 23968 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_210
timestamp 1669390400
transform 1 0 24864 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_214
timestamp 1669390400
transform 1 0 25312 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_218
timestamp 1669390400
transform 1 0 25760 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_220
timestamp 1669390400
transform 1 0 25984 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_227
timestamp 1669390400
transform 1 0 26768 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_231
timestamp 1669390400
transform 1 0 27216 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_239
timestamp 1669390400
transform 1 0 28112 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1669390400
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_250
timestamp 1669390400
transform 1 0 29344 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_253
timestamp 1669390400
transform 1 0 29680 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_265
timestamp 1669390400
transform 1 0 31024 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_269
timestamp 1669390400
transform 1 0 31472 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_273
timestamp 1669390400
transform 1 0 31920 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_289
timestamp 1669390400
transform 1 0 33712 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_295
timestamp 1669390400
transform 1 0 34384 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_299
timestamp 1669390400
transform 1 0 34832 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_303
timestamp 1669390400
transform 1 0 35280 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_316
timestamp 1669390400
transform 1 0 36736 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1669390400
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_321
timestamp 1669390400
transform 1 0 37296 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_328
timestamp 1669390400
transform 1 0 38080 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_332
timestamp 1669390400
transform 1 0 38528 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_334
timestamp 1669390400
transform 1 0 38752 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_341
timestamp 1669390400
transform 1 0 39536 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_345
timestamp 1669390400
transform 1 0 39984 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_347
timestamp 1669390400
transform 1 0 40208 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_354
timestamp 1669390400
transform 1 0 40992 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_358
timestamp 1669390400
transform 1 0 41440 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_362
timestamp 1669390400
transform 1 0 41888 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_375
timestamp 1669390400
transform 1 0 43344 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_383
timestamp 1669390400
transform 1 0 44240 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_387
timestamp 1669390400
transform 1 0 44688 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1669390400
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_392
timestamp 1669390400
transform 1 0 45248 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_398
timestamp 1669390400
transform 1 0 45920 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_400
timestamp 1669390400
transform 1 0 46144 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_403
timestamp 1669390400
transform 1 0 46480 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_407
timestamp 1669390400
transform 1 0 46928 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_411
timestamp 1669390400
transform 1 0 47376 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_415
timestamp 1669390400
transform 1 0 47824 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_419
timestamp 1669390400
transform 1 0 48272 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_425
timestamp 1669390400
transform 1 0 48944 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_427
timestamp 1669390400
transform 1 0 49168 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_434
timestamp 1669390400
transform 1 0 49952 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_438
timestamp 1669390400
transform 1 0 50400 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_442
timestamp 1669390400
transform 1 0 50848 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_446
timestamp 1669390400
transform 1 0 51296 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_448
timestamp 1669390400
transform 1 0 51520 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_459
timestamp 1669390400
transform 1 0 52752 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_463
timestamp 1669390400
transform 1 0 53200 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_471
timestamp 1669390400
transform 1 0 54096 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_475
timestamp 1669390400
transform 1 0 54544 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_491
timestamp 1669390400
transform 1 0 56336 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_499
timestamp 1669390400
transform 1 0 57232 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_14_507
timestamp 1669390400
transform 1 0 58128 0 1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_2
timestamp 1669390400
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_8
timestamp 1669390400
transform 1 0 2240 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_12
timestamp 1669390400
transform 1 0 2688 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_20
timestamp 1669390400
transform 1 0 3584 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_28
timestamp 1669390400
transform 1 0 4480 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_30
timestamp 1669390400
transform 1 0 4704 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_33
timestamp 1669390400
transform 1 0 5040 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_41
timestamp 1669390400
transform 1 0 5936 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_57
timestamp 1669390400
transform 1 0 7728 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_59
timestamp 1669390400
transform 1 0 7952 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_62
timestamp 1669390400
transform 1 0 8288 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_66
timestamp 1669390400
transform 1 0 8736 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1669390400
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_73
timestamp 1669390400
transform 1 0 9520 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_79
timestamp 1669390400
transform 1 0 10192 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_92
timestamp 1669390400
transform 1 0 11648 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_126
timestamp 1669390400
transform 1 0 15456 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_136
timestamp 1669390400
transform 1 0 16576 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_138
timestamp 1669390400
transform 1 0 16800 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1669390400
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_144
timestamp 1669390400
transform 1 0 17472 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_146
timestamp 1669390400
transform 1 0 17696 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_156
timestamp 1669390400
transform 1 0 18816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_160
timestamp 1669390400
transform 1 0 19264 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_184
timestamp 1669390400
transform 1 0 21952 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_190
timestamp 1669390400
transform 1 0 22624 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_198
timestamp 1669390400
transform 1 0 23520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_202
timestamp 1669390400
transform 1 0 23968 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_206
timestamp 1669390400
transform 1 0 24416 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1669390400
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_215
timestamp 1669390400
transform 1 0 25424 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_219
timestamp 1669390400
transform 1 0 25872 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_221
timestamp 1669390400
transform 1 0 26096 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_228
timestamp 1669390400
transform 1 0 26880 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_232
timestamp 1669390400
transform 1 0 27328 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_240
timestamp 1669390400
transform 1 0 28224 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_244
timestamp 1669390400
transform 1 0 28672 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_247
timestamp 1669390400
transform 1 0 29008 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_251
timestamp 1669390400
transform 1 0 29456 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_265
timestamp 1669390400
transform 1 0 31024 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_269
timestamp 1669390400
transform 1 0 31472 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_273
timestamp 1669390400
transform 1 0 31920 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1669390400
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_286
timestamp 1669390400
transform 1 0 33376 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_292
timestamp 1669390400
transform 1 0 34048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_296
timestamp 1669390400
transform 1 0 34496 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_298
timestamp 1669390400
transform 1 0 34720 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_301
timestamp 1669390400
transform 1 0 35056 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_305
timestamp 1669390400
transform 1 0 35504 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_315
timestamp 1669390400
transform 1 0 36624 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_323
timestamp 1669390400
transform 1 0 37520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_331
timestamp 1669390400
transform 1 0 38416 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_335
timestamp 1669390400
transform 1 0 38864 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_339
timestamp 1669390400
transform 1 0 39312 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_343
timestamp 1669390400
transform 1 0 39760 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_347
timestamp 1669390400
transform 1 0 40208 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_349
timestamp 1669390400
transform 1 0 40432 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_352
timestamp 1669390400
transform 1 0 40768 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1669390400
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_357
timestamp 1669390400
transform 1 0 41328 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_360
timestamp 1669390400
transform 1 0 41664 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_373
timestamp 1669390400
transform 1 0 43120 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_385
timestamp 1669390400
transform 1 0 44464 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_395
timestamp 1669390400
transform 1 0 45584 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_403
timestamp 1669390400
transform 1 0 46480 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_409
timestamp 1669390400
transform 1 0 47152 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_413
timestamp 1669390400
transform 1 0 47600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_423
timestamp 1669390400
transform 1 0 48720 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_425
timestamp 1669390400
transform 1 0 48944 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_428
timestamp 1669390400
transform 1 0 49280 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_431
timestamp 1669390400
transform 1 0 49616 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_433
timestamp 1669390400
transform 1 0 49840 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_444
timestamp 1669390400
transform 1 0 51072 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_448
timestamp 1669390400
transform 1 0 51520 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_458
timestamp 1669390400
transform 1 0 52640 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_466
timestamp 1669390400
transform 1 0 53536 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_470
timestamp 1669390400
transform 1 0 53984 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_480
timestamp 1669390400
transform 1 0 55104 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_496
timestamp 1669390400
transform 1 0 56896 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_499
timestamp 1669390400
transform 1 0 57232 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_506
timestamp 1669390400
transform 1 0 58016 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_508
timestamp 1669390400
transform 1 0 58240 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_2
timestamp 1669390400
transform 1 0 1568 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_6
timestamp 1669390400
transform 1 0 2016 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_10
timestamp 1669390400
transform 1 0 2464 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_14
timestamp 1669390400
transform 1 0 2912 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_18
timestamp 1669390400
transform 1 0 3360 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_22
timestamp 1669390400
transform 1 0 3808 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_26
timestamp 1669390400
transform 1 0 4256 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_30
timestamp 1669390400
transform 1 0 4704 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_34
timestamp 1669390400
transform 1 0 5152 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_37
timestamp 1669390400
transform 1 0 5488 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_44
timestamp 1669390400
transform 1 0 6272 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_48
timestamp 1669390400
transform 1 0 6720 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_60
timestamp 1669390400
transform 1 0 8064 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_64
timestamp 1669390400
transform 1 0 8512 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_68
timestamp 1669390400
transform 1 0 8960 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_76
timestamp 1669390400
transform 1 0 9856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_82
timestamp 1669390400
transform 1 0 10528 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_92
timestamp 1669390400
transform 1 0 11648 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_94
timestamp 1669390400
transform 1 0 11872 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_97
timestamp 1669390400
transform 1 0 12208 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_101
timestamp 1669390400
transform 1 0 12656 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1669390400
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_108
timestamp 1669390400
transform 1 0 13440 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_114
timestamp 1669390400
transform 1 0 14112 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_116
timestamp 1669390400
transform 1 0 14336 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_119
timestamp 1669390400
transform 1 0 14672 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_123
timestamp 1669390400
transform 1 0 15120 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_126
timestamp 1669390400
transform 1 0 15456 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_135
timestamp 1669390400
transform 1 0 16464 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_155
timestamp 1669390400
transform 1 0 18704 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_165
timestamp 1669390400
transform 1 0 19824 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_169
timestamp 1669390400
transform 1 0 20272 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_172
timestamp 1669390400
transform 1 0 20608 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1669390400
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_179
timestamp 1669390400
transform 1 0 21392 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_189
timestamp 1669390400
transform 1 0 22512 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_191
timestamp 1669390400
transform 1 0 22736 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_202
timestamp 1669390400
transform 1 0 23968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_206
timestamp 1669390400
transform 1 0 24416 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_209
timestamp 1669390400
transform 1 0 24752 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_217
timestamp 1669390400
transform 1 0 25648 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_227
timestamp 1669390400
transform 1 0 26768 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_231
timestamp 1669390400
transform 1 0 27216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_243
timestamp 1669390400
transform 1 0 28560 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1669390400
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_250
timestamp 1669390400
transform 1 0 29344 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_257
timestamp 1669390400
transform 1 0 30128 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_261
timestamp 1669390400
transform 1 0 30576 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_265
timestamp 1669390400
transform 1 0 31024 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_269
timestamp 1669390400
transform 1 0 31472 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_276
timestamp 1669390400
transform 1 0 32256 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_284
timestamp 1669390400
transform 1 0 33152 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_290
timestamp 1669390400
transform 1 0 33824 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_294
timestamp 1669390400
transform 1 0 34272 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_298
timestamp 1669390400
transform 1 0 34720 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_308
timestamp 1669390400
transform 1 0 35840 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_310
timestamp 1669390400
transform 1 0 36064 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_316
timestamp 1669390400
transform 1 0 36736 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1669390400
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_321
timestamp 1669390400
transform 1 0 37296 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_333
timestamp 1669390400
transform 1 0 38640 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_335
timestamp 1669390400
transform 1 0 38864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_342
timestamp 1669390400
transform 1 0 39648 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_346
timestamp 1669390400
transform 1 0 40096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_350
timestamp 1669390400
transform 1 0 40544 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_359
timestamp 1669390400
transform 1 0 41552 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_361
timestamp 1669390400
transform 1 0 41776 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_368
timestamp 1669390400
transform 1 0 42560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_372
timestamp 1669390400
transform 1 0 43008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_379
timestamp 1669390400
transform 1 0 43792 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_383
timestamp 1669390400
transform 1 0 44240 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_387
timestamp 1669390400
transform 1 0 44688 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1669390400
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_392
timestamp 1669390400
transform 1 0 45248 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_401
timestamp 1669390400
transform 1 0 46256 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_409
timestamp 1669390400
transform 1 0 47152 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_417
timestamp 1669390400
transform 1 0 48048 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_421
timestamp 1669390400
transform 1 0 48496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_432
timestamp 1669390400
transform 1 0 49728 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_442
timestamp 1669390400
transform 1 0 50848 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_444
timestamp 1669390400
transform 1 0 51072 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_460
timestamp 1669390400
transform 1 0 52864 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_463
timestamp 1669390400
transform 1 0 53200 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_474
timestamp 1669390400
transform 1 0 54432 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_478
timestamp 1669390400
transform 1 0 54880 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_490
timestamp 1669390400
transform 1 0 56224 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_498
timestamp 1669390400
transform 1 0 57120 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_502
timestamp 1669390400
transform 1 0 57568 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_16_506
timestamp 1669390400
transform 1 0 58016 0 1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_508
timestamp 1669390400
transform 1 0 58240 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_2
timestamp 1669390400
transform 1 0 1568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_8
timestamp 1669390400
transform 1 0 2240 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_12
timestamp 1669390400
transform 1 0 2688 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_16
timestamp 1669390400
transform 1 0 3136 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_20
timestamp 1669390400
transform 1 0 3584 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_24
timestamp 1669390400
transform 1 0 4032 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_32
timestamp 1669390400
transform 1 0 4928 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_47
timestamp 1669390400
transform 1 0 6608 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_60
timestamp 1669390400
transform 1 0 8064 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_66
timestamp 1669390400
transform 1 0 8736 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1669390400
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_73
timestamp 1669390400
transform 1 0 9520 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_80
timestamp 1669390400
transform 1 0 10304 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_88
timestamp 1669390400
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_92
timestamp 1669390400
transform 1 0 11648 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_95
timestamp 1669390400
transform 1 0 11984 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_99
timestamp 1669390400
transform 1 0 12432 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_119
timestamp 1669390400
transform 1 0 14672 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_127
timestamp 1669390400
transform 1 0 15568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_133
timestamp 1669390400
transform 1 0 16240 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_137
timestamp 1669390400
transform 1 0 16688 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1669390400
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_144
timestamp 1669390400
transform 1 0 17472 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_152
timestamp 1669390400
transform 1 0 18368 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_158
timestamp 1669390400
transform 1 0 19040 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_170
timestamp 1669390400
transform 1 0 20384 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_172
timestamp 1669390400
transform 1 0 20608 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_175
timestamp 1669390400
transform 1 0 20944 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_185
timestamp 1669390400
transform 1 0 22064 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_205
timestamp 1669390400
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_209
timestamp 1669390400
transform 1 0 24752 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1669390400
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_215
timestamp 1669390400
transform 1 0 25424 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_218
timestamp 1669390400
transform 1 0 25760 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_222
timestamp 1669390400
transform 1 0 26208 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_228
timestamp 1669390400
transform 1 0 26880 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_230
timestamp 1669390400
transform 1 0 27104 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_233
timestamp 1669390400
transform 1 0 27440 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_237
timestamp 1669390400
transform 1 0 27888 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_241
timestamp 1669390400
transform 1 0 28336 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_245
timestamp 1669390400
transform 1 0 28784 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_253
timestamp 1669390400
transform 1 0 29680 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_257
timestamp 1669390400
transform 1 0 30128 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_261
timestamp 1669390400
transform 1 0 30576 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_264
timestamp 1669390400
transform 1 0 30912 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_268
timestamp 1669390400
transform 1 0 31360 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_272
timestamp 1669390400
transform 1 0 31808 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_282
timestamp 1669390400
transform 1 0 32928 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_286
timestamp 1669390400
transform 1 0 33376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_292
timestamp 1669390400
transform 1 0 34048 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_296
timestamp 1669390400
transform 1 0 34496 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_300
timestamp 1669390400
transform 1 0 34944 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_313
timestamp 1669390400
transform 1 0 36400 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_317
timestamp 1669390400
transform 1 0 36848 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_321
timestamp 1669390400
transform 1 0 37296 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_325
timestamp 1669390400
transform 1 0 37744 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_329
timestamp 1669390400
transform 1 0 38192 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_339
timestamp 1669390400
transform 1 0 39312 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_341
timestamp 1669390400
transform 1 0 39536 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_352
timestamp 1669390400
transform 1 0 40768 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1669390400
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_357
timestamp 1669390400
transform 1 0 41328 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_360
timestamp 1669390400
transform 1 0 41664 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_364
timestamp 1669390400
transform 1 0 42112 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_368
timestamp 1669390400
transform 1 0 42560 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_372
timestamp 1669390400
transform 1 0 43008 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_374
timestamp 1669390400
transform 1 0 43232 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_377
timestamp 1669390400
transform 1 0 43568 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_381
timestamp 1669390400
transform 1 0 44016 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_388
timestamp 1669390400
transform 1 0 44800 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_398
timestamp 1669390400
transform 1 0 45920 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_402
timestamp 1669390400
transform 1 0 46368 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_404
timestamp 1669390400
transform 1 0 46592 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_411
timestamp 1669390400
transform 1 0 47376 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_413
timestamp 1669390400
transform 1 0 47600 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_422
timestamp 1669390400
transform 1 0 48608 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_428
timestamp 1669390400
transform 1 0 49280 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_446
timestamp 1669390400
transform 1 0 51296 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_450
timestamp 1669390400
transform 1 0 51744 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_454
timestamp 1669390400
transform 1 0 52192 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_456
timestamp 1669390400
transform 1 0 52416 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_471
timestamp 1669390400
transform 1 0 54096 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_481
timestamp 1669390400
transform 1 0 55216 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_485
timestamp 1669390400
transform 1 0 55664 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_492
timestamp 1669390400
transform 1 0 56448 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_496
timestamp 1669390400
transform 1 0 56896 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_499
timestamp 1669390400
transform 1 0 57232 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_506
timestamp 1669390400
transform 1 0 58016 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_508
timestamp 1669390400
transform 1 0 58240 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1669390400
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_19
timestamp 1669390400
transform 1 0 3472 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_23
timestamp 1669390400
transform 1 0 3920 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_26
timestamp 1669390400
transform 1 0 4256 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_30
timestamp 1669390400
transform 1 0 4704 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_34
timestamp 1669390400
transform 1 0 5152 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_37
timestamp 1669390400
transform 1 0 5488 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_43
timestamp 1669390400
transform 1 0 6160 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_47
timestamp 1669390400
transform 1 0 6608 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_58
timestamp 1669390400
transform 1 0 7840 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_71
timestamp 1669390400
transform 1 0 9296 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_81
timestamp 1669390400
transform 1 0 10416 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_95
timestamp 1669390400
transform 1 0 11984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_101
timestamp 1669390400
transform 1 0 12656 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1669390400
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_108
timestamp 1669390400
transform 1 0 13440 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_118
timestamp 1669390400
transform 1 0 14560 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_138
timestamp 1669390400
transform 1 0 16800 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_140
timestamp 1669390400
transform 1 0 17024 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_143
timestamp 1669390400
transform 1 0 17360 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_153
timestamp 1669390400
transform 1 0 18480 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_161
timestamp 1669390400
transform 1 0 19376 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_168
timestamp 1669390400
transform 1 0 20160 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_172
timestamp 1669390400
transform 1 0 20608 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1669390400
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_179
timestamp 1669390400
transform 1 0 21392 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_185
timestamp 1669390400
transform 1 0 22064 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_191
timestamp 1669390400
transform 1 0 22736 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_203
timestamp 1669390400
transform 1 0 24080 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_205
timestamp 1669390400
transform 1 0 24304 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_208
timestamp 1669390400
transform 1 0 24640 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_215
timestamp 1669390400
transform 1 0 25424 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_219
timestamp 1669390400
transform 1 0 25872 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_221
timestamp 1669390400
transform 1 0 26096 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_227
timestamp 1669390400
transform 1 0 26768 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_234
timestamp 1669390400
transform 1 0 27552 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_242
timestamp 1669390400
transform 1 0 28448 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_244
timestamp 1669390400
transform 1 0 28672 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1669390400
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_250
timestamp 1669390400
transform 1 0 29344 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_256
timestamp 1669390400
transform 1 0 30016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_262
timestamp 1669390400
transform 1 0 30688 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_269
timestamp 1669390400
transform 1 0 31472 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_281
timestamp 1669390400
transform 1 0 32816 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_289
timestamp 1669390400
transform 1 0 33712 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_293
timestamp 1669390400
transform 1 0 34160 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_299
timestamp 1669390400
transform 1 0 34832 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_301
timestamp 1669390400
transform 1 0 35056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_310
timestamp 1669390400
transform 1 0 36064 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_314
timestamp 1669390400
transform 1 0 36512 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1669390400
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_321
timestamp 1669390400
transform 1 0 37296 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_324
timestamp 1669390400
transform 1 0 37632 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_333
timestamp 1669390400
transform 1 0 38640 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_335
timestamp 1669390400
transform 1 0 38864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_338
timestamp 1669390400
transform 1 0 39200 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_344
timestamp 1669390400
transform 1 0 39872 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_346
timestamp 1669390400
transform 1 0 40096 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_359
timestamp 1669390400
transform 1 0 41552 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_369
timestamp 1669390400
transform 1 0 42672 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_373
timestamp 1669390400
transform 1 0 43120 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_377
timestamp 1669390400
transform 1 0 43568 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1669390400
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_392
timestamp 1669390400
transform 1 0 45248 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_399
timestamp 1669390400
transform 1 0 46032 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_403
timestamp 1669390400
transform 1 0 46480 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_407
timestamp 1669390400
transform 1 0 46928 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_411
timestamp 1669390400
transform 1 0 47376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_421
timestamp 1669390400
transform 1 0 48496 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_425
timestamp 1669390400
transform 1 0 48944 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_429
timestamp 1669390400
transform 1 0 49392 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_433
timestamp 1669390400
transform 1 0 49840 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_437
timestamp 1669390400
transform 1 0 50288 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_440
timestamp 1669390400
transform 1 0 50624 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_444
timestamp 1669390400
transform 1 0 51072 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_448
timestamp 1669390400
transform 1 0 51520 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_452
timestamp 1669390400
transform 1 0 51968 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_456
timestamp 1669390400
transform 1 0 52416 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_460
timestamp 1669390400
transform 1 0 52864 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_463
timestamp 1669390400
transform 1 0 53200 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_470
timestamp 1669390400
transform 1 0 53984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_480
timestamp 1669390400
transform 1 0 55104 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_487
timestamp 1669390400
transform 1 0 55888 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_497
timestamp 1669390400
transform 1 0 57008 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_505
timestamp 1669390400
transform 1 0 57904 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_2
timestamp 1669390400
transform 1 0 1568 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_5
timestamp 1669390400
transform 1 0 1904 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_9
timestamp 1669390400
transform 1 0 2352 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_13
timestamp 1669390400
transform 1 0 2800 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_23
timestamp 1669390400
transform 1 0 3920 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_35
timestamp 1669390400
transform 1 0 5264 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_45
timestamp 1669390400
transform 1 0 6384 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_55
timestamp 1669390400
transform 1 0 7504 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_66
timestamp 1669390400
transform 1 0 8736 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1669390400
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_73
timestamp 1669390400
transform 1 0 9520 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_76
timestamp 1669390400
transform 1 0 9856 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_86
timestamp 1669390400
transform 1 0 10976 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_92
timestamp 1669390400
transform 1 0 11648 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_96
timestamp 1669390400
transform 1 0 12096 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_100
timestamp 1669390400
transform 1 0 12544 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_104
timestamp 1669390400
transform 1 0 12992 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_108
timestamp 1669390400
transform 1 0 13440 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_115
timestamp 1669390400
transform 1 0 14224 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_122
timestamp 1669390400
transform 1 0 15008 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_134
timestamp 1669390400
transform 1 0 16352 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_138
timestamp 1669390400
transform 1 0 16800 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1669390400
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_144
timestamp 1669390400
transform 1 0 17472 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_169
timestamp 1669390400
transform 1 0 20272 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_179
timestamp 1669390400
transform 1 0 21392 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_187
timestamp 1669390400
transform 1 0 22288 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_193
timestamp 1669390400
transform 1 0 22960 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_207
timestamp 1669390400
transform 1 0 24528 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_209
timestamp 1669390400
transform 1 0 24752 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1669390400
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_215
timestamp 1669390400
transform 1 0 25424 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_219
timestamp 1669390400
transform 1 0 25872 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_227
timestamp 1669390400
transform 1 0 26768 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_231
timestamp 1669390400
transform 1 0 27216 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_239
timestamp 1669390400
transform 1 0 28112 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_243
timestamp 1669390400
transform 1 0 28560 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_247
timestamp 1669390400
transform 1 0 29008 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_255
timestamp 1669390400
transform 1 0 29904 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_259
timestamp 1669390400
transform 1 0 30352 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_261
timestamp 1669390400
transform 1 0 30576 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_272
timestamp 1669390400
transform 1 0 31808 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_282
timestamp 1669390400
transform 1 0 32928 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_286
timestamp 1669390400
transform 1 0 33376 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_297
timestamp 1669390400
transform 1 0 34608 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_301
timestamp 1669390400
transform 1 0 35056 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_305
timestamp 1669390400
transform 1 0 35504 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_311
timestamp 1669390400
transform 1 0 36176 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_313
timestamp 1669390400
transform 1 0 36400 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_324
timestamp 1669390400
transform 1 0 37632 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_328
timestamp 1669390400
transform 1 0 38080 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_331
timestamp 1669390400
transform 1 0 38416 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_339
timestamp 1669390400
transform 1 0 39312 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_343
timestamp 1669390400
transform 1 0 39760 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_345
timestamp 1669390400
transform 1 0 39984 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1669390400
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_357
timestamp 1669390400
transform 1 0 41328 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_359
timestamp 1669390400
transform 1 0 41552 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_369
timestamp 1669390400
transform 1 0 42672 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_373
timestamp 1669390400
transform 1 0 43120 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_377
timestamp 1669390400
transform 1 0 43568 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_379
timestamp 1669390400
transform 1 0 43792 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_385
timestamp 1669390400
transform 1 0 44464 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_389
timestamp 1669390400
transform 1 0 44912 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_401
timestamp 1669390400
transform 1 0 46256 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_409
timestamp 1669390400
transform 1 0 47152 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_415
timestamp 1669390400
transform 1 0 47824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_425
timestamp 1669390400
transform 1 0 48944 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_428
timestamp 1669390400
transform 1 0 49280 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_435
timestamp 1669390400
transform 1 0 50064 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_439
timestamp 1669390400
transform 1 0 50512 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_443
timestamp 1669390400
transform 1 0 50960 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_453
timestamp 1669390400
transform 1 0 52080 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_461
timestamp 1669390400
transform 1 0 52976 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_465
timestamp 1669390400
transform 1 0 53424 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_469
timestamp 1669390400
transform 1 0 53872 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_471
timestamp 1669390400
transform 1 0 54096 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_480
timestamp 1669390400
transform 1 0 55104 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_495
timestamp 1669390400
transform 1 0 56784 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_499
timestamp 1669390400
transform 1 0 57232 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_506
timestamp 1669390400
transform 1 0 58016 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_508
timestamp 1669390400
transform 1 0 58240 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_2
timestamp 1669390400
transform 1 0 1568 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_6
timestamp 1669390400
transform 1 0 2016 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_10
timestamp 1669390400
transform 1 0 2464 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_14
timestamp 1669390400
transform 1 0 2912 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_18
timestamp 1669390400
transform 1 0 3360 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_22
timestamp 1669390400
transform 1 0 3808 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_26
timestamp 1669390400
transform 1 0 4256 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_34
timestamp 1669390400
transform 1 0 5152 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_37
timestamp 1669390400
transform 1 0 5488 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_44
timestamp 1669390400
transform 1 0 6272 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_52
timestamp 1669390400
transform 1 0 7168 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_58
timestamp 1669390400
transform 1 0 7840 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_62
timestamp 1669390400
transform 1 0 8288 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_70
timestamp 1669390400
transform 1 0 9184 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_87
timestamp 1669390400
transform 1 0 11088 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_91
timestamp 1669390400
transform 1 0 11536 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_95
timestamp 1669390400
transform 1 0 11984 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1669390400
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_108
timestamp 1669390400
transform 1 0 13440 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_117
timestamp 1669390400
transform 1 0 14448 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_121
timestamp 1669390400
transform 1 0 14896 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_128
timestamp 1669390400
transform 1 0 15680 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_134
timestamp 1669390400
transform 1 0 16352 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_138
timestamp 1669390400
transform 1 0 16800 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_142
timestamp 1669390400
transform 1 0 17248 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_152
timestamp 1669390400
transform 1 0 18368 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_156
timestamp 1669390400
transform 1 0 18816 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1669390400
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_179
timestamp 1669390400
transform 1 0 21392 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_186
timestamp 1669390400
transform 1 0 22176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_200
timestamp 1669390400
transform 1 0 23744 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_202
timestamp 1669390400
transform 1 0 23968 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_205
timestamp 1669390400
transform 1 0 24304 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_209
timestamp 1669390400
transform 1 0 24752 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_212
timestamp 1669390400
transform 1 0 25088 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_216
timestamp 1669390400
transform 1 0 25536 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_220
timestamp 1669390400
transform 1 0 25984 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_230
timestamp 1669390400
transform 1 0 27104 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_239
timestamp 1669390400
transform 1 0 28112 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1669390400
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_250
timestamp 1669390400
transform 1 0 29344 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_257
timestamp 1669390400
transform 1 0 30128 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_264
timestamp 1669390400
transform 1 0 30912 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_268
timestamp 1669390400
transform 1 0 31360 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_274
timestamp 1669390400
transform 1 0 32032 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_276
timestamp 1669390400
transform 1 0 32256 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_279
timestamp 1669390400
transform 1 0 32592 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_283
timestamp 1669390400
transform 1 0 33040 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_287
timestamp 1669390400
transform 1 0 33488 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_291
timestamp 1669390400
transform 1 0 33936 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_295
timestamp 1669390400
transform 1 0 34384 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_305
timestamp 1669390400
transform 1 0 35504 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1669390400
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_321
timestamp 1669390400
transform 1 0 37296 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_331
timestamp 1669390400
transform 1 0 38416 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_346
timestamp 1669390400
transform 1 0 40096 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_354
timestamp 1669390400
transform 1 0 40992 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_356
timestamp 1669390400
transform 1 0 41216 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_365
timestamp 1669390400
transform 1 0 42224 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_369
timestamp 1669390400
transform 1 0 42672 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_373
timestamp 1669390400
transform 1 0 43120 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1669390400
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_392
timestamp 1669390400
transform 1 0 45248 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_405
timestamp 1669390400
transform 1 0 46704 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_409
timestamp 1669390400
transform 1 0 47152 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_430
timestamp 1669390400
transform 1 0 49504 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_438
timestamp 1669390400
transform 1 0 50400 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_442
timestamp 1669390400
transform 1 0 50848 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_457
timestamp 1669390400
transform 1 0 52528 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_463
timestamp 1669390400
transform 1 0 53200 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_474
timestamp 1669390400
transform 1 0 54432 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_478
timestamp 1669390400
transform 1 0 54880 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_488
timestamp 1669390400
transform 1 0 56000 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_492
timestamp 1669390400
transform 1 0 56448 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_494
timestamp 1669390400
transform 1 0 56672 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_20_501
timestamp 1669390400
transform 1 0 57456 0 1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_505
timestamp 1669390400
transform 1 0 57904 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_2
timestamp 1669390400
transform 1 0 1568 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_8
timestamp 1669390400
transform 1 0 2240 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_12
timestamp 1669390400
transform 1 0 2688 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_20
timestamp 1669390400
transform 1 0 3584 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_36
timestamp 1669390400
transform 1 0 5376 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_40
timestamp 1669390400
transform 1 0 5824 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_44
timestamp 1669390400
transform 1 0 6272 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_65
timestamp 1669390400
transform 1 0 8624 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_67
timestamp 1669390400
transform 1 0 8848 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1669390400
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_73
timestamp 1669390400
transform 1 0 9520 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_89
timestamp 1669390400
transform 1 0 11312 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_101
timestamp 1669390400
transform 1 0 12656 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_129
timestamp 1669390400
transform 1 0 15792 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_139
timestamp 1669390400
transform 1 0 16912 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1669390400
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_144
timestamp 1669390400
transform 1 0 17472 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_150
timestamp 1669390400
transform 1 0 18144 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_160
timestamp 1669390400
transform 1 0 19264 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_162
timestamp 1669390400
transform 1 0 19488 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_180
timestamp 1669390400
transform 1 0 21504 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_182
timestamp 1669390400
transform 1 0 21728 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_185
timestamp 1669390400
transform 1 0 22064 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_195
timestamp 1669390400
transform 1 0 23184 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_210
timestamp 1669390400
transform 1 0 24864 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1669390400
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_215
timestamp 1669390400
transform 1 0 25424 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_226
timestamp 1669390400
transform 1 0 26656 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_230
timestamp 1669390400
transform 1 0 27104 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_234
timestamp 1669390400
transform 1 0 27552 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_238
timestamp 1669390400
transform 1 0 28000 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_241
timestamp 1669390400
transform 1 0 28336 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_245
timestamp 1669390400
transform 1 0 28784 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_249
timestamp 1669390400
transform 1 0 29232 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_261
timestamp 1669390400
transform 1 0 30576 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_265
timestamp 1669390400
transform 1 0 31024 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_269
timestamp 1669390400
transform 1 0 31472 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_273
timestamp 1669390400
transform 1 0 31920 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_279
timestamp 1669390400
transform 1 0 32592 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1669390400
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_286
timestamp 1669390400
transform 1 0 33376 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_294
timestamp 1669390400
transform 1 0 34272 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_304
timestamp 1669390400
transform 1 0 35392 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_312
timestamp 1669390400
transform 1 0 36288 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_314
timestamp 1669390400
transform 1 0 36512 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_321
timestamp 1669390400
transform 1 0 37296 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_325
timestamp 1669390400
transform 1 0 37744 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_329
timestamp 1669390400
transform 1 0 38192 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_333
timestamp 1669390400
transform 1 0 38640 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_335
timestamp 1669390400
transform 1 0 38864 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_343
timestamp 1669390400
transform 1 0 39760 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_347
timestamp 1669390400
transform 1 0 40208 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_349
timestamp 1669390400
transform 1 0 40432 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_352
timestamp 1669390400
transform 1 0 40768 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1669390400
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_357
timestamp 1669390400
transform 1 0 41328 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_366
timestamp 1669390400
transform 1 0 42336 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_374
timestamp 1669390400
transform 1 0 43232 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_378
timestamp 1669390400
transform 1 0 43680 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_380
timestamp 1669390400
transform 1 0 43904 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_394
timestamp 1669390400
transform 1 0 45472 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_402
timestamp 1669390400
transform 1 0 46368 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_406
timestamp 1669390400
transform 1 0 46816 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_414
timestamp 1669390400
transform 1 0 47712 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_416
timestamp 1669390400
transform 1 0 47936 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_425
timestamp 1669390400
transform 1 0 48944 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_428
timestamp 1669390400
transform 1 0 49280 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_445
timestamp 1669390400
transform 1 0 51184 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_453
timestamp 1669390400
transform 1 0 52080 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_457
timestamp 1669390400
transform 1 0 52528 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_467
timestamp 1669390400
transform 1 0 53648 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_477
timestamp 1669390400
transform 1 0 54768 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_481
timestamp 1669390400
transform 1 0 55216 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_490
timestamp 1669390400
transform 1 0 56224 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_496
timestamp 1669390400
transform 1 0 56896 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_499
timestamp 1669390400
transform 1 0 57232 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_506
timestamp 1669390400
transform 1 0 58016 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_508
timestamp 1669390400
transform 1 0 58240 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_2
timestamp 1669390400
transform 1 0 1568 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_6
timestamp 1669390400
transform 1 0 2016 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_10
timestamp 1669390400
transform 1 0 2464 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_14
timestamp 1669390400
transform 1 0 2912 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_18
timestamp 1669390400
transform 1 0 3360 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_22
timestamp 1669390400
transform 1 0 3808 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_26
timestamp 1669390400
transform 1 0 4256 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_30
timestamp 1669390400
transform 1 0 4704 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1669390400
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_37
timestamp 1669390400
transform 1 0 5488 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_49
timestamp 1669390400
transform 1 0 6832 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_87
timestamp 1669390400
transform 1 0 11088 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_93
timestamp 1669390400
transform 1 0 11760 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_104
timestamp 1669390400
transform 1 0 12992 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_108
timestamp 1669390400
transform 1 0 13440 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_111
timestamp 1669390400
transform 1 0 13776 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_122
timestamp 1669390400
transform 1 0 15008 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_124
timestamp 1669390400
transform 1 0 15232 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_127
timestamp 1669390400
transform 1 0 15568 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_131
timestamp 1669390400
transform 1 0 16016 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_141
timestamp 1669390400
transform 1 0 17136 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_145
timestamp 1669390400
transform 1 0 17584 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_148
timestamp 1669390400
transform 1 0 17920 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_152
timestamp 1669390400
transform 1 0 18368 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_156
timestamp 1669390400
transform 1 0 18816 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_160
timestamp 1669390400
transform 1 0 19264 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_164
timestamp 1669390400
transform 1 0 19712 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1669390400
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_179
timestamp 1669390400
transform 1 0 21392 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_185
timestamp 1669390400
transform 1 0 22064 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_189
timestamp 1669390400
transform 1 0 22512 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_201
timestamp 1669390400
transform 1 0 23856 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_203
timestamp 1669390400
transform 1 0 24080 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_210
timestamp 1669390400
transform 1 0 24864 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_220
timestamp 1669390400
transform 1 0 25984 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_226
timestamp 1669390400
transform 1 0 26656 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_246
timestamp 1669390400
transform 1 0 28896 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_250
timestamp 1669390400
transform 1 0 29344 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_253
timestamp 1669390400
transform 1 0 29680 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_261
timestamp 1669390400
transform 1 0 30576 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_265
timestamp 1669390400
transform 1 0 31024 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_269
timestamp 1669390400
transform 1 0 31472 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_273
timestamp 1669390400
transform 1 0 31920 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_277
timestamp 1669390400
transform 1 0 32368 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_281
timestamp 1669390400
transform 1 0 32816 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_292
timestamp 1669390400
transform 1 0 34048 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_296
timestamp 1669390400
transform 1 0 34496 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_300
timestamp 1669390400
transform 1 0 34944 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_302
timestamp 1669390400
transform 1 0 35168 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_305
timestamp 1669390400
transform 1 0 35504 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_309
timestamp 1669390400
transform 1 0 35952 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_313
timestamp 1669390400
transform 1 0 36400 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_317
timestamp 1669390400
transform 1 0 36848 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_321
timestamp 1669390400
transform 1 0 37296 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_333
timestamp 1669390400
transform 1 0 38640 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_337
timestamp 1669390400
transform 1 0 39088 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_341
timestamp 1669390400
transform 1 0 39536 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_350
timestamp 1669390400
transform 1 0 40544 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_354
timestamp 1669390400
transform 1 0 40992 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_363
timestamp 1669390400
transform 1 0 42000 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_365
timestamp 1669390400
transform 1 0 42224 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_374
timestamp 1669390400
transform 1 0 43232 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_382
timestamp 1669390400
transform 1 0 44128 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_386
timestamp 1669390400
transform 1 0 44576 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_392
timestamp 1669390400
transform 1 0 45248 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_395
timestamp 1669390400
transform 1 0 45584 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_399
timestamp 1669390400
transform 1 0 46032 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_401
timestamp 1669390400
transform 1 0 46256 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_407
timestamp 1669390400
transform 1 0 46928 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_409
timestamp 1669390400
transform 1 0 47152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_416
timestamp 1669390400
transform 1 0 47936 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_420
timestamp 1669390400
transform 1 0 48384 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_424
timestamp 1669390400
transform 1 0 48832 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_428
timestamp 1669390400
transform 1 0 49280 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_432
timestamp 1669390400
transform 1 0 49728 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_436
timestamp 1669390400
transform 1 0 50176 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_440
timestamp 1669390400
transform 1 0 50624 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_444
timestamp 1669390400
transform 1 0 51072 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_453
timestamp 1669390400
transform 1 0 52080 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_457
timestamp 1669390400
transform 1 0 52528 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_463
timestamp 1669390400
transform 1 0 53200 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_466
timestamp 1669390400
transform 1 0 53536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_475
timestamp 1669390400
transform 1 0 54544 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_491
timestamp 1669390400
transform 1 0 56336 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_495
timestamp 1669390400
transform 1 0 56784 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_497
timestamp 1669390400
transform 1 0 57008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_502
timestamp 1669390400
transform 1 0 57568 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_22_506
timestamp 1669390400
transform 1 0 58016 0 1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_508
timestamp 1669390400
transform 1 0 58240 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_2
timestamp 1669390400
transform 1 0 1568 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_8
timestamp 1669390400
transform 1 0 2240 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_25
timestamp 1669390400
transform 1 0 4144 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_40
timestamp 1669390400
transform 1 0 5824 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_42
timestamp 1669390400
transform 1 0 6048 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_49
timestamp 1669390400
transform 1 0 6832 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_63
timestamp 1669390400
transform 1 0 8400 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_67
timestamp 1669390400
transform 1 0 8848 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_70
timestamp 1669390400
transform 1 0 9184 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_73
timestamp 1669390400
transform 1 0 9520 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_84
timestamp 1669390400
transform 1 0 10752 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_109
timestamp 1669390400
transform 1 0 13552 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_113
timestamp 1669390400
transform 1 0 14000 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_116
timestamp 1669390400
transform 1 0 14336 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_126
timestamp 1669390400
transform 1 0 15456 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_134
timestamp 1669390400
transform 1 0 16352 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1669390400
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_144
timestamp 1669390400
transform 1 0 17472 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_155
timestamp 1669390400
transform 1 0 18704 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_163
timestamp 1669390400
transform 1 0 19600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_169
timestamp 1669390400
transform 1 0 20272 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_182
timestamp 1669390400
transform 1 0 21728 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_192
timestamp 1669390400
transform 1 0 22848 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_194
timestamp 1669390400
transform 1 0 23072 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_200
timestamp 1669390400
transform 1 0 23744 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_204
timestamp 1669390400
transform 1 0 24192 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_208
timestamp 1669390400
transform 1 0 24640 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1669390400
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_215
timestamp 1669390400
transform 1 0 25424 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_221
timestamp 1669390400
transform 1 0 26096 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_231
timestamp 1669390400
transform 1 0 27216 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_243
timestamp 1669390400
transform 1 0 28560 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_253
timestamp 1669390400
transform 1 0 29680 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_261
timestamp 1669390400
transform 1 0 30576 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_265
timestamp 1669390400
transform 1 0 31024 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_269
timestamp 1669390400
transform 1 0 31472 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_275
timestamp 1669390400
transform 1 0 32144 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1669390400
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_286
timestamp 1669390400
transform 1 0 33376 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_300
timestamp 1669390400
transform 1 0 34944 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_302
timestamp 1669390400
transform 1 0 35168 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_313
timestamp 1669390400
transform 1 0 36400 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_317
timestamp 1669390400
transform 1 0 36848 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_321
timestamp 1669390400
transform 1 0 37296 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_325
timestamp 1669390400
transform 1 0 37744 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_329
timestamp 1669390400
transform 1 0 38192 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_331
timestamp 1669390400
transform 1 0 38416 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_334
timestamp 1669390400
transform 1 0 38752 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_338
timestamp 1669390400
transform 1 0 39200 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_342
timestamp 1669390400
transform 1 0 39648 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_352
timestamp 1669390400
transform 1 0 40768 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1669390400
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_357
timestamp 1669390400
transform 1 0 41328 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_360
timestamp 1669390400
transform 1 0 41664 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_364
timestamp 1669390400
transform 1 0 42112 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_406
timestamp 1669390400
transform 1 0 46816 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_418
timestamp 1669390400
transform 1 0 48160 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_422
timestamp 1669390400
transform 1 0 48608 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_428
timestamp 1669390400
transform 1 0 49280 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_431
timestamp 1669390400
transform 1 0 49616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_435
timestamp 1669390400
transform 1 0 50064 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_444
timestamp 1669390400
transform 1 0 51072 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_456
timestamp 1669390400
transform 1 0 52416 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_460
timestamp 1669390400
transform 1 0 52864 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_470
timestamp 1669390400
transform 1 0 53984 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_474
timestamp 1669390400
transform 1 0 54432 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_478
timestamp 1669390400
transform 1 0 54880 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_486
timestamp 1669390400
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_496
timestamp 1669390400
transform 1 0 56896 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_499
timestamp 1669390400
transform 1 0 57232 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_506
timestamp 1669390400
transform 1 0 58016 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_508
timestamp 1669390400
transform 1 0 58240 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_2
timestamp 1669390400
transform 1 0 1568 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_17
timestamp 1669390400
transform 1 0 3248 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_27
timestamp 1669390400
transform 1 0 4368 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_31
timestamp 1669390400
transform 1 0 4816 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1669390400
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_37
timestamp 1669390400
transform 1 0 5488 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_41
timestamp 1669390400
transform 1 0 5936 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_48
timestamp 1669390400
transform 1 0 6720 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_58
timestamp 1669390400
transform 1 0 7840 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_62
timestamp 1669390400
transform 1 0 8288 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_66
timestamp 1669390400
transform 1 0 8736 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_73
timestamp 1669390400
transform 1 0 9520 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_77
timestamp 1669390400
transform 1 0 9968 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_85
timestamp 1669390400
transform 1 0 10864 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_95
timestamp 1669390400
transform 1 0 11984 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_101
timestamp 1669390400
transform 1 0 12656 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1669390400
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_108
timestamp 1669390400
transform 1 0 13440 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_112
timestamp 1669390400
transform 1 0 13888 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_127
timestamp 1669390400
transform 1 0 15568 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_134
timestamp 1669390400
transform 1 0 16352 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_141
timestamp 1669390400
transform 1 0 17136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_145
timestamp 1669390400
transform 1 0 17584 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_148
timestamp 1669390400
transform 1 0 17920 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_161
timestamp 1669390400
transform 1 0 19376 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_165
timestamp 1669390400
transform 1 0 19824 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_174
timestamp 1669390400
transform 1 0 20832 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1669390400
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_179
timestamp 1669390400
transform 1 0 21392 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_194
timestamp 1669390400
transform 1 0 23072 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_196
timestamp 1669390400
transform 1 0 23296 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_203
timestamp 1669390400
transform 1 0 24080 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_238
timestamp 1669390400
transform 1 0 28000 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_245
timestamp 1669390400
transform 1 0 28784 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1669390400
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_250
timestamp 1669390400
transform 1 0 29344 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_259
timestamp 1669390400
transform 1 0 30352 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_263
timestamp 1669390400
transform 1 0 30800 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_269
timestamp 1669390400
transform 1 0 31472 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_280
timestamp 1669390400
transform 1 0 32704 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_282
timestamp 1669390400
transform 1 0 32928 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_289
timestamp 1669390400
transform 1 0 33712 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_291
timestamp 1669390400
transform 1 0 33936 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_298
timestamp 1669390400
transform 1 0 34720 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_302
timestamp 1669390400
transform 1 0 35168 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1669390400
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_321
timestamp 1669390400
transform 1 0 37296 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_332
timestamp 1669390400
transform 1 0 38528 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_342
timestamp 1669390400
transform 1 0 39648 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_352
timestamp 1669390400
transform 1 0 40768 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_356
timestamp 1669390400
transform 1 0 41216 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_360
timestamp 1669390400
transform 1 0 41664 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_375
timestamp 1669390400
transform 1 0 43344 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_383
timestamp 1669390400
transform 1 0 44240 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_387
timestamp 1669390400
transform 1 0 44688 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1669390400
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_392
timestamp 1669390400
transform 1 0 45248 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_404
timestamp 1669390400
transform 1 0 46592 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_414
timestamp 1669390400
transform 1 0 47712 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_418
timestamp 1669390400
transform 1 0 48160 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_427
timestamp 1669390400
transform 1 0 49168 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_429
timestamp 1669390400
transform 1 0 49392 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_443
timestamp 1669390400
transform 1 0 50960 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_457
timestamp 1669390400
transform 1 0 52528 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_463
timestamp 1669390400
transform 1 0 53200 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_470
timestamp 1669390400
transform 1 0 53984 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_474
timestamp 1669390400
transform 1 0 54432 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_490
timestamp 1669390400
transform 1 0 56224 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_498
timestamp 1669390400
transform 1 0 57120 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_506
timestamp 1669390400
transform 1 0 58016 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_508
timestamp 1669390400
transform 1 0 58240 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1669390400
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_5
timestamp 1669390400
transform 1 0 1904 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_9
timestamp 1669390400
transform 1 0 2352 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_58
timestamp 1669390400
transform 1 0 7840 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_66
timestamp 1669390400
transform 1 0 8736 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_70
timestamp 1669390400
transform 1 0 9184 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_73
timestamp 1669390400
transform 1 0 9520 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_114
timestamp 1669390400
transform 1 0 14112 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_131
timestamp 1669390400
transform 1 0 16016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_137
timestamp 1669390400
transform 1 0 16688 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1669390400
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_144
timestamp 1669390400
transform 1 0 17472 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_153
timestamp 1669390400
transform 1 0 18480 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_157
timestamp 1669390400
transform 1 0 18928 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_160
timestamp 1669390400
transform 1 0 19264 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_164
timestamp 1669390400
transform 1 0 19712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_179
timestamp 1669390400
transform 1 0 21392 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_188
timestamp 1669390400
transform 1 0 22400 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_192
timestamp 1669390400
transform 1 0 22848 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_196
timestamp 1669390400
transform 1 0 23296 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_206
timestamp 1669390400
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1669390400
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_215
timestamp 1669390400
transform 1 0 25424 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_224
timestamp 1669390400
transform 1 0 26432 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_241
timestamp 1669390400
transform 1 0 28336 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_249
timestamp 1669390400
transform 1 0 29232 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_253
timestamp 1669390400
transform 1 0 29680 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_257
timestamp 1669390400
transform 1 0 30128 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_261
timestamp 1669390400
transform 1 0 30576 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_274
timestamp 1669390400
transform 1 0 32032 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1669390400
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_286
timestamp 1669390400
transform 1 0 33376 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_289
timestamp 1669390400
transform 1 0 33712 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_293
timestamp 1669390400
transform 1 0 34160 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_303
timestamp 1669390400
transform 1 0 35280 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_316
timestamp 1669390400
transform 1 0 36736 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_320
timestamp 1669390400
transform 1 0 37184 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_330
timestamp 1669390400
transform 1 0 38304 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_334
timestamp 1669390400
transform 1 0 38752 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_338
timestamp 1669390400
transform 1 0 39200 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_350
timestamp 1669390400
transform 1 0 40544 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1669390400
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_357
timestamp 1669390400
transform 1 0 41328 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_364
timestamp 1669390400
transform 1 0 42112 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_368
timestamp 1669390400
transform 1 0 42560 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_380
timestamp 1669390400
transform 1 0 43904 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_382
timestamp 1669390400
transform 1 0 44128 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_388
timestamp 1669390400
transform 1 0 44800 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_395
timestamp 1669390400
transform 1 0 45584 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_399
timestamp 1669390400
transform 1 0 46032 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_401
timestamp 1669390400
transform 1 0 46256 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_408
timestamp 1669390400
transform 1 0 47040 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_412
timestamp 1669390400
transform 1 0 47488 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_416
timestamp 1669390400
transform 1 0 47936 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_420
timestamp 1669390400
transform 1 0 48384 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_424
timestamp 1669390400
transform 1 0 48832 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_428
timestamp 1669390400
transform 1 0 49280 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_436
timestamp 1669390400
transform 1 0 50176 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_438
timestamp 1669390400
transform 1 0 50400 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_445
timestamp 1669390400
transform 1 0 51184 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_449
timestamp 1669390400
transform 1 0 51632 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_453
timestamp 1669390400
transform 1 0 52080 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_470
timestamp 1669390400
transform 1 0 53984 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_477
timestamp 1669390400
transform 1 0 54768 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_484
timestamp 1669390400
transform 1 0 55552 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_494
timestamp 1669390400
transform 1 0 56672 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_496
timestamp 1669390400
transform 1 0 56896 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_499
timestamp 1669390400
transform 1 0 57232 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_506
timestamp 1669390400
transform 1 0 58016 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_508
timestamp 1669390400
transform 1 0 58240 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_2
timestamp 1669390400
transform 1 0 1568 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_11
timestamp 1669390400
transform 1 0 2576 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_21
timestamp 1669390400
transform 1 0 3696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_25
timestamp 1669390400
transform 1 0 4144 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1669390400
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_37
timestamp 1669390400
transform 1 0 5488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_43
timestamp 1669390400
transform 1 0 6160 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_53
timestamp 1669390400
transform 1 0 7280 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_61
timestamp 1669390400
transform 1 0 8176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_65
timestamp 1669390400
transform 1 0 8624 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_68
timestamp 1669390400
transform 1 0 8960 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_86
timestamp 1669390400
transform 1 0 10976 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_102
timestamp 1669390400
transform 1 0 12768 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_108
timestamp 1669390400
transform 1 0 13440 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_115
timestamp 1669390400
transform 1 0 14224 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_123
timestamp 1669390400
transform 1 0 15120 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_130
timestamp 1669390400
transform 1 0 15904 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_132
timestamp 1669390400
transform 1 0 16128 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_144
timestamp 1669390400
transform 1 0 17472 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_156
timestamp 1669390400
transform 1 0 18816 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_158
timestamp 1669390400
transform 1 0 19040 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_169
timestamp 1669390400
transform 1 0 20272 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1669390400
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_179
timestamp 1669390400
transform 1 0 21392 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_182
timestamp 1669390400
transform 1 0 21728 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_197
timestamp 1669390400
transform 1 0 23408 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_222
timestamp 1669390400
transform 1 0 26208 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_226
timestamp 1669390400
transform 1 0 26656 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_229
timestamp 1669390400
transform 1 0 26992 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_233
timestamp 1669390400
transform 1 0 27440 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_240
timestamp 1669390400
transform 1 0 28224 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_246
timestamp 1669390400
transform 1 0 28896 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_250
timestamp 1669390400
transform 1 0 29344 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_253
timestamp 1669390400
transform 1 0 29680 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_257
timestamp 1669390400
transform 1 0 30128 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_259
timestamp 1669390400
transform 1 0 30352 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_273
timestamp 1669390400
transform 1 0 31920 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_277
timestamp 1669390400
transform 1 0 32368 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_280
timestamp 1669390400
transform 1 0 32704 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_292
timestamp 1669390400
transform 1 0 34048 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_299
timestamp 1669390400
transform 1 0 34832 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_301
timestamp 1669390400
transform 1 0 35056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_308
timestamp 1669390400
transform 1 0 35840 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_312
timestamp 1669390400
transform 1 0 36288 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_316
timestamp 1669390400
transform 1 0 36736 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1669390400
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_321
timestamp 1669390400
transform 1 0 37296 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_324
timestamp 1669390400
transform 1 0 37632 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_328
timestamp 1669390400
transform 1 0 38080 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_332
timestamp 1669390400
transform 1 0 38528 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_334
timestamp 1669390400
transform 1 0 38752 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_337
timestamp 1669390400
transform 1 0 39088 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_341
timestamp 1669390400
transform 1 0 39536 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_345
timestamp 1669390400
transform 1 0 39984 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_349
timestamp 1669390400
transform 1 0 40432 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_353
timestamp 1669390400
transform 1 0 40880 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_357
timestamp 1669390400
transform 1 0 41328 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_361
timestamp 1669390400
transform 1 0 41776 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_365
timestamp 1669390400
transform 1 0 42224 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_375
timestamp 1669390400
transform 1 0 43344 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_379
timestamp 1669390400
transform 1 0 43792 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_383
timestamp 1669390400
transform 1 0 44240 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_387
timestamp 1669390400
transform 1 0 44688 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1669390400
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_392
timestamp 1669390400
transform 1 0 45248 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_401
timestamp 1669390400
transform 1 0 46256 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_403
timestamp 1669390400
transform 1 0 46480 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_412
timestamp 1669390400
transform 1 0 47488 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_416
timestamp 1669390400
transform 1 0 47936 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_426
timestamp 1669390400
transform 1 0 49056 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_435
timestamp 1669390400
transform 1 0 50064 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_443
timestamp 1669390400
transform 1 0 50960 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_453
timestamp 1669390400
transform 1 0 52080 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_457
timestamp 1669390400
transform 1 0 52528 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_463
timestamp 1669390400
transform 1 0 53200 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_472
timestamp 1669390400
transform 1 0 54208 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_476
timestamp 1669390400
transform 1 0 54656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_490
timestamp 1669390400
transform 1 0 56224 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_502
timestamp 1669390400
transform 1 0 57568 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_506
timestamp 1669390400
transform 1 0 58016 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_508
timestamp 1669390400
transform 1 0 58240 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_2
timestamp 1669390400
transform 1 0 1568 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_6
timestamp 1669390400
transform 1 0 2016 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_10
timestamp 1669390400
transform 1 0 2464 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_20
timestamp 1669390400
transform 1 0 3584 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_65
timestamp 1669390400
transform 1 0 8624 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_67
timestamp 1669390400
transform 1 0 8848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_70
timestamp 1669390400
transform 1 0 9184 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_73
timestamp 1669390400
transform 1 0 9520 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_88
timestamp 1669390400
transform 1 0 11200 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_92
timestamp 1669390400
transform 1 0 11648 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_104
timestamp 1669390400
transform 1 0 12992 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_106
timestamp 1669390400
transform 1 0 13216 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_115
timestamp 1669390400
transform 1 0 14224 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_121
timestamp 1669390400
transform 1 0 14896 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_125
timestamp 1669390400
transform 1 0 15344 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_129
timestamp 1669390400
transform 1 0 15792 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_133
timestamp 1669390400
transform 1 0 16240 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_137
timestamp 1669390400
transform 1 0 16688 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1669390400
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_144
timestamp 1669390400
transform 1 0 17472 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_152
timestamp 1669390400
transform 1 0 18368 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_154
timestamp 1669390400
transform 1 0 18592 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_157
timestamp 1669390400
transform 1 0 18928 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_161
timestamp 1669390400
transform 1 0 19376 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_165
timestamp 1669390400
transform 1 0 19824 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_207
timestamp 1669390400
transform 1 0 24528 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_209
timestamp 1669390400
transform 1 0 24752 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1669390400
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_215
timestamp 1669390400
transform 1 0 25424 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_222
timestamp 1669390400
transform 1 0 26208 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_226
timestamp 1669390400
transform 1 0 26656 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_235
timestamp 1669390400
transform 1 0 27664 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_245
timestamp 1669390400
transform 1 0 28784 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_253
timestamp 1669390400
transform 1 0 29680 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_257
timestamp 1669390400
transform 1 0 30128 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_261
timestamp 1669390400
transform 1 0 30576 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_265
timestamp 1669390400
transform 1 0 31024 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_269
timestamp 1669390400
transform 1 0 31472 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_272
timestamp 1669390400
transform 1 0 31808 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_276
timestamp 1669390400
transform 1 0 32256 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_279
timestamp 1669390400
transform 1 0 32592 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1669390400
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_286
timestamp 1669390400
transform 1 0 33376 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_289
timestamp 1669390400
transform 1 0 33712 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_293
timestamp 1669390400
transform 1 0 34160 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_297
timestamp 1669390400
transform 1 0 34608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_303
timestamp 1669390400
transform 1 0 35280 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_307
timestamp 1669390400
transform 1 0 35728 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_311
timestamp 1669390400
transform 1 0 36176 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_315
timestamp 1669390400
transform 1 0 36624 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_317
timestamp 1669390400
transform 1 0 36848 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_327
timestamp 1669390400
transform 1 0 37968 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_331
timestamp 1669390400
transform 1 0 38416 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_333
timestamp 1669390400
transform 1 0 38640 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_336
timestamp 1669390400
transform 1 0 38976 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_350
timestamp 1669390400
transform 1 0 40544 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1669390400
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_357
timestamp 1669390400
transform 1 0 41328 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_360
timestamp 1669390400
transform 1 0 41664 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_364
timestamp 1669390400
transform 1 0 42112 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_368
timestamp 1669390400
transform 1 0 42560 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_375
timestamp 1669390400
transform 1 0 43344 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_400
timestamp 1669390400
transform 1 0 46144 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_420
timestamp 1669390400
transform 1 0 48384 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_424
timestamp 1669390400
transform 1 0 48832 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_428
timestamp 1669390400
transform 1 0 49280 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_452
timestamp 1669390400
transform 1 0 51968 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_454
timestamp 1669390400
transform 1 0 52192 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_463
timestamp 1669390400
transform 1 0 53200 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_474
timestamp 1669390400
transform 1 0 54432 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_482
timestamp 1669390400
transform 1 0 55328 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_484
timestamp 1669390400
transform 1 0 55552 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_491
timestamp 1669390400
transform 1 0 56336 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_495
timestamp 1669390400
transform 1 0 56784 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_499
timestamp 1669390400
transform 1 0 57232 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_508
timestamp 1669390400
transform 1 0 58240 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_2
timestamp 1669390400
transform 1 0 1568 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_6
timestamp 1669390400
transform 1 0 2016 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_10
timestamp 1669390400
transform 1 0 2464 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_14
timestamp 1669390400
transform 1 0 2912 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_18
timestamp 1669390400
transform 1 0 3360 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_22
timestamp 1669390400
transform 1 0 3808 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_26
timestamp 1669390400
transform 1 0 4256 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_30
timestamp 1669390400
transform 1 0 4704 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1669390400
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_37
timestamp 1669390400
transform 1 0 5488 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_44
timestamp 1669390400
transform 1 0 6272 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_69
timestamp 1669390400
transform 1 0 9072 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_71
timestamp 1669390400
transform 1 0 9296 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_74
timestamp 1669390400
transform 1 0 9632 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_84
timestamp 1669390400
transform 1 0 10752 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_94
timestamp 1669390400
transform 1 0 11872 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_98
timestamp 1669390400
transform 1 0 12320 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_101
timestamp 1669390400
transform 1 0 12656 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1669390400
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_108
timestamp 1669390400
transform 1 0 13440 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_119
timestamp 1669390400
transform 1 0 14672 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_128
timestamp 1669390400
transform 1 0 15680 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_132
timestamp 1669390400
transform 1 0 16128 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_136
timestamp 1669390400
transform 1 0 16576 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_140
timestamp 1669390400
transform 1 0 17024 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_148
timestamp 1669390400
transform 1 0 17920 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_154
timestamp 1669390400
transform 1 0 18592 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_158
timestamp 1669390400
transform 1 0 19040 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_170
timestamp 1669390400
transform 1 0 20384 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1669390400
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_179
timestamp 1669390400
transform 1 0 21392 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_187
timestamp 1669390400
transform 1 0 22288 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_191
timestamp 1669390400
transform 1 0 22736 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_201
timestamp 1669390400
transform 1 0 23856 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_211
timestamp 1669390400
transform 1 0 24976 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_218
timestamp 1669390400
transform 1 0 25760 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_225
timestamp 1669390400
transform 1 0 26544 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_229
timestamp 1669390400
transform 1 0 26992 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_238
timestamp 1669390400
transform 1 0 28000 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_242
timestamp 1669390400
transform 1 0 28448 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_244
timestamp 1669390400
transform 1 0 28672 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1669390400
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_250
timestamp 1669390400
transform 1 0 29344 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_253
timestamp 1669390400
transform 1 0 29680 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_257
timestamp 1669390400
transform 1 0 30128 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_261
timestamp 1669390400
transform 1 0 30576 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_270
timestamp 1669390400
transform 1 0 31584 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_278
timestamp 1669390400
transform 1 0 32480 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_282
timestamp 1669390400
transform 1 0 32928 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_284
timestamp 1669390400
transform 1 0 33152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_291
timestamp 1669390400
transform 1 0 33936 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_303
timestamp 1669390400
transform 1 0 35280 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_310
timestamp 1669390400
transform 1 0 36064 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_312
timestamp 1669390400
transform 1 0 36288 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1669390400
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_321
timestamp 1669390400
transform 1 0 37296 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_332
timestamp 1669390400
transform 1 0 38528 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_336
timestamp 1669390400
transform 1 0 38976 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_338
timestamp 1669390400
transform 1 0 39200 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_343
timestamp 1669390400
transform 1 0 39760 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_356
timestamp 1669390400
transform 1 0 41216 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_360
timestamp 1669390400
transform 1 0 41664 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_364
timestamp 1669390400
transform 1 0 42112 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_366
timestamp 1669390400
transform 1 0 42336 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_376
timestamp 1669390400
transform 1 0 43456 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_383
timestamp 1669390400
transform 1 0 44240 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_387
timestamp 1669390400
transform 1 0 44688 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1669390400
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_392
timestamp 1669390400
transform 1 0 45248 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_401
timestamp 1669390400
transform 1 0 46256 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_409
timestamp 1669390400
transform 1 0 47152 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_413
timestamp 1669390400
transform 1 0 47600 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_415
timestamp 1669390400
transform 1 0 47824 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_421
timestamp 1669390400
transform 1 0 48496 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_429
timestamp 1669390400
transform 1 0 49392 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_449
timestamp 1669390400
transform 1 0 51632 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_453
timestamp 1669390400
transform 1 0 52080 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_457
timestamp 1669390400
transform 1 0 52528 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_463
timestamp 1669390400
transform 1 0 53200 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_28_500
timestamp 1669390400
transform 1 0 57344 0 1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_508
timestamp 1669390400
transform 1 0 58240 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_2
timestamp 1669390400
transform 1 0 1568 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_8
timestamp 1669390400
transform 1 0 2240 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_12
timestamp 1669390400
transform 1 0 2688 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_16
timestamp 1669390400
transform 1 0 3136 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_24
timestamp 1669390400
transform 1 0 4032 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_32
timestamp 1669390400
transform 1 0 4928 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_34
timestamp 1669390400
transform 1 0 5152 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_37
timestamp 1669390400
transform 1 0 5488 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_41
timestamp 1669390400
transform 1 0 5936 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_45
timestamp 1669390400
transform 1 0 6384 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_55
timestamp 1669390400
transform 1 0 7504 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_57
timestamp 1669390400
transform 1 0 7728 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_60
timestamp 1669390400
transform 1 0 8064 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1669390400
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_73
timestamp 1669390400
transform 1 0 9520 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_79
timestamp 1669390400
transform 1 0 10192 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_89
timestamp 1669390400
transform 1 0 11312 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_95
timestamp 1669390400
transform 1 0 11984 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_99
timestamp 1669390400
transform 1 0 12432 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_111
timestamp 1669390400
transform 1 0 13776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_115
timestamp 1669390400
transform 1 0 14224 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_122
timestamp 1669390400
transform 1 0 15008 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_129
timestamp 1669390400
transform 1 0 15792 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1669390400
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_144
timestamp 1669390400
transform 1 0 17472 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_150
timestamp 1669390400
transform 1 0 18144 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_164
timestamp 1669390400
transform 1 0 19712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_208
timestamp 1669390400
transform 1 0 24640 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1669390400
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_215
timestamp 1669390400
transform 1 0 25424 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_224
timestamp 1669390400
transform 1 0 26432 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_228
timestamp 1669390400
transform 1 0 26880 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_237
timestamp 1669390400
transform 1 0 27888 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_245
timestamp 1669390400
transform 1 0 28784 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_249
timestamp 1669390400
transform 1 0 29232 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_253
timestamp 1669390400
transform 1 0 29680 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_257
timestamp 1669390400
transform 1 0 30128 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_261
timestamp 1669390400
transform 1 0 30576 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_280
timestamp 1669390400
transform 1 0 32704 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_286
timestamp 1669390400
transform 1 0 33376 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_289
timestamp 1669390400
transform 1 0 33712 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_301
timestamp 1669390400
transform 1 0 35056 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_311
timestamp 1669390400
transform 1 0 36176 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_315
timestamp 1669390400
transform 1 0 36624 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_319
timestamp 1669390400
transform 1 0 37072 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_331
timestamp 1669390400
transform 1 0 38416 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_341
timestamp 1669390400
transform 1 0 39536 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_343
timestamp 1669390400
transform 1 0 39760 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1669390400
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_357
timestamp 1669390400
transform 1 0 41328 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_366
timestamp 1669390400
transform 1 0 42336 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_376
timestamp 1669390400
transform 1 0 43456 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_385
timestamp 1669390400
transform 1 0 44464 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_387
timestamp 1669390400
transform 1 0 44688 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_393
timestamp 1669390400
transform 1 0 45360 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_397
timestamp 1669390400
transform 1 0 45808 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_401
timestamp 1669390400
transform 1 0 46256 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_409
timestamp 1669390400
transform 1 0 47152 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_419
timestamp 1669390400
transform 1 0 48272 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_423
timestamp 1669390400
transform 1 0 48720 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_425
timestamp 1669390400
transform 1 0 48944 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_428
timestamp 1669390400
transform 1 0 49280 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_430
timestamp 1669390400
transform 1 0 49504 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_439
timestamp 1669390400
transform 1 0 50512 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_443
timestamp 1669390400
transform 1 0 50960 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_447
timestamp 1669390400
transform 1 0 51408 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_451
timestamp 1669390400
transform 1 0 51856 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_455
timestamp 1669390400
transform 1 0 52304 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_462
timestamp 1669390400
transform 1 0 53088 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_472
timestamp 1669390400
transform 1 0 54208 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_476
timestamp 1669390400
transform 1 0 54656 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_491
timestamp 1669390400
transform 1 0 56336 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_495
timestamp 1669390400
transform 1 0 56784 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_499
timestamp 1669390400
transform 1 0 57232 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_508
timestamp 1669390400
transform 1 0 58240 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_2
timestamp 1669390400
transform 1 0 1568 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_8
timestamp 1669390400
transform 1 0 2240 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_12
timestamp 1669390400
transform 1 0 2688 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_16
timestamp 1669390400
transform 1 0 3136 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_20
timestamp 1669390400
transform 1 0 3584 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_24
timestamp 1669390400
transform 1 0 4032 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_34
timestamp 1669390400
transform 1 0 5152 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_37
timestamp 1669390400
transform 1 0 5488 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_46
timestamp 1669390400
transform 1 0 6496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_55
timestamp 1669390400
transform 1 0 7504 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_61
timestamp 1669390400
transform 1 0 8176 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_65
timestamp 1669390400
transform 1 0 8624 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_69
timestamp 1669390400
transform 1 0 9072 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_73
timestamp 1669390400
transform 1 0 9520 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_84
timestamp 1669390400
transform 1 0 10752 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_92
timestamp 1669390400
transform 1 0 11648 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_96
timestamp 1669390400
transform 1 0 12096 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1669390400
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_108
timestamp 1669390400
transform 1 0 13440 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_110
timestamp 1669390400
transform 1 0 13664 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_113
timestamp 1669390400
transform 1 0 14000 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_127
timestamp 1669390400
transform 1 0 15568 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_129
timestamp 1669390400
transform 1 0 15792 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_132
timestamp 1669390400
transform 1 0 16128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_143
timestamp 1669390400
transform 1 0 17360 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_147
timestamp 1669390400
transform 1 0 17808 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_150
timestamp 1669390400
transform 1 0 18144 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_154
timestamp 1669390400
transform 1 0 18592 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_158
timestamp 1669390400
transform 1 0 19040 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_162
timestamp 1669390400
transform 1 0 19488 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1669390400
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_179
timestamp 1669390400
transform 1 0 21392 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_183
timestamp 1669390400
transform 1 0 21840 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_187
timestamp 1669390400
transform 1 0 22288 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_191
timestamp 1669390400
transform 1 0 22736 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_203
timestamp 1669390400
transform 1 0 24080 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_213
timestamp 1669390400
transform 1 0 25200 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_233
timestamp 1669390400
transform 1 0 27440 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_237
timestamp 1669390400
transform 1 0 27888 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_241
timestamp 1669390400
transform 1 0 28336 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_245
timestamp 1669390400
transform 1 0 28784 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1669390400
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_250
timestamp 1669390400
transform 1 0 29344 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_254
timestamp 1669390400
transform 1 0 29792 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_261
timestamp 1669390400
transform 1 0 30576 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_273
timestamp 1669390400
transform 1 0 31920 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_281
timestamp 1669390400
transform 1 0 32816 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_285
timestamp 1669390400
transform 1 0 33264 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_297
timestamp 1669390400
transform 1 0 34608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_301
timestamp 1669390400
transform 1 0 35056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_304
timestamp 1669390400
transform 1 0 35392 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_308
timestamp 1669390400
transform 1 0 35840 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_312
timestamp 1669390400
transform 1 0 36288 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_316
timestamp 1669390400
transform 1 0 36736 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1669390400
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_321
timestamp 1669390400
transform 1 0 37296 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_328
timestamp 1669390400
transform 1 0 38080 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_335
timestamp 1669390400
transform 1 0 38864 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_339
timestamp 1669390400
transform 1 0 39312 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_343
timestamp 1669390400
transform 1 0 39760 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_363
timestamp 1669390400
transform 1 0 42000 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_367
timestamp 1669390400
transform 1 0 42448 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_371
timestamp 1669390400
transform 1 0 42896 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_386
timestamp 1669390400
transform 1 0 44576 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_392
timestamp 1669390400
transform 1 0 45248 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_399
timestamp 1669390400
transform 1 0 46032 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_403
timestamp 1669390400
transform 1 0 46480 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_413
timestamp 1669390400
transform 1 0 47600 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_417
timestamp 1669390400
transform 1 0 48048 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_421
timestamp 1669390400
transform 1 0 48496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_431
timestamp 1669390400
transform 1 0 49616 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_438
timestamp 1669390400
transform 1 0 50400 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_442
timestamp 1669390400
transform 1 0 50848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_446
timestamp 1669390400
transform 1 0 51296 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_453
timestamp 1669390400
transform 1 0 52080 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_457
timestamp 1669390400
transform 1 0 52528 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_463
timestamp 1669390400
transform 1 0 53200 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_465
timestamp 1669390400
transform 1 0 53424 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_482
timestamp 1669390400
transform 1 0 55328 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_492
timestamp 1669390400
transform 1 0 56448 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_496
timestamp 1669390400
transform 1 0 56896 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_503
timestamp 1669390400
transform 1 0 57680 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_507
timestamp 1669390400
transform 1 0 58128 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_2
timestamp 1669390400
transform 1 0 1568 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_5
timestamp 1669390400
transform 1 0 1904 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_9
timestamp 1669390400
transform 1 0 2352 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_13
timestamp 1669390400
transform 1 0 2800 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_17
timestamp 1669390400
transform 1 0 3248 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_21
timestamp 1669390400
transform 1 0 3696 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_25
timestamp 1669390400
transform 1 0 4144 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_29
timestamp 1669390400
transform 1 0 4592 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_33
timestamp 1669390400
transform 1 0 5040 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_37
timestamp 1669390400
transform 1 0 5488 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_41
timestamp 1669390400
transform 1 0 5936 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_49
timestamp 1669390400
transform 1 0 6832 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_60
timestamp 1669390400
transform 1 0 8064 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1669390400
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_73
timestamp 1669390400
transform 1 0 9520 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_76
timestamp 1669390400
transform 1 0 9856 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_80
timestamp 1669390400
transform 1 0 10304 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_84
timestamp 1669390400
transform 1 0 10752 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_99
timestamp 1669390400
transform 1 0 12432 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_111
timestamp 1669390400
transform 1 0 13776 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_118
timestamp 1669390400
transform 1 0 14560 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_122
timestamp 1669390400
transform 1 0 15008 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_125
timestamp 1669390400
transform 1 0 15344 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_129
timestamp 1669390400
transform 1 0 15792 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_133
timestamp 1669390400
transform 1 0 16240 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_140
timestamp 1669390400
transform 1 0 17024 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_144
timestamp 1669390400
transform 1 0 17472 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_147
timestamp 1669390400
transform 1 0 17808 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_151
timestamp 1669390400
transform 1 0 18256 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_161
timestamp 1669390400
transform 1 0 19376 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_171
timestamp 1669390400
transform 1 0 20496 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_196
timestamp 1669390400
transform 1 0 23296 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_204
timestamp 1669390400
transform 1 0 24192 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_211
timestamp 1669390400
transform 1 0 24976 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_215
timestamp 1669390400
transform 1 0 25424 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_218
timestamp 1669390400
transform 1 0 25760 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_235
timestamp 1669390400
transform 1 0 27664 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_242
timestamp 1669390400
transform 1 0 28448 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_246
timestamp 1669390400
transform 1 0 28896 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_254
timestamp 1669390400
transform 1 0 29792 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_258
timestamp 1669390400
transform 1 0 30240 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_260
timestamp 1669390400
transform 1 0 30464 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_269
timestamp 1669390400
transform 1 0 31472 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_273
timestamp 1669390400
transform 1 0 31920 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_277
timestamp 1669390400
transform 1 0 32368 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_281
timestamp 1669390400
transform 1 0 32816 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1669390400
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_286
timestamp 1669390400
transform 1 0 33376 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_303
timestamp 1669390400
transform 1 0 35280 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_307
timestamp 1669390400
transform 1 0 35728 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_311
timestamp 1669390400
transform 1 0 36176 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_335
timestamp 1669390400
transform 1 0 38864 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_342
timestamp 1669390400
transform 1 0 39648 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_344
timestamp 1669390400
transform 1 0 39872 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_347
timestamp 1669390400
transform 1 0 40208 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_351
timestamp 1669390400
transform 1 0 40656 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_357
timestamp 1669390400
transform 1 0 41328 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_366
timestamp 1669390400
transform 1 0 42336 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_376
timestamp 1669390400
transform 1 0 43456 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_378
timestamp 1669390400
transform 1 0 43680 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_394
timestamp 1669390400
transform 1 0 45472 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_411
timestamp 1669390400
transform 1 0 47376 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_423
timestamp 1669390400
transform 1 0 48720 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_425
timestamp 1669390400
transform 1 0 48944 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_428
timestamp 1669390400
transform 1 0 49280 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_435
timestamp 1669390400
transform 1 0 50064 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_443
timestamp 1669390400
transform 1 0 50960 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_447
timestamp 1669390400
transform 1 0 51408 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_449
timestamp 1669390400
transform 1 0 51632 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_456
timestamp 1669390400
transform 1 0 52416 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_494
timestamp 1669390400
transform 1 0 56672 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_496
timestamp 1669390400
transform 1 0 56896 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_499
timestamp 1669390400
transform 1 0 57232 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_506
timestamp 1669390400
transform 1 0 58016 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_508
timestamp 1669390400
transform 1 0 58240 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1669390400
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_17
timestamp 1669390400
transform 1 0 3248 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_19
timestamp 1669390400
transform 1 0 3472 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_22
timestamp 1669390400
transform 1 0 3808 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_26
timestamp 1669390400
transform 1 0 4256 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_30
timestamp 1669390400
transform 1 0 4704 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_34
timestamp 1669390400
transform 1 0 5152 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_37
timestamp 1669390400
transform 1 0 5488 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_45
timestamp 1669390400
transform 1 0 6384 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_59
timestamp 1669390400
transform 1 0 7952 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_63
timestamp 1669390400
transform 1 0 8400 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_66
timestamp 1669390400
transform 1 0 8736 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_101
timestamp 1669390400
transform 1 0 12656 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1669390400
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_108
timestamp 1669390400
transform 1 0 13440 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_122
timestamp 1669390400
transform 1 0 15008 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_134
timestamp 1669390400
transform 1 0 16352 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_151
timestamp 1669390400
transform 1 0 18256 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_168
timestamp 1669390400
transform 1 0 20160 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_172
timestamp 1669390400
transform 1 0 20608 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1669390400
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_179
timestamp 1669390400
transform 1 0 21392 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_183
timestamp 1669390400
transform 1 0 21840 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_187
timestamp 1669390400
transform 1 0 22288 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_191
timestamp 1669390400
transform 1 0 22736 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_195
timestamp 1669390400
transform 1 0 23184 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_205
timestamp 1669390400
transform 1 0 24304 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_213
timestamp 1669390400
transform 1 0 25200 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_217
timestamp 1669390400
transform 1 0 25648 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_220
timestamp 1669390400
transform 1 0 25984 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_224
timestamp 1669390400
transform 1 0 26432 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_234
timestamp 1669390400
transform 1 0 27552 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_242
timestamp 1669390400
transform 1 0 28448 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_246
timestamp 1669390400
transform 1 0 28896 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_250
timestamp 1669390400
transform 1 0 29344 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_254
timestamp 1669390400
transform 1 0 29792 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_256
timestamp 1669390400
transform 1 0 30016 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_263
timestamp 1669390400
transform 1 0 30800 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_270
timestamp 1669390400
transform 1 0 31584 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_272
timestamp 1669390400
transform 1 0 31808 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_279
timestamp 1669390400
transform 1 0 32592 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_293
timestamp 1669390400
transform 1 0 34160 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_302
timestamp 1669390400
transform 1 0 35168 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_306
timestamp 1669390400
transform 1 0 35616 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_310
timestamp 1669390400
transform 1 0 36064 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_312
timestamp 1669390400
transform 1 0 36288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1669390400
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_321
timestamp 1669390400
transform 1 0 37296 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_332
timestamp 1669390400
transform 1 0 38528 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_336
timestamp 1669390400
transform 1 0 38976 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_340
timestamp 1669390400
transform 1 0 39424 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_344
timestamp 1669390400
transform 1 0 39872 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_348
timestamp 1669390400
transform 1 0 40320 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1669390400
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_392
timestamp 1669390400
transform 1 0 45248 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_395
timestamp 1669390400
transform 1 0 45584 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_397
timestamp 1669390400
transform 1 0 45808 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_416
timestamp 1669390400
transform 1 0 47936 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_436
timestamp 1669390400
transform 1 0 50176 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_438
timestamp 1669390400
transform 1 0 50400 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_447
timestamp 1669390400
transform 1 0 51408 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_460
timestamp 1669390400
transform 1 0 52864 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_463
timestamp 1669390400
transform 1 0 53200 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_474
timestamp 1669390400
transform 1 0 54432 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_478
timestamp 1669390400
transform 1 0 54880 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_485
timestamp 1669390400
transform 1 0 55664 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_495
timestamp 1669390400
transform 1 0 56784 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_505
timestamp 1669390400
transform 1 0 57904 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_2
timestamp 1669390400
transform 1 0 1568 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_8
timestamp 1669390400
transform 1 0 2240 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_12
timestamp 1669390400
transform 1 0 2688 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_16
timestamp 1669390400
transform 1 0 3136 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_20
timestamp 1669390400
transform 1 0 3584 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_24
timestamp 1669390400
transform 1 0 4032 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_28
timestamp 1669390400
transform 1 0 4480 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_32
timestamp 1669390400
transform 1 0 4928 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_42
timestamp 1669390400
transform 1 0 6048 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_48
timestamp 1669390400
transform 1 0 6720 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_57
timestamp 1669390400
transform 1 0 7728 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_61
timestamp 1669390400
transform 1 0 8176 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1669390400
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_73
timestamp 1669390400
transform 1 0 9520 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_75
timestamp 1669390400
transform 1 0 9744 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_78
timestamp 1669390400
transform 1 0 10080 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_88
timestamp 1669390400
transform 1 0 11200 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_130
timestamp 1669390400
transform 1 0 15904 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_140
timestamp 1669390400
transform 1 0 17024 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_144
timestamp 1669390400
transform 1 0 17472 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_156
timestamp 1669390400
transform 1 0 18816 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_158
timestamp 1669390400
transform 1 0 19040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_161
timestamp 1669390400
transform 1 0 19376 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_165
timestamp 1669390400
transform 1 0 19824 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_173
timestamp 1669390400
transform 1 0 20720 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_177
timestamp 1669390400
transform 1 0 21168 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_181
timestamp 1669390400
transform 1 0 21616 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_185
timestamp 1669390400
transform 1 0 22064 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_193
timestamp 1669390400
transform 1 0 22960 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1669390400
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_215
timestamp 1669390400
transform 1 0 25424 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_224
timestamp 1669390400
transform 1 0 26432 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_228
timestamp 1669390400
transform 1 0 26880 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_236
timestamp 1669390400
transform 1 0 27776 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_240
timestamp 1669390400
transform 1 0 28224 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_254
timestamp 1669390400
transform 1 0 29792 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_269
timestamp 1669390400
transform 1 0 31472 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_273
timestamp 1669390400
transform 1 0 31920 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1669390400
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_286
timestamp 1669390400
transform 1 0 33376 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_289
timestamp 1669390400
transform 1 0 33712 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_291
timestamp 1669390400
transform 1 0 33936 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_300
timestamp 1669390400
transform 1 0 34944 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_304
timestamp 1669390400
transform 1 0 35392 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_323
timestamp 1669390400
transform 1 0 37520 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_333
timestamp 1669390400
transform 1 0 38640 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_343
timestamp 1669390400
transform 1 0 39760 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_353
timestamp 1669390400
transform 1 0 40880 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_357
timestamp 1669390400
transform 1 0 41328 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_364
timestamp 1669390400
transform 1 0 42112 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_368
timestamp 1669390400
transform 1 0 42560 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_412
timestamp 1669390400
transform 1 0 47488 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_419
timestamp 1669390400
transform 1 0 48272 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_425
timestamp 1669390400
transform 1 0 48944 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_428
timestamp 1669390400
transform 1 0 49280 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_430
timestamp 1669390400
transform 1 0 49504 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_437
timestamp 1669390400
transform 1 0 50288 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_449
timestamp 1669390400
transform 1 0 51632 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_451
timestamp 1669390400
transform 1 0 51856 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_470
timestamp 1669390400
transform 1 0 53984 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_474
timestamp 1669390400
transform 1 0 54432 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_486
timestamp 1669390400
transform 1 0 55776 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_496
timestamp 1669390400
transform 1 0 56896 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_499
timestamp 1669390400
transform 1 0 57232 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_506
timestamp 1669390400
transform 1 0 58016 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_508
timestamp 1669390400
transform 1 0 58240 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_2
timestamp 1669390400
transform 1 0 1568 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_6
timestamp 1669390400
transform 1 0 2016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_10
timestamp 1669390400
transform 1 0 2464 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_14
timestamp 1669390400
transform 1 0 2912 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_18
timestamp 1669390400
transform 1 0 3360 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_22
timestamp 1669390400
transform 1 0 3808 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_26
timestamp 1669390400
transform 1 0 4256 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_30
timestamp 1669390400
transform 1 0 4704 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_34
timestamp 1669390400
transform 1 0 5152 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_37
timestamp 1669390400
transform 1 0 5488 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_50
timestamp 1669390400
transform 1 0 6944 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_54
timestamp 1669390400
transform 1 0 7392 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_57
timestamp 1669390400
transform 1 0 7728 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_67
timestamp 1669390400
transform 1 0 8848 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_71
timestamp 1669390400
transform 1 0 9296 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_75
timestamp 1669390400
transform 1 0 9744 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_79
timestamp 1669390400
transform 1 0 10192 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_83
timestamp 1669390400
transform 1 0 10640 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_90
timestamp 1669390400
transform 1 0 11424 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_94
timestamp 1669390400
transform 1 0 11872 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_96
timestamp 1669390400
transform 1 0 12096 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1669390400
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_108
timestamp 1669390400
transform 1 0 13440 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_120
timestamp 1669390400
transform 1 0 14784 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_130
timestamp 1669390400
transform 1 0 15904 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_134
timestamp 1669390400
transform 1 0 16352 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_136
timestamp 1669390400
transform 1 0 16576 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_139
timestamp 1669390400
transform 1 0 16912 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_149
timestamp 1669390400
transform 1 0 18032 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_157
timestamp 1669390400
transform 1 0 18928 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_161
timestamp 1669390400
transform 1 0 19376 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_168
timestamp 1669390400
transform 1 0 20160 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1669390400
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_179
timestamp 1669390400
transform 1 0 21392 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_187
timestamp 1669390400
transform 1 0 22288 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_210
timestamp 1669390400
transform 1 0 24864 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_216
timestamp 1669390400
transform 1 0 25536 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_220
timestamp 1669390400
transform 1 0 25984 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_224
timestamp 1669390400
transform 1 0 26432 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_232
timestamp 1669390400
transform 1 0 27328 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_236
timestamp 1669390400
transform 1 0 27776 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_240
timestamp 1669390400
transform 1 0 28224 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_247
timestamp 1669390400
transform 1 0 29008 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_250
timestamp 1669390400
transform 1 0 29344 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_256
timestamp 1669390400
transform 1 0 30016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_266
timestamp 1669390400
transform 1 0 31136 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_274
timestamp 1669390400
transform 1 0 32032 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_278
timestamp 1669390400
transform 1 0 32480 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_280
timestamp 1669390400
transform 1 0 32704 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1669390400
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_321
timestamp 1669390400
transform 1 0 37296 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_328
timestamp 1669390400
transform 1 0 38080 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_354
timestamp 1669390400
transform 1 0 40992 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_358
timestamp 1669390400
transform 1 0 41440 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_370
timestamp 1669390400
transform 1 0 42784 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_374
timestamp 1669390400
transform 1 0 43232 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_378
timestamp 1669390400
transform 1 0 43680 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_388
timestamp 1669390400
transform 1 0 44800 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_392
timestamp 1669390400
transform 1 0 45248 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_398
timestamp 1669390400
transform 1 0 45920 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_402
timestamp 1669390400
transform 1 0 46368 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_406
timestamp 1669390400
transform 1 0 46816 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_434
timestamp 1669390400
transform 1 0 49952 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_438
timestamp 1669390400
transform 1 0 50400 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_440
timestamp 1669390400
transform 1 0 50624 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_460
timestamp 1669390400
transform 1 0 52864 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_463
timestamp 1669390400
transform 1 0 53200 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_466
timestamp 1669390400
transform 1 0 53536 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_470
timestamp 1669390400
transform 1 0 53984 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_474
timestamp 1669390400
transform 1 0 54432 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_478
timestamp 1669390400
transform 1 0 54880 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_482
timestamp 1669390400
transform 1 0 55328 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_486
timestamp 1669390400
transform 1 0 55776 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_488
timestamp 1669390400
transform 1 0 56000 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_502
timestamp 1669390400
transform 1 0 57568 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_506
timestamp 1669390400
transform 1 0 58016 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_508
timestamp 1669390400
transform 1 0 58240 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_2
timestamp 1669390400
transform 1 0 1568 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_6
timestamp 1669390400
transform 1 0 2016 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_10
timestamp 1669390400
transform 1 0 2464 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_14
timestamp 1669390400
transform 1 0 2912 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_18
timestamp 1669390400
transform 1 0 3360 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_22
timestamp 1669390400
transform 1 0 3808 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_26
timestamp 1669390400
transform 1 0 4256 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_30
timestamp 1669390400
transform 1 0 4704 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_38
timestamp 1669390400
transform 1 0 5600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_42
timestamp 1669390400
transform 1 0 6048 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_45
timestamp 1669390400
transform 1 0 6384 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_49
timestamp 1669390400
transform 1 0 6832 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_53
timestamp 1669390400
transform 1 0 7280 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_57
timestamp 1669390400
transform 1 0 7728 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_69
timestamp 1669390400
transform 1 0 9072 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_73
timestamp 1669390400
transform 1 0 9520 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_76
timestamp 1669390400
transform 1 0 9856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_80
timestamp 1669390400
transform 1 0 10304 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_83
timestamp 1669390400
transform 1 0 10640 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_87
timestamp 1669390400
transform 1 0 11088 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_91
timestamp 1669390400
transform 1 0 11536 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_99
timestamp 1669390400
transform 1 0 12432 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_103
timestamp 1669390400
transform 1 0 12880 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_107
timestamp 1669390400
transform 1 0 13328 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_113
timestamp 1669390400
transform 1 0 14000 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_117
timestamp 1669390400
transform 1 0 14448 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_121
timestamp 1669390400
transform 1 0 14896 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_125
timestamp 1669390400
transform 1 0 15344 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_129
timestamp 1669390400
transform 1 0 15792 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_132
timestamp 1669390400
transform 1 0 16128 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_134
timestamp 1669390400
transform 1 0 16352 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_137
timestamp 1669390400
transform 1 0 16688 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1669390400
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_144
timestamp 1669390400
transform 1 0 17472 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_147
timestamp 1669390400
transform 1 0 17808 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_153
timestamp 1669390400
transform 1 0 18480 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_157
timestamp 1669390400
transform 1 0 18928 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_159
timestamp 1669390400
transform 1 0 19152 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_184
timestamp 1669390400
transform 1 0 21952 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_194
timestamp 1669390400
transform 1 0 23072 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_198
timestamp 1669390400
transform 1 0 23520 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_201
timestamp 1669390400
transform 1 0 23856 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_205
timestamp 1669390400
transform 1 0 24304 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_212
timestamp 1669390400
transform 1 0 25088 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_215
timestamp 1669390400
transform 1 0 25424 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_224
timestamp 1669390400
transform 1 0 26432 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_237
timestamp 1669390400
transform 1 0 27888 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_241
timestamp 1669390400
transform 1 0 28336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_245
timestamp 1669390400
transform 1 0 28784 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_247
timestamp 1669390400
transform 1 0 29008 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_261
timestamp 1669390400
transform 1 0 30576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_271
timestamp 1669390400
transform 1 0 31696 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_275
timestamp 1669390400
transform 1 0 32144 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_283
timestamp 1669390400
transform 1 0 33040 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_286
timestamp 1669390400
transform 1 0 33376 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_298
timestamp 1669390400
transform 1 0 34720 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_302
timestamp 1669390400
transform 1 0 35168 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_304
timestamp 1669390400
transform 1 0 35392 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_345
timestamp 1669390400
transform 1 0 39984 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1669390400
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_357
timestamp 1669390400
transform 1 0 41328 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_360
timestamp 1669390400
transform 1 0 41664 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_362
timestamp 1669390400
transform 1 0 41888 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_375
timestamp 1669390400
transform 1 0 43344 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_385
timestamp 1669390400
transform 1 0 44464 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_395
timestamp 1669390400
transform 1 0 45584 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_399
timestamp 1669390400
transform 1 0 46032 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_403
timestamp 1669390400
transform 1 0 46480 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_425
timestamp 1669390400
transform 1 0 48944 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_428
timestamp 1669390400
transform 1 0 49280 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_436
timestamp 1669390400
transform 1 0 50176 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_445
timestamp 1669390400
transform 1 0 51184 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_487
timestamp 1669390400
transform 1 0 55888 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_489
timestamp 1669390400
transform 1 0 56112 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_496
timestamp 1669390400
transform 1 0 56896 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_499
timestamp 1669390400
transform 1 0 57232 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_506
timestamp 1669390400
transform 1 0 58016 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_508
timestamp 1669390400
transform 1 0 58240 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_2
timestamp 1669390400
transform 1 0 1568 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_6
timestamp 1669390400
transform 1 0 2016 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_10
timestamp 1669390400
transform 1 0 2464 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_14
timestamp 1669390400
transform 1 0 2912 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_18
timestamp 1669390400
transform 1 0 3360 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_22
timestamp 1669390400
transform 1 0 3808 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_26
timestamp 1669390400
transform 1 0 4256 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_30
timestamp 1669390400
transform 1 0 4704 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1669390400
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_37
timestamp 1669390400
transform 1 0 5488 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_40
timestamp 1669390400
transform 1 0 5824 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_44
timestamp 1669390400
transform 1 0 6272 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_48
timestamp 1669390400
transform 1 0 6720 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_52
timestamp 1669390400
transform 1 0 7168 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_73
timestamp 1669390400
transform 1 0 9520 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_83
timestamp 1669390400
transform 1 0 10640 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_87
timestamp 1669390400
transform 1 0 11088 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_101
timestamp 1669390400
transform 1 0 12656 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1669390400
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_108
timestamp 1669390400
transform 1 0 13440 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_119
timestamp 1669390400
transform 1 0 14672 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_135
timestamp 1669390400
transform 1 0 16464 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_137
timestamp 1669390400
transform 1 0 16688 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_164
timestamp 1669390400
transform 1 0 19712 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_172
timestamp 1669390400
transform 1 0 20608 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1669390400
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_179
timestamp 1669390400
transform 1 0 21392 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_188
timestamp 1669390400
transform 1 0 22400 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_192
timestamp 1669390400
transform 1 0 22848 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_203
timestamp 1669390400
transform 1 0 24080 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_211
timestamp 1669390400
transform 1 0 24976 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_241
timestamp 1669390400
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_245
timestamp 1669390400
transform 1 0 28784 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_247
timestamp 1669390400
transform 1 0 29008 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_250
timestamp 1669390400
transform 1 0 29344 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_258
timestamp 1669390400
transform 1 0 30240 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_260
timestamp 1669390400
transform 1 0 30464 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_263
timestamp 1669390400
transform 1 0 30800 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_265
timestamp 1669390400
transform 1 0 31024 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_36_270
timestamp 1669390400
transform 1 0 31584 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_278
timestamp 1669390400
transform 1 0 32480 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_282
timestamp 1669390400
transform 1 0 32928 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_296
timestamp 1669390400
transform 1 0 34496 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_300
timestamp 1669390400
transform 1 0 34944 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_302
timestamp 1669390400
transform 1 0 35168 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_308
timestamp 1669390400
transform 1 0 35840 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1669390400
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_321
timestamp 1669390400
transform 1 0 37296 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_330
timestamp 1669390400
transform 1 0 38304 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_334
timestamp 1669390400
transform 1 0 38752 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_336
timestamp 1669390400
transform 1 0 38976 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_345
timestamp 1669390400
transform 1 0 39984 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_355
timestamp 1669390400
transform 1 0 41104 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_365
timestamp 1669390400
transform 1 0 42224 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_375
timestamp 1669390400
transform 1 0 43344 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_379
timestamp 1669390400
transform 1 0 43792 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1669390400
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_392
timestamp 1669390400
transform 1 0 45248 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_408
timestamp 1669390400
transform 1 0 47040 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_425
timestamp 1669390400
transform 1 0 48944 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_440
timestamp 1669390400
transform 1 0 50624 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_448
timestamp 1669390400
transform 1 0 51520 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_460
timestamp 1669390400
transform 1 0 52864 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_463
timestamp 1669390400
transform 1 0 53200 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_470
timestamp 1669390400
transform 1 0 53984 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_486
timestamp 1669390400
transform 1 0 55776 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_497
timestamp 1669390400
transform 1 0 57008 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_507
timestamp 1669390400
transform 1 0 58128 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_2
timestamp 1669390400
transform 1 0 1568 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_10
timestamp 1669390400
transform 1 0 2464 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_14
timestamp 1669390400
transform 1 0 2912 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_16
timestamp 1669390400
transform 1 0 3136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_19
timestamp 1669390400
transform 1 0 3472 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_23
timestamp 1669390400
transform 1 0 3920 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_27
timestamp 1669390400
transform 1 0 4368 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_40
timestamp 1669390400
transform 1 0 5824 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_48
timestamp 1669390400
transform 1 0 6720 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_52
timestamp 1669390400
transform 1 0 7168 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_60
timestamp 1669390400
transform 1 0 8064 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1669390400
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_73
timestamp 1669390400
transform 1 0 9520 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_76
timestamp 1669390400
transform 1 0 9856 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_80
timestamp 1669390400
transform 1 0 10304 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_86
timestamp 1669390400
transform 1 0 10976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_90
timestamp 1669390400
transform 1 0 11424 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_104
timestamp 1669390400
transform 1 0 12992 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_114
timestamp 1669390400
transform 1 0 14112 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_118
timestamp 1669390400
transform 1 0 14560 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_125
timestamp 1669390400
transform 1 0 15344 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_140
timestamp 1669390400
transform 1 0 17024 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_144
timestamp 1669390400
transform 1 0 17472 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_151
timestamp 1669390400
transform 1 0 18256 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_166
timestamp 1669390400
transform 1 0 19936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_174
timestamp 1669390400
transform 1 0 20832 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_176
timestamp 1669390400
transform 1 0 21056 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_179
timestamp 1669390400
transform 1 0 21392 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_186
timestamp 1669390400
transform 1 0 22176 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_193
timestamp 1669390400
transform 1 0 22960 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_207
timestamp 1669390400
transform 1 0 24528 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_211
timestamp 1669390400
transform 1 0 24976 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_215
timestamp 1669390400
transform 1 0 25424 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_217
timestamp 1669390400
transform 1 0 25648 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_223
timestamp 1669390400
transform 1 0 26320 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_233
timestamp 1669390400
transform 1 0 27440 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_237
timestamp 1669390400
transform 1 0 27888 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_241
timestamp 1669390400
transform 1 0 28336 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_257
timestamp 1669390400
transform 1 0 30128 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_259
timestamp 1669390400
transform 1 0 30352 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_262
timestamp 1669390400
transform 1 0 30688 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_266
timestamp 1669390400
transform 1 0 31136 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_274
timestamp 1669390400
transform 1 0 32032 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_278
timestamp 1669390400
transform 1 0 32480 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_280
timestamp 1669390400
transform 1 0 32704 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_283
timestamp 1669390400
transform 1 0 33040 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_286
timestamp 1669390400
transform 1 0 33376 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_294
timestamp 1669390400
transform 1 0 34272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_298
timestamp 1669390400
transform 1 0 34720 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_301
timestamp 1669390400
transform 1 0 35056 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_326
timestamp 1669390400
transform 1 0 37856 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_330
timestamp 1669390400
transform 1 0 38304 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_334
timestamp 1669390400
transform 1 0 38752 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_346
timestamp 1669390400
transform 1 0 40096 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_350
timestamp 1669390400
transform 1 0 40544 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1669390400
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_357
timestamp 1669390400
transform 1 0 41328 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_366
timestamp 1669390400
transform 1 0 42336 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_370
timestamp 1669390400
transform 1 0 42784 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_374
timestamp 1669390400
transform 1 0 43232 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_385
timestamp 1669390400
transform 1 0 44464 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_395
timestamp 1669390400
transform 1 0 45584 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_405
timestamp 1669390400
transform 1 0 46704 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_412
timestamp 1669390400
transform 1 0 47488 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_422
timestamp 1669390400
transform 1 0 48608 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_428
timestamp 1669390400
transform 1 0 49280 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_438
timestamp 1669390400
transform 1 0 50400 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_446
timestamp 1669390400
transform 1 0 51296 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_450
timestamp 1669390400
transform 1 0 51744 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_462
timestamp 1669390400
transform 1 0 53088 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_475
timestamp 1669390400
transform 1 0 54544 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_491
timestamp 1669390400
transform 1 0 56336 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_495
timestamp 1669390400
transform 1 0 56784 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_499
timestamp 1669390400
transform 1 0 57232 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_506
timestamp 1669390400
transform 1 0 58016 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_508
timestamp 1669390400
transform 1 0 58240 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_2
timestamp 1669390400
transform 1 0 1568 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_18
timestamp 1669390400
transform 1 0 3360 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_20
timestamp 1669390400
transform 1 0 3584 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1669390400
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_37
timestamp 1669390400
transform 1 0 5488 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_56
timestamp 1669390400
transform 1 0 7616 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_68
timestamp 1669390400
transform 1 0 8960 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_72
timestamp 1669390400
transform 1 0 9408 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_76
timestamp 1669390400
transform 1 0 9856 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_92
timestamp 1669390400
transform 1 0 11648 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_101
timestamp 1669390400
transform 1 0 12656 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1669390400
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_108
timestamp 1669390400
transform 1 0 13440 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_115
timestamp 1669390400
transform 1 0 14224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_119
timestamp 1669390400
transform 1 0 14672 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_121
timestamp 1669390400
transform 1 0 14896 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_124
timestamp 1669390400
transform 1 0 15232 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_128
timestamp 1669390400
transform 1 0 15680 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_130
timestamp 1669390400
transform 1 0 15904 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_139
timestamp 1669390400
transform 1 0 16912 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_143
timestamp 1669390400
transform 1 0 17360 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_147
timestamp 1669390400
transform 1 0 17808 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_155
timestamp 1669390400
transform 1 0 18704 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_161
timestamp 1669390400
transform 1 0 19376 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_163
timestamp 1669390400
transform 1 0 19600 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_166
timestamp 1669390400
transform 1 0 19936 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1669390400
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_179
timestamp 1669390400
transform 1 0 21392 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_183
timestamp 1669390400
transform 1 0 21840 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_187
timestamp 1669390400
transform 1 0 22288 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_202
timestamp 1669390400
transform 1 0 23968 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_229
timestamp 1669390400
transform 1 0 26992 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_239
timestamp 1669390400
transform 1 0 28112 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_247
timestamp 1669390400
transform 1 0 29008 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_250
timestamp 1669390400
transform 1 0 29344 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_260
timestamp 1669390400
transform 1 0 30464 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_268
timestamp 1669390400
transform 1 0 31360 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_272
timestamp 1669390400
transform 1 0 31808 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_281
timestamp 1669390400
transform 1 0 32816 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_295
timestamp 1669390400
transform 1 0 34384 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_299
timestamp 1669390400
transform 1 0 34832 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_305
timestamp 1669390400
transform 1 0 35504 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_307
timestamp 1669390400
transform 1 0 35728 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_314
timestamp 1669390400
transform 1 0 36512 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_318
timestamp 1669390400
transform 1 0 36960 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_321
timestamp 1669390400
transform 1 0 37296 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_324
timestamp 1669390400
transform 1 0 37632 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_328
timestamp 1669390400
transform 1 0 38080 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_332
timestamp 1669390400
transform 1 0 38528 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_336
timestamp 1669390400
transform 1 0 38976 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_347
timestamp 1669390400
transform 1 0 40208 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_351
timestamp 1669390400
transform 1 0 40656 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_355
timestamp 1669390400
transform 1 0 41104 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_357
timestamp 1669390400
transform 1 0 41328 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_368
timestamp 1669390400
transform 1 0 42560 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_372
timestamp 1669390400
transform 1 0 43008 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_376
timestamp 1669390400
transform 1 0 43456 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_380
timestamp 1669390400
transform 1 0 43904 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_384
timestamp 1669390400
transform 1 0 44352 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_388
timestamp 1669390400
transform 1 0 44800 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_392
timestamp 1669390400
transform 1 0 45248 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_399
timestamp 1669390400
transform 1 0 46032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_403
timestamp 1669390400
transform 1 0 46480 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_407
timestamp 1669390400
transform 1 0 46928 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_411
timestamp 1669390400
transform 1 0 47376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_428
timestamp 1669390400
transform 1 0 49280 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_432
timestamp 1669390400
transform 1 0 49728 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_444
timestamp 1669390400
transform 1 0 51072 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_452
timestamp 1669390400
transform 1 0 51968 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_460
timestamp 1669390400
transform 1 0 52864 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_463
timestamp 1669390400
transform 1 0 53200 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_466
timestamp 1669390400
transform 1 0 53536 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_468
timestamp 1669390400
transform 1 0 53760 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_483
timestamp 1669390400
transform 1 0 55440 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_493
timestamp 1669390400
transform 1 0 56560 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_503
timestamp 1669390400
transform 1 0 57680 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_507
timestamp 1669390400
transform 1 0 58128 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_2
timestamp 1669390400
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_18
timestamp 1669390400
transform 1 0 3360 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_26
timestamp 1669390400
transform 1 0 4256 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_30
timestamp 1669390400
transform 1 0 4704 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_34
timestamp 1669390400
transform 1 0 5152 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_38
timestamp 1669390400
transform 1 0 5600 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_47
timestamp 1669390400
transform 1 0 6608 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_55
timestamp 1669390400
transform 1 0 7504 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_61
timestamp 1669390400
transform 1 0 8176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_65
timestamp 1669390400
transform 1 0 8624 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_67
timestamp 1669390400
transform 1 0 8848 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1669390400
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_73
timestamp 1669390400
transform 1 0 9520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_84
timestamp 1669390400
transform 1 0 10752 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_91
timestamp 1669390400
transform 1 0 11536 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_99
timestamp 1669390400
transform 1 0 12432 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_101
timestamp 1669390400
transform 1 0 12656 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_104
timestamp 1669390400
transform 1 0 12992 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_108
timestamp 1669390400
transform 1 0 13440 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_116
timestamp 1669390400
transform 1 0 14336 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_120
timestamp 1669390400
transform 1 0 14784 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_124
timestamp 1669390400
transform 1 0 15232 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_130
timestamp 1669390400
transform 1 0 15904 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_138
timestamp 1669390400
transform 1 0 16800 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_144
timestamp 1669390400
transform 1 0 17472 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_146
timestamp 1669390400
transform 1 0 17696 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_159
timestamp 1669390400
transform 1 0 19152 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_174
timestamp 1669390400
transform 1 0 20832 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_176
timestamp 1669390400
transform 1 0 21056 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_211
timestamp 1669390400
transform 1 0 24976 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_215
timestamp 1669390400
transform 1 0 25424 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_227
timestamp 1669390400
transform 1 0 26768 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_231
timestamp 1669390400
transform 1 0 27216 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_239
timestamp 1669390400
transform 1 0 28112 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_247
timestamp 1669390400
transform 1 0 29008 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_249
timestamp 1669390400
transform 1 0 29232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_252
timestamp 1669390400
transform 1 0 29568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_259
timestamp 1669390400
transform 1 0 30352 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_269
timestamp 1669390400
transform 1 0 31472 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_273
timestamp 1669390400
transform 1 0 31920 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_281
timestamp 1669390400
transform 1 0 32816 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_283
timestamp 1669390400
transform 1 0 33040 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_286
timestamp 1669390400
transform 1 0 33376 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_299
timestamp 1669390400
transform 1 0 34832 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_303
timestamp 1669390400
transform 1 0 35280 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_305
timestamp 1669390400
transform 1 0 35504 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_314
timestamp 1669390400
transform 1 0 36512 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_333
timestamp 1669390400
transform 1 0 38640 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_337
timestamp 1669390400
transform 1 0 39088 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1669390400
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_357
timestamp 1669390400
transform 1 0 41328 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_373
timestamp 1669390400
transform 1 0 43120 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_375
timestamp 1669390400
transform 1 0 43344 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_399
timestamp 1669390400
transform 1 0 46032 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_407
timestamp 1669390400
transform 1 0 46928 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_415
timestamp 1669390400
transform 1 0 47824 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_419
timestamp 1669390400
transform 1 0 48272 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_423
timestamp 1669390400
transform 1 0 48720 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_425
timestamp 1669390400
transform 1 0 48944 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_428
timestamp 1669390400
transform 1 0 49280 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_438
timestamp 1669390400
transform 1 0 50400 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_442
timestamp 1669390400
transform 1 0 50848 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_444
timestamp 1669390400
transform 1 0 51072 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_453
timestamp 1669390400
transform 1 0 52080 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_461
timestamp 1669390400
transform 1 0 52976 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_470
timestamp 1669390400
transform 1 0 53984 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_480
timestamp 1669390400
transform 1 0 55104 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_487
timestamp 1669390400
transform 1 0 55888 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_489
timestamp 1669390400
transform 1 0 56112 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_496
timestamp 1669390400
transform 1 0 56896 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_499
timestamp 1669390400
transform 1 0 57232 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_504
timestamp 1669390400
transform 1 0 57792 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_508
timestamp 1669390400
transform 1 0 58240 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_2
timestamp 1669390400
transform 1 0 1568 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_17
timestamp 1669390400
transform 1 0 3248 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_21
timestamp 1669390400
transform 1 0 3696 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_25
timestamp 1669390400
transform 1 0 4144 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1669390400
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_37
timestamp 1669390400
transform 1 0 5488 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_49
timestamp 1669390400
transform 1 0 6832 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_51
timestamp 1669390400
transform 1 0 7056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_54
timestamp 1669390400
transform 1 0 7392 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_67
timestamp 1669390400
transform 1 0 8848 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_71
timestamp 1669390400
transform 1 0 9296 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_75
timestamp 1669390400
transform 1 0 9744 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_85
timestamp 1669390400
transform 1 0 10864 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_99
timestamp 1669390400
transform 1 0 12432 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1669390400
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_108
timestamp 1669390400
transform 1 0 13440 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_122
timestamp 1669390400
transform 1 0 15008 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_134
timestamp 1669390400
transform 1 0 16352 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_138
timestamp 1669390400
transform 1 0 16800 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_158
timestamp 1669390400
transform 1 0 19040 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_162
timestamp 1669390400
transform 1 0 19488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1669390400
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1669390400
transform 1 0 21392 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_186
timestamp 1669390400
transform 1 0 22176 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_190
timestamp 1669390400
transform 1 0 22624 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_194
timestamp 1669390400
transform 1 0 23072 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_197
timestamp 1669390400
transform 1 0 23408 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_203
timestamp 1669390400
transform 1 0 24080 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_239
timestamp 1669390400
transform 1 0 28112 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_243
timestamp 1669390400
transform 1 0 28560 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1669390400
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1669390400
transform 1 0 29344 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_273
timestamp 1669390400
transform 1 0 31920 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_280
timestamp 1669390400
transform 1 0 32704 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_284
timestamp 1669390400
transform 1 0 33152 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_286
timestamp 1669390400
transform 1 0 33376 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_292
timestamp 1669390400
transform 1 0 34048 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_296
timestamp 1669390400
transform 1 0 34496 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_304
timestamp 1669390400
transform 1 0 35392 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_307
timestamp 1669390400
transform 1 0 35728 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_315
timestamp 1669390400
transform 1 0 36624 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_321
timestamp 1669390400
transform 1 0 37296 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_328
timestamp 1669390400
transform 1 0 38080 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_330
timestamp 1669390400
transform 1 0 38304 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_340
timestamp 1669390400
transform 1 0 39424 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_377
timestamp 1669390400
transform 1 0 43568 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_381
timestamp 1669390400
transform 1 0 44016 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_385
timestamp 1669390400
transform 1 0 44464 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1669390400
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_392
timestamp 1669390400
transform 1 0 45248 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_395
timestamp 1669390400
transform 1 0 45584 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_397
timestamp 1669390400
transform 1 0 45808 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_404
timestamp 1669390400
transform 1 0 46592 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_408
timestamp 1669390400
transform 1 0 47040 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_412
timestamp 1669390400
transform 1 0 47488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_416
timestamp 1669390400
transform 1 0 47936 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_454
timestamp 1669390400
transform 1 0 52192 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_458
timestamp 1669390400
transform 1 0 52640 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_460
timestamp 1669390400
transform 1 0 52864 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_463
timestamp 1669390400
transform 1 0 53200 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_470
timestamp 1669390400
transform 1 0 53984 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_478
timestamp 1669390400
transform 1 0 54880 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_480
timestamp 1669390400
transform 1 0 55104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_487
timestamp 1669390400
transform 1 0 55888 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_491
timestamp 1669390400
transform 1 0 56336 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_504
timestamp 1669390400
transform 1 0 57792 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_508
timestamp 1669390400
transform 1 0 58240 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_2
timestamp 1669390400
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_18
timestamp 1669390400
transform 1 0 3360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_38
timestamp 1669390400
transform 1 0 5600 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_44
timestamp 1669390400
transform 1 0 6272 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_54
timestamp 1669390400
transform 1 0 7392 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_56
timestamp 1669390400
transform 1 0 7616 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_59
timestamp 1669390400
transform 1 0 7952 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_63
timestamp 1669390400
transform 1 0 8400 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1669390400
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_73
timestamp 1669390400
transform 1 0 9520 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_85
timestamp 1669390400
transform 1 0 10864 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_91
timestamp 1669390400
transform 1 0 11536 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_95
timestamp 1669390400
transform 1 0 11984 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_97
timestamp 1669390400
transform 1 0 12208 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_100
timestamp 1669390400
transform 1 0 12544 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_108
timestamp 1669390400
transform 1 0 13440 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_127
timestamp 1669390400
transform 1 0 15568 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_133
timestamp 1669390400
transform 1 0 16240 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1669390400
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1669390400
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_151
timestamp 1669390400
transform 1 0 18256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_155
timestamp 1669390400
transform 1 0 18704 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_158
timestamp 1669390400
transform 1 0 19040 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_162
timestamp 1669390400
transform 1 0 19488 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_172
timestamp 1669390400
transform 1 0 20608 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_176
timestamp 1669390400
transform 1 0 21056 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_180
timestamp 1669390400
transform 1 0 21504 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_184
timestamp 1669390400
transform 1 0 21952 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_200
timestamp 1669390400
transform 1 0 23744 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_210
timestamp 1669390400
transform 1 0 24864 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1669390400
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_215
timestamp 1669390400
transform 1 0 25424 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_218
timestamp 1669390400
transform 1 0 25760 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_222
timestamp 1669390400
transform 1 0 26208 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_254
timestamp 1669390400
transform 1 0 29792 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_264
timestamp 1669390400
transform 1 0 30912 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_274
timestamp 1669390400
transform 1 0 32032 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_278
timestamp 1669390400
transform 1 0 32480 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_282
timestamp 1669390400
transform 1 0 32928 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_286
timestamp 1669390400
transform 1 0 33376 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_294
timestamp 1669390400
transform 1 0 34272 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_300
timestamp 1669390400
transform 1 0 34944 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_308
timestamp 1669390400
transform 1 0 35840 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_310
timestamp 1669390400
transform 1 0 36064 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_316
timestamp 1669390400
transform 1 0 36736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_320
timestamp 1669390400
transform 1 0 37184 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_324
timestamp 1669390400
transform 1 0 37632 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_337
timestamp 1669390400
transform 1 0 39088 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_354
timestamp 1669390400
transform 1 0 40992 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_357
timestamp 1669390400
transform 1 0 41328 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_360
timestamp 1669390400
transform 1 0 41664 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_364
timestamp 1669390400
transform 1 0 42112 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_384
timestamp 1669390400
transform 1 0 44352 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_388
timestamp 1669390400
transform 1 0 44800 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_398
timestamp 1669390400
transform 1 0 45920 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_408
timestamp 1669390400
transform 1 0 47040 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_412
timestamp 1669390400
transform 1 0 47488 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_415
timestamp 1669390400
transform 1 0 47824 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_425
timestamp 1669390400
transform 1 0 48944 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_428
timestamp 1669390400
transform 1 0 49280 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_431
timestamp 1669390400
transform 1 0 49616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_435
timestamp 1669390400
transform 1 0 50064 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_446
timestamp 1669390400
transform 1 0 51296 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_455
timestamp 1669390400
transform 1 0 52304 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_463
timestamp 1669390400
transform 1 0 53200 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_465
timestamp 1669390400
transform 1 0 53424 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_491
timestamp 1669390400
transform 1 0 56336 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_495
timestamp 1669390400
transform 1 0 56784 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_499
timestamp 1669390400
transform 1 0 57232 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_508
timestamp 1669390400
transform 1 0 58240 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_2
timestamp 1669390400
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_18
timestamp 1669390400
transform 1 0 3360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_26
timestamp 1669390400
transform 1 0 4256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_30
timestamp 1669390400
transform 1 0 4704 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1669390400
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_37
timestamp 1669390400
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_43
timestamp 1669390400
transform 1 0 6160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_47
timestamp 1669390400
transform 1 0 6608 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_51
timestamp 1669390400
transform 1 0 7056 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_55
timestamp 1669390400
transform 1 0 7504 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_69
timestamp 1669390400
transform 1 0 9072 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_77
timestamp 1669390400
transform 1 0 9968 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_81
timestamp 1669390400
transform 1 0 10416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_87
timestamp 1669390400
transform 1 0 11088 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_97
timestamp 1669390400
transform 1 0 12208 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_101
timestamp 1669390400
transform 1 0 12656 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1669390400
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_108
timestamp 1669390400
transform 1 0 13440 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_110
timestamp 1669390400
transform 1 0 13664 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_113
timestamp 1669390400
transform 1 0 14000 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_125
timestamp 1669390400
transform 1 0 15344 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_129
timestamp 1669390400
transform 1 0 15792 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_131
timestamp 1669390400
transform 1 0 16016 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_134
timestamp 1669390400
transform 1 0 16352 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_138
timestamp 1669390400
transform 1 0 16800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_144
timestamp 1669390400
transform 1 0 17472 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_148
timestamp 1669390400
transform 1 0 17920 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_152
timestamp 1669390400
transform 1 0 18368 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_156
timestamp 1669390400
transform 1 0 18816 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_160
timestamp 1669390400
transform 1 0 19264 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_172
timestamp 1669390400
transform 1 0 20608 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1669390400
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1669390400
transform 1 0 21392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_42_186
timestamp 1669390400
transform 1 0 22176 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_194
timestamp 1669390400
transform 1 0 23072 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_198
timestamp 1669390400
transform 1 0 23520 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_202
timestamp 1669390400
transform 1 0 23968 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_214
timestamp 1669390400
transform 1 0 25312 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_218
timestamp 1669390400
transform 1 0 25760 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_222
timestamp 1669390400
transform 1 0 26208 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_232
timestamp 1669390400
transform 1 0 27328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_250
timestamp 1669390400
transform 1 0 29344 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_268
timestamp 1669390400
transform 1 0 31360 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_272
timestamp 1669390400
transform 1 0 31808 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_286
timestamp 1669390400
transform 1 0 33376 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_290
timestamp 1669390400
transform 1 0 33824 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_306
timestamp 1669390400
transform 1 0 35616 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_310
timestamp 1669390400
transform 1 0 36064 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_312
timestamp 1669390400
transform 1 0 36288 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_315
timestamp 1669390400
transform 1 0 36624 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_321
timestamp 1669390400
transform 1 0 37296 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_324
timestamp 1669390400
transform 1 0 37632 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_326
timestamp 1669390400
transform 1 0 37856 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_329
timestamp 1669390400
transform 1 0 38192 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_336
timestamp 1669390400
transform 1 0 38976 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_340
timestamp 1669390400
transform 1 0 39424 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_344
timestamp 1669390400
transform 1 0 39872 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_348
timestamp 1669390400
transform 1 0 40320 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_352
timestamp 1669390400
transform 1 0 40768 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_356
timestamp 1669390400
transform 1 0 41216 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_360
timestamp 1669390400
transform 1 0 41664 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_364
timestamp 1669390400
transform 1 0 42112 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_368
timestamp 1669390400
transform 1 0 42560 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_376
timestamp 1669390400
transform 1 0 43456 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_384
timestamp 1669390400
transform 1 0 44352 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_388
timestamp 1669390400
transform 1 0 44800 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_392
timestamp 1669390400
transform 1 0 45248 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_401
timestamp 1669390400
transform 1 0 46256 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_403
timestamp 1669390400
transform 1 0 46480 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_412
timestamp 1669390400
transform 1 0 47488 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_450
timestamp 1669390400
transform 1 0 51744 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_460
timestamp 1669390400
transform 1 0 52864 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_463
timestamp 1669390400
transform 1 0 53200 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_474
timestamp 1669390400
transform 1 0 54432 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_478
timestamp 1669390400
transform 1 0 54880 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_482
timestamp 1669390400
transform 1 0 55328 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_486
timestamp 1669390400
transform 1 0 55776 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_492
timestamp 1669390400
transform 1 0 56448 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_506
timestamp 1669390400
transform 1 0 58016 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_508
timestamp 1669390400
transform 1 0 58240 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_2
timestamp 1669390400
transform 1 0 1568 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_18
timestamp 1669390400
transform 1 0 3360 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_22
timestamp 1669390400
transform 1 0 3808 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_25
timestamp 1669390400
transform 1 0 4144 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_36
timestamp 1669390400
transform 1 0 5376 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_40
timestamp 1669390400
transform 1 0 5824 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_46
timestamp 1669390400
transform 1 0 6496 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_57
timestamp 1669390400
transform 1 0 7728 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_61
timestamp 1669390400
transform 1 0 8176 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_69
timestamp 1669390400
transform 1 0 9072 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_73
timestamp 1669390400
transform 1 0 9520 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_83
timestamp 1669390400
transform 1 0 10640 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_87
timestamp 1669390400
transform 1 0 11088 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_91
timestamp 1669390400
transform 1 0 11536 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_99
timestamp 1669390400
transform 1 0 12432 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_101
timestamp 1669390400
transform 1 0 12656 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_104
timestamp 1669390400
transform 1 0 12992 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_113
timestamp 1669390400
transform 1 0 14000 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_131
timestamp 1669390400
transform 1 0 16016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1669390400
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_144
timestamp 1669390400
transform 1 0 17472 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_147
timestamp 1669390400
transform 1 0 17808 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_159
timestamp 1669390400
transform 1 0 19152 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_186
timestamp 1669390400
transform 1 0 22176 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_192
timestamp 1669390400
transform 1 0 22848 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_212
timestamp 1669390400
transform 1 0 25088 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_215
timestamp 1669390400
transform 1 0 25424 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_221
timestamp 1669390400
transform 1 0 26096 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_225
timestamp 1669390400
transform 1 0 26544 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_229
timestamp 1669390400
transform 1 0 26992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_236
timestamp 1669390400
transform 1 0 27776 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_240
timestamp 1669390400
transform 1 0 28224 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_257
timestamp 1669390400
transform 1 0 30128 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_261
timestamp 1669390400
transform 1 0 30576 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_276
timestamp 1669390400
transform 1 0 32256 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1669390400
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_286
timestamp 1669390400
transform 1 0 33376 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_299
timestamp 1669390400
transform 1 0 34832 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_313
timestamp 1669390400
transform 1 0 36400 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_323
timestamp 1669390400
transform 1 0 37520 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_325
timestamp 1669390400
transform 1 0 37744 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_328
timestamp 1669390400
transform 1 0 38080 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_332
timestamp 1669390400
transform 1 0 38528 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_336
timestamp 1669390400
transform 1 0 38976 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_346
timestamp 1669390400
transform 1 0 40096 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_350
timestamp 1669390400
transform 1 0 40544 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_354
timestamp 1669390400
transform 1 0 40992 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_357
timestamp 1669390400
transform 1 0 41328 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_368
timestamp 1669390400
transform 1 0 42560 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_372
timestamp 1669390400
transform 1 0 43008 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_376
timestamp 1669390400
transform 1 0 43456 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_378
timestamp 1669390400
transform 1 0 43680 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_387
timestamp 1669390400
transform 1 0 44688 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_391
timestamp 1669390400
transform 1 0 45136 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_395
timestamp 1669390400
transform 1 0 45584 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_399
timestamp 1669390400
transform 1 0 46032 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_407
timestamp 1669390400
transform 1 0 46928 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_424
timestamp 1669390400
transform 1 0 48832 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_428
timestamp 1669390400
transform 1 0 49280 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_431
timestamp 1669390400
transform 1 0 49616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_442
timestamp 1669390400
transform 1 0 50848 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_446
timestamp 1669390400
transform 1 0 51296 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_450
timestamp 1669390400
transform 1 0 51744 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_477
timestamp 1669390400
transform 1 0 54768 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_493
timestamp 1669390400
transform 1 0 56560 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_499
timestamp 1669390400
transform 1 0 57232 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_502
timestamp 1669390400
transform 1 0 57568 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_506
timestamp 1669390400
transform 1 0 58016 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_508
timestamp 1669390400
transform 1 0 58240 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_2
timestamp 1669390400
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_18
timestamp 1669390400
transform 1 0 3360 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_21
timestamp 1669390400
transform 1 0 3696 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1669390400
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_37
timestamp 1669390400
transform 1 0 5488 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_47
timestamp 1669390400
transform 1 0 6608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_63
timestamp 1669390400
transform 1 0 8400 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_67
timestamp 1669390400
transform 1 0 8848 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_71
timestamp 1669390400
transform 1 0 9296 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_81
timestamp 1669390400
transform 1 0 10416 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_92
timestamp 1669390400
transform 1 0 11648 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_94
timestamp 1669390400
transform 1 0 11872 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1669390400
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_108
timestamp 1669390400
transform 1 0 13440 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_126
timestamp 1669390400
transform 1 0 15456 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_138
timestamp 1669390400
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_150
timestamp 1669390400
transform 1 0 18144 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_158
timestamp 1669390400
transform 1 0 19040 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_160
timestamp 1669390400
transform 1 0 19264 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_169
timestamp 1669390400
transform 1 0 20272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_173
timestamp 1669390400
transform 1 0 20720 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1669390400
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1669390400
transform 1 0 21392 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_182
timestamp 1669390400
transform 1 0 21728 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_190
timestamp 1669390400
transform 1 0 22624 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_194
timestamp 1669390400
transform 1 0 23072 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_197
timestamp 1669390400
transform 1 0 23408 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_232
timestamp 1669390400
transform 1 0 27328 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_246
timestamp 1669390400
transform 1 0 28896 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_250
timestamp 1669390400
transform 1 0 29344 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_259
timestamp 1669390400
transform 1 0 30352 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_267
timestamp 1669390400
transform 1 0 31248 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_274
timestamp 1669390400
transform 1 0 32032 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_278
timestamp 1669390400
transform 1 0 32480 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_282
timestamp 1669390400
transform 1 0 32928 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_294
timestamp 1669390400
transform 1 0 34272 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_305
timestamp 1669390400
transform 1 0 35504 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_318
timestamp 1669390400
transform 1 0 36960 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_321
timestamp 1669390400
transform 1 0 37296 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_327
timestamp 1669390400
transform 1 0 37968 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_333
timestamp 1669390400
transform 1 0 38640 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_341
timestamp 1669390400
transform 1 0 39536 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_355
timestamp 1669390400
transform 1 0 41104 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_365
timestamp 1669390400
transform 1 0 42224 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_379
timestamp 1669390400
transform 1 0 43792 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_383
timestamp 1669390400
transform 1 0 44240 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_387
timestamp 1669390400
transform 1 0 44688 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1669390400
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_392
timestamp 1669390400
transform 1 0 45248 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_398
timestamp 1669390400
transform 1 0 45920 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_402
timestamp 1669390400
transform 1 0 46368 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_406
timestamp 1669390400
transform 1 0 46816 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_410
timestamp 1669390400
transform 1 0 47264 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_414
timestamp 1669390400
transform 1 0 47712 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_417
timestamp 1669390400
transform 1 0 48048 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_421
timestamp 1669390400
transform 1 0 48496 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_425
timestamp 1669390400
transform 1 0 48944 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_427
timestamp 1669390400
transform 1 0 49168 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_430
timestamp 1669390400
transform 1 0 49504 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_434
timestamp 1669390400
transform 1 0 49952 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_438
timestamp 1669390400
transform 1 0 50400 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_442
timestamp 1669390400
transform 1 0 50848 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_446
timestamp 1669390400
transform 1 0 51296 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_460
timestamp 1669390400
transform 1 0 52864 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_463
timestamp 1669390400
transform 1 0 53200 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_466
timestamp 1669390400
transform 1 0 53536 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_470
timestamp 1669390400
transform 1 0 53984 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_474
timestamp 1669390400
transform 1 0 54432 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_481
timestamp 1669390400
transform 1 0 55216 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_496
timestamp 1669390400
transform 1 0 56896 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_506
timestamp 1669390400
transform 1 0 58016 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_508
timestamp 1669390400
transform 1 0 58240 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_2
timestamp 1669390400
transform 1 0 1568 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_18
timestamp 1669390400
transform 1 0 3360 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_22
timestamp 1669390400
transform 1 0 3808 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_26
timestamp 1669390400
transform 1 0 4256 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_39
timestamp 1669390400
transform 1 0 5712 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_45
timestamp 1669390400
transform 1 0 6384 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_49
timestamp 1669390400
transform 1 0 6832 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_58
timestamp 1669390400
transform 1 0 7840 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_62
timestamp 1669390400
transform 1 0 8288 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1669390400
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_73
timestamp 1669390400
transform 1 0 9520 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_79
timestamp 1669390400
transform 1 0 10192 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_92
timestamp 1669390400
transform 1 0 11648 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_94
timestamp 1669390400
transform 1 0 11872 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_97
timestamp 1669390400
transform 1 0 12208 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_101
timestamp 1669390400
transform 1 0 12656 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_105
timestamp 1669390400
transform 1 0 13104 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_109
timestamp 1669390400
transform 1 0 13552 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_123
timestamp 1669390400
transform 1 0 15120 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_130
timestamp 1669390400
transform 1 0 15904 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_134
timestamp 1669390400
transform 1 0 16352 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1669390400
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_144
timestamp 1669390400
transform 1 0 17472 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_156
timestamp 1669390400
transform 1 0 18816 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_158
timestamp 1669390400
transform 1 0 19040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_161
timestamp 1669390400
transform 1 0 19376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_167
timestamp 1669390400
transform 1 0 20048 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_171
timestamp 1669390400
transform 1 0 20496 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_179
timestamp 1669390400
transform 1 0 21392 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_191
timestamp 1669390400
transform 1 0 22736 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_195
timestamp 1669390400
transform 1 0 23184 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_201
timestamp 1669390400
transform 1 0 23856 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_208
timestamp 1669390400
transform 1 0 24640 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1669390400
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_215
timestamp 1669390400
transform 1 0 25424 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_234
timestamp 1669390400
transform 1 0 27552 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_238
timestamp 1669390400
transform 1 0 28000 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_242
timestamp 1669390400
transform 1 0 28448 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_263
timestamp 1669390400
transform 1 0 30800 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_279
timestamp 1669390400
transform 1 0 32592 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1669390400
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_286
timestamp 1669390400
transform 1 0 33376 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_297
timestamp 1669390400
transform 1 0 34608 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_307
timestamp 1669390400
transform 1 0 35728 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_317
timestamp 1669390400
transform 1 0 36848 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_321
timestamp 1669390400
transform 1 0 37296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_333
timestamp 1669390400
transform 1 0 38640 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_343
timestamp 1669390400
transform 1 0 39760 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_345
timestamp 1669390400
transform 1 0 39984 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_348
timestamp 1669390400
transform 1 0 40320 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_352
timestamp 1669390400
transform 1 0 40768 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_354
timestamp 1669390400
transform 1 0 40992 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_357
timestamp 1669390400
transform 1 0 41328 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_365
timestamp 1669390400
transform 1 0 42224 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_369
timestamp 1669390400
transform 1 0 42672 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_371
timestamp 1669390400
transform 1 0 42896 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_391
timestamp 1669390400
transform 1 0 45136 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_401
timestamp 1669390400
transform 1 0 46256 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_405
timestamp 1669390400
transform 1 0 46704 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_409
timestamp 1669390400
transform 1 0 47152 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_415
timestamp 1669390400
transform 1 0 47824 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_422
timestamp 1669390400
transform 1 0 48608 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_428
timestamp 1669390400
transform 1 0 49280 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_441
timestamp 1669390400
transform 1 0 50736 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_445
timestamp 1669390400
transform 1 0 51184 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_449
timestamp 1669390400
transform 1 0 51632 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_453
timestamp 1669390400
transform 1 0 52080 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_457
timestamp 1669390400
transform 1 0 52528 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_461
timestamp 1669390400
transform 1 0 52976 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_475
timestamp 1669390400
transform 1 0 54544 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_479
timestamp 1669390400
transform 1 0 54992 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_483
timestamp 1669390400
transform 1 0 55440 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_495
timestamp 1669390400
transform 1 0 56784 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_499
timestamp 1669390400
transform 1 0 57232 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_505
timestamp 1669390400
transform 1 0 57904 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_2
timestamp 1669390400
transform 1 0 1568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_6
timestamp 1669390400
transform 1 0 2016 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_14
timestamp 1669390400
transform 1 0 2912 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_18
timestamp 1669390400
transform 1 0 3360 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_22
timestamp 1669390400
transform 1 0 3808 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1669390400
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_37
timestamp 1669390400
transform 1 0 5488 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_50
timestamp 1669390400
transform 1 0 6944 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_54
timestamp 1669390400
transform 1 0 7392 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_58
timestamp 1669390400
transform 1 0 7840 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_70
timestamp 1669390400
transform 1 0 9184 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_74
timestamp 1669390400
transform 1 0 9632 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_77
timestamp 1669390400
transform 1 0 9968 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_85
timestamp 1669390400
transform 1 0 10864 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_89
timestamp 1669390400
transform 1 0 11312 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_93
timestamp 1669390400
transform 1 0 11760 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_97
timestamp 1669390400
transform 1 0 12208 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_101
timestamp 1669390400
transform 1 0 12656 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1669390400
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_108
timestamp 1669390400
transform 1 0 13440 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_119
timestamp 1669390400
transform 1 0 14672 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_121
timestamp 1669390400
transform 1 0 14896 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_124
timestamp 1669390400
transform 1 0 15232 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_128
timestamp 1669390400
transform 1 0 15680 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_130
timestamp 1669390400
transform 1 0 15904 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_133
timestamp 1669390400
transform 1 0 16240 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_139
timestamp 1669390400
transform 1 0 16912 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_143
timestamp 1669390400
transform 1 0 17360 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_151
timestamp 1669390400
transform 1 0 18256 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_155
timestamp 1669390400
transform 1 0 18704 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_159
timestamp 1669390400
transform 1 0 19152 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1669390400
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1669390400
transform 1 0 21392 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_188
timestamp 1669390400
transform 1 0 22400 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_190
timestamp 1669390400
transform 1 0 22624 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_193
timestamp 1669390400
transform 1 0 22960 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_197
timestamp 1669390400
transform 1 0 23408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_205
timestamp 1669390400
transform 1 0 24304 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_207
timestamp 1669390400
transform 1 0 24528 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_210
timestamp 1669390400
transform 1 0 24864 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_216
timestamp 1669390400
transform 1 0 25536 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_220
timestamp 1669390400
transform 1 0 25984 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_236
timestamp 1669390400
transform 1 0 27776 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_244
timestamp 1669390400
transform 1 0 28672 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_250
timestamp 1669390400
transform 1 0 29344 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_257
timestamp 1669390400
transform 1 0 30128 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_263
timestamp 1669390400
transform 1 0 30800 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_278
timestamp 1669390400
transform 1 0 32480 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_293
timestamp 1669390400
transform 1 0 34160 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_301
timestamp 1669390400
transform 1 0 35056 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_303
timestamp 1669390400
transform 1 0 35280 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_309
timestamp 1669390400
transform 1 0 35952 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_313
timestamp 1669390400
transform 1 0 36400 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_317
timestamp 1669390400
transform 1 0 36848 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_321
timestamp 1669390400
transform 1 0 37296 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_323
timestamp 1669390400
transform 1 0 37520 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_329
timestamp 1669390400
transform 1 0 38192 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_341
timestamp 1669390400
transform 1 0 39536 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_345
timestamp 1669390400
transform 1 0 39984 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_349
timestamp 1669390400
transform 1 0 40432 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_353
timestamp 1669390400
transform 1 0 40880 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_357
timestamp 1669390400
transform 1 0 41328 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_361
timestamp 1669390400
transform 1 0 41776 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_365
timestamp 1669390400
transform 1 0 42224 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_377
timestamp 1669390400
transform 1 0 43568 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_383
timestamp 1669390400
transform 1 0 44240 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_387
timestamp 1669390400
transform 1 0 44688 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_389
timestamp 1669390400
transform 1 0 44912 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_392
timestamp 1669390400
transform 1 0 45248 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_395
timestamp 1669390400
transform 1 0 45584 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_397
timestamp 1669390400
transform 1 0 45808 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_408
timestamp 1669390400
transform 1 0 47040 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_412
timestamp 1669390400
transform 1 0 47488 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_419
timestamp 1669390400
transform 1 0 48272 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_423
timestamp 1669390400
transform 1 0 48720 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_425
timestamp 1669390400
transform 1 0 48944 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_460
timestamp 1669390400
transform 1 0 52864 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_463
timestamp 1669390400
transform 1 0 53200 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_466
timestamp 1669390400
transform 1 0 53536 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_470
timestamp 1669390400
transform 1 0 53984 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_474
timestamp 1669390400
transform 1 0 54432 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_476
timestamp 1669390400
transform 1 0 54656 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_482
timestamp 1669390400
transform 1 0 55328 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_492
timestamp 1669390400
transform 1 0 56448 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_506
timestamp 1669390400
transform 1 0 58016 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_508
timestamp 1669390400
transform 1 0 58240 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_2
timestamp 1669390400
transform 1 0 1568 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_17
timestamp 1669390400
transform 1 0 3248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_25
timestamp 1669390400
transform 1 0 4144 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_29
timestamp 1669390400
transform 1 0 4592 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_31
timestamp 1669390400
transform 1 0 4816 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_34
timestamp 1669390400
transform 1 0 5152 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_38
timestamp 1669390400
transform 1 0 5600 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_42
timestamp 1669390400
transform 1 0 6048 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_46
timestamp 1669390400
transform 1 0 6496 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_50
timestamp 1669390400
transform 1 0 6944 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_63
timestamp 1669390400
transform 1 0 8400 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_67
timestamp 1669390400
transform 1 0 8848 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1669390400
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_73
timestamp 1669390400
transform 1 0 9520 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_82
timestamp 1669390400
transform 1 0 10528 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_86
timestamp 1669390400
transform 1 0 10976 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_89
timestamp 1669390400
transform 1 0 11312 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_93
timestamp 1669390400
transform 1 0 11760 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_107
timestamp 1669390400
transform 1 0 13328 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_119
timestamp 1669390400
transform 1 0 14672 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_123
timestamp 1669390400
transform 1 0 15120 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_126
timestamp 1669390400
transform 1 0 15456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_136
timestamp 1669390400
transform 1 0 16576 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_140
timestamp 1669390400
transform 1 0 17024 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_144
timestamp 1669390400
transform 1 0 17472 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_148
timestamp 1669390400
transform 1 0 17920 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_152
timestamp 1669390400
transform 1 0 18368 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_156
timestamp 1669390400
transform 1 0 18816 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_166
timestamp 1669390400
transform 1 0 19936 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_176
timestamp 1669390400
transform 1 0 21056 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_178
timestamp 1669390400
transform 1 0 21280 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_184
timestamp 1669390400
transform 1 0 21952 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_188
timestamp 1669390400
transform 1 0 22400 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_192
timestamp 1669390400
transform 1 0 22848 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_198
timestamp 1669390400
transform 1 0 23520 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_212
timestamp 1669390400
transform 1 0 25088 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_215
timestamp 1669390400
transform 1 0 25424 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_222
timestamp 1669390400
transform 1 0 26208 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_238
timestamp 1669390400
transform 1 0 28000 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_252
timestamp 1669390400
transform 1 0 29568 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_254
timestamp 1669390400
transform 1 0 29792 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_257
timestamp 1669390400
transform 1 0 30128 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_272
timestamp 1669390400
transform 1 0 31808 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_280
timestamp 1669390400
transform 1 0 32704 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_286
timestamp 1669390400
transform 1 0 33376 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_292
timestamp 1669390400
transform 1 0 34048 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_296
timestamp 1669390400
transform 1 0 34496 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_305
timestamp 1669390400
transform 1 0 35504 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_315
timestamp 1669390400
transform 1 0 36624 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_319
timestamp 1669390400
transform 1 0 37072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_323
timestamp 1669390400
transform 1 0 37520 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_335
timestamp 1669390400
transform 1 0 38864 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_339
timestamp 1669390400
transform 1 0 39312 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_343
timestamp 1669390400
transform 1 0 39760 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_347
timestamp 1669390400
transform 1 0 40208 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_351
timestamp 1669390400
transform 1 0 40656 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_357
timestamp 1669390400
transform 1 0 41328 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_366
timestamp 1669390400
transform 1 0 42336 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_368
timestamp 1669390400
transform 1 0 42560 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_376
timestamp 1669390400
transform 1 0 43456 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_378
timestamp 1669390400
transform 1 0 43680 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_389
timestamp 1669390400
transform 1 0 44912 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_393
timestamp 1669390400
transform 1 0 45360 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_397
timestamp 1669390400
transform 1 0 45808 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_399
timestamp 1669390400
transform 1 0 46032 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_415
timestamp 1669390400
transform 1 0 47824 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_425
timestamp 1669390400
transform 1 0 48944 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_428
timestamp 1669390400
transform 1 0 49280 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_435
timestamp 1669390400
transform 1 0 50064 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_439
timestamp 1669390400
transform 1 0 50512 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_443
timestamp 1669390400
transform 1 0 50960 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_447
timestamp 1669390400
transform 1 0 51408 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_449
timestamp 1669390400
transform 1 0 51632 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_460
timestamp 1669390400
transform 1 0 52864 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_464
timestamp 1669390400
transform 1 0 53312 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_468
timestamp 1669390400
transform 1 0 53760 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_475
timestamp 1669390400
transform 1 0 54544 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_477
timestamp 1669390400
transform 1 0 54768 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_482
timestamp 1669390400
transform 1 0 55328 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_496
timestamp 1669390400
transform 1 0 56896 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_499
timestamp 1669390400
transform 1 0 57232 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_502
timestamp 1669390400
transform 1 0 57568 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_506
timestamp 1669390400
transform 1 0 58016 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_508
timestamp 1669390400
transform 1 0 58240 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_2
timestamp 1669390400
transform 1 0 1568 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_4
timestamp 1669390400
transform 1 0 1792 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_17
timestamp 1669390400
transform 1 0 3248 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_25
timestamp 1669390400
transform 1 0 4144 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_33
timestamp 1669390400
transform 1 0 5040 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_37
timestamp 1669390400
transform 1 0 5488 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_48
timestamp 1669390400
transform 1 0 6720 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_54
timestamp 1669390400
transform 1 0 7392 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_65
timestamp 1669390400
transform 1 0 8624 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_77
timestamp 1669390400
transform 1 0 9968 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_87
timestamp 1669390400
transform 1 0 11088 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_93
timestamp 1669390400
transform 1 0 11760 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_97
timestamp 1669390400
transform 1 0 12208 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_101
timestamp 1669390400
transform 1 0 12656 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1669390400
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_108
timestamp 1669390400
transform 1 0 13440 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_117
timestamp 1669390400
transform 1 0 14448 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_121
timestamp 1669390400
transform 1 0 14896 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_124
timestamp 1669390400
transform 1 0 15232 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_139
timestamp 1669390400
transform 1 0 16912 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_153
timestamp 1669390400
transform 1 0 18480 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_157
timestamp 1669390400
transform 1 0 18928 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_165
timestamp 1669390400
transform 1 0 19824 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_169
timestamp 1669390400
transform 1 0 20272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_173
timestamp 1669390400
transform 1 0 20720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1669390400
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1669390400
transform 1 0 21392 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_188
timestamp 1669390400
transform 1 0 22400 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_196
timestamp 1669390400
transform 1 0 23296 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_227
timestamp 1669390400
transform 1 0 26768 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_234
timestamp 1669390400
transform 1 0 27552 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_238
timestamp 1669390400
transform 1 0 28000 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_247
timestamp 1669390400
transform 1 0 29008 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_250
timestamp 1669390400
transform 1 0 29344 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_259
timestamp 1669390400
transform 1 0 30352 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_267
timestamp 1669390400
transform 1 0 31248 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_274
timestamp 1669390400
transform 1 0 32032 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_282
timestamp 1669390400
transform 1 0 32928 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_286
timestamp 1669390400
transform 1 0 33376 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_296
timestamp 1669390400
transform 1 0 34496 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_315
timestamp 1669390400
transform 1 0 36624 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_321
timestamp 1669390400
transform 1 0 37296 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_324
timestamp 1669390400
transform 1 0 37632 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_328
timestamp 1669390400
transform 1 0 38080 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_339
timestamp 1669390400
transform 1 0 39312 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_347
timestamp 1669390400
transform 1 0 40208 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_351
timestamp 1669390400
transform 1 0 40656 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_361
timestamp 1669390400
transform 1 0 41776 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_373
timestamp 1669390400
transform 1 0 43120 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_381
timestamp 1669390400
transform 1 0 44016 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_389
timestamp 1669390400
transform 1 0 44912 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_392
timestamp 1669390400
transform 1 0 45248 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_395
timestamp 1669390400
transform 1 0 45584 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_399
timestamp 1669390400
transform 1 0 46032 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_408
timestamp 1669390400
transform 1 0 47040 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_412
timestamp 1669390400
transform 1 0 47488 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_419
timestamp 1669390400
transform 1 0 48272 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_423
timestamp 1669390400
transform 1 0 48720 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_430
timestamp 1669390400
transform 1 0 49504 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_434
timestamp 1669390400
transform 1 0 49952 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_438
timestamp 1669390400
transform 1 0 50400 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_442
timestamp 1669390400
transform 1 0 50848 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_448
timestamp 1669390400
transform 1 0 51520 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_452
timestamp 1669390400
transform 1 0 51968 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_456
timestamp 1669390400
transform 1 0 52416 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_460
timestamp 1669390400
transform 1 0 52864 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_463
timestamp 1669390400
transform 1 0 53200 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_487
timestamp 1669390400
transform 1 0 55888 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_494
timestamp 1669390400
transform 1 0 56672 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_498
timestamp 1669390400
transform 1 0 57120 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_502
timestamp 1669390400
transform 1 0 57568 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_506
timestamp 1669390400
transform 1 0 58016 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_508
timestamp 1669390400
transform 1 0 58240 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_2
timestamp 1669390400
transform 1 0 1568 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_26
timestamp 1669390400
transform 1 0 4256 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_34
timestamp 1669390400
transform 1 0 5152 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_43
timestamp 1669390400
transform 1 0 6160 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_52
timestamp 1669390400
transform 1 0 7168 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_60
timestamp 1669390400
transform 1 0 8064 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_64
timestamp 1669390400
transform 1 0 8512 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_67
timestamp 1669390400
transform 1 0 8848 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_73
timestamp 1669390400
transform 1 0 9520 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_80
timestamp 1669390400
transform 1 0 10304 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_86
timestamp 1669390400
transform 1 0 10976 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_90
timestamp 1669390400
transform 1 0 11424 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_94
timestamp 1669390400
transform 1 0 11872 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_96
timestamp 1669390400
transform 1 0 12096 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_109
timestamp 1669390400
transform 1 0 13552 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_119
timestamp 1669390400
transform 1 0 14672 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_123
timestamp 1669390400
transform 1 0 15120 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_125
timestamp 1669390400
transform 1 0 15344 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1669390400
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_144
timestamp 1669390400
transform 1 0 17472 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_147
timestamp 1669390400
transform 1 0 17808 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_151
timestamp 1669390400
transform 1 0 18256 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_155
timestamp 1669390400
transform 1 0 18704 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_159
timestamp 1669390400
transform 1 0 19152 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_163
timestamp 1669390400
transform 1 0 19600 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_169
timestamp 1669390400
transform 1 0 20272 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_176
timestamp 1669390400
transform 1 0 21056 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_180
timestamp 1669390400
transform 1 0 21504 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_212
timestamp 1669390400
transform 1 0 25088 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_215
timestamp 1669390400
transform 1 0 25424 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_224
timestamp 1669390400
transform 1 0 26432 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_228
timestamp 1669390400
transform 1 0 26880 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_260
timestamp 1669390400
transform 1 0 30464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_264
timestamp 1669390400
transform 1 0 30912 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_279
timestamp 1669390400
transform 1 0 32592 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_283
timestamp 1669390400
transform 1 0 33040 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_286
timestamp 1669390400
transform 1 0 33376 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_289
timestamp 1669390400
transform 1 0 33712 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_303
timestamp 1669390400
transform 1 0 35280 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_313
timestamp 1669390400
transform 1 0 36400 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_323
timestamp 1669390400
transform 1 0 37520 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_330
timestamp 1669390400
transform 1 0 38304 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_341
timestamp 1669390400
transform 1 0 39536 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_351
timestamp 1669390400
transform 1 0 40656 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_357
timestamp 1669390400
transform 1 0 41328 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_395
timestamp 1669390400
transform 1 0 45584 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_397
timestamp 1669390400
transform 1 0 45808 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_408
timestamp 1669390400
transform 1 0 47040 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_425
timestamp 1669390400
transform 1 0 48944 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_428
timestamp 1669390400
transform 1 0 49280 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_430
timestamp 1669390400
transform 1 0 49504 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_445
timestamp 1669390400
transform 1 0 51184 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_449
timestamp 1669390400
transform 1 0 51632 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_451
timestamp 1669390400
transform 1 0 51856 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_458
timestamp 1669390400
transform 1 0 52640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_464
timestamp 1669390400
transform 1 0 53312 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_468
timestamp 1669390400
transform 1 0 53760 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_472
timestamp 1669390400
transform 1 0 54208 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_474
timestamp 1669390400
transform 1 0 54432 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_477
timestamp 1669390400
transform 1 0 54768 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_479
timestamp 1669390400
transform 1 0 54992 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_486
timestamp 1669390400
transform 1 0 55776 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_496
timestamp 1669390400
transform 1 0 56896 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_499
timestamp 1669390400
transform 1 0 57232 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_502
timestamp 1669390400
transform 1 0 57568 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_506
timestamp 1669390400
transform 1 0 58016 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_508
timestamp 1669390400
transform 1 0 58240 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_2
timestamp 1669390400
transform 1 0 1568 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_10
timestamp 1669390400
transform 1 0 2464 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_12
timestamp 1669390400
transform 1 0 2688 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_21
timestamp 1669390400
transform 1 0 3696 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_29
timestamp 1669390400
transform 1 0 4592 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1669390400
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_37
timestamp 1669390400
transform 1 0 5488 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_41
timestamp 1669390400
transform 1 0 5936 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_55
timestamp 1669390400
transform 1 0 7504 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_59
timestamp 1669390400
transform 1 0 7952 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_75
timestamp 1669390400
transform 1 0 9744 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_83
timestamp 1669390400
transform 1 0 10640 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_92
timestamp 1669390400
transform 1 0 11648 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_96
timestamp 1669390400
transform 1 0 12096 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_100
timestamp 1669390400
transform 1 0 12544 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_102
timestamp 1669390400
transform 1 0 12768 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1669390400
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_108
timestamp 1669390400
transform 1 0 13440 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_116
timestamp 1669390400
transform 1 0 14336 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_118
timestamp 1669390400
transform 1 0 14560 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_121
timestamp 1669390400
transform 1 0 14896 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_131
timestamp 1669390400
transform 1 0 16016 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_135
timestamp 1669390400
transform 1 0 16464 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_141
timestamp 1669390400
transform 1 0 17136 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_147
timestamp 1669390400
transform 1 0 17808 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_151
timestamp 1669390400
transform 1 0 18256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_157
timestamp 1669390400
transform 1 0 18928 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_159
timestamp 1669390400
transform 1 0 19152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_166
timestamp 1669390400
transform 1 0 19936 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_172
timestamp 1669390400
transform 1 0 20608 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1669390400
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_179
timestamp 1669390400
transform 1 0 21392 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_200
timestamp 1669390400
transform 1 0 23744 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_208
timestamp 1669390400
transform 1 0 24640 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_216
timestamp 1669390400
transform 1 0 25536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_220
timestamp 1669390400
transform 1 0 25984 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_222
timestamp 1669390400
transform 1 0 26208 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_225
timestamp 1669390400
transform 1 0 26544 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_233
timestamp 1669390400
transform 1 0 27440 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1669390400
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_250
timestamp 1669390400
transform 1 0 29344 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_252
timestamp 1669390400
transform 1 0 29568 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_263
timestamp 1669390400
transform 1 0 30800 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_275
timestamp 1669390400
transform 1 0 32144 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_285
timestamp 1669390400
transform 1 0 33264 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_289
timestamp 1669390400
transform 1 0 33712 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_293
timestamp 1669390400
transform 1 0 34160 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_297
timestamp 1669390400
transform 1 0 34608 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_300
timestamp 1669390400
transform 1 0 34944 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_308
timestamp 1669390400
transform 1 0 35840 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_312
timestamp 1669390400
transform 1 0 36288 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_314
timestamp 1669390400
transform 1 0 36512 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_317
timestamp 1669390400
transform 1 0 36848 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_321
timestamp 1669390400
transform 1 0 37296 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_333
timestamp 1669390400
transform 1 0 38640 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_337
timestamp 1669390400
transform 1 0 39088 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_349
timestamp 1669390400
transform 1 0 40432 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_359
timestamp 1669390400
transform 1 0 41552 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_363
timestamp 1669390400
transform 1 0 42000 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_367
timestamp 1669390400
transform 1 0 42448 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_378
timestamp 1669390400
transform 1 0 43680 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_386
timestamp 1669390400
transform 1 0 44576 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_392
timestamp 1669390400
transform 1 0 45248 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_394
timestamp 1669390400
transform 1 0 45472 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_406
timestamp 1669390400
transform 1 0 46816 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_410
timestamp 1669390400
transform 1 0 47264 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_414
timestamp 1669390400
transform 1 0 47712 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_418
timestamp 1669390400
transform 1 0 48160 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_422
timestamp 1669390400
transform 1 0 48608 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_426
timestamp 1669390400
transform 1 0 49056 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_430
timestamp 1669390400
transform 1 0 49504 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_434
timestamp 1669390400
transform 1 0 49952 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_451
timestamp 1669390400
transform 1 0 51856 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_459
timestamp 1669390400
transform 1 0 52752 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_463
timestamp 1669390400
transform 1 0 53200 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_466
timestamp 1669390400
transform 1 0 53536 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_473
timestamp 1669390400
transform 1 0 54320 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_483
timestamp 1669390400
transform 1 0 55440 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_497
timestamp 1669390400
transform 1 0 57008 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_501
timestamp 1669390400
transform 1 0 57456 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_505
timestamp 1669390400
transform 1 0 57904 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_2
timestamp 1669390400
transform 1 0 1568 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_10
timestamp 1669390400
transform 1 0 2464 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_45
timestamp 1669390400
transform 1 0 6384 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_54
timestamp 1669390400
transform 1 0 7392 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_58
timestamp 1669390400
transform 1 0 7840 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_66
timestamp 1669390400
transform 1 0 8736 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1669390400
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_73
timestamp 1669390400
transform 1 0 9520 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_76
timestamp 1669390400
transform 1 0 9856 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_90
timestamp 1669390400
transform 1 0 11424 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_102
timestamp 1669390400
transform 1 0 12768 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_104
timestamp 1669390400
transform 1 0 12992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_107
timestamp 1669390400
transform 1 0 13328 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_111
timestamp 1669390400
transform 1 0 13776 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_117
timestamp 1669390400
transform 1 0 14448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_131
timestamp 1669390400
transform 1 0 16016 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_140
timestamp 1669390400
transform 1 0 17024 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_144
timestamp 1669390400
transform 1 0 17472 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_146
timestamp 1669390400
transform 1 0 17696 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_155
timestamp 1669390400
transform 1 0 18704 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_163
timestamp 1669390400
transform 1 0 19600 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_165
timestamp 1669390400
transform 1 0 19824 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_177
timestamp 1669390400
transform 1 0 21168 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_181
timestamp 1669390400
transform 1 0 21616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_185
timestamp 1669390400
transform 1 0 22064 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_189
timestamp 1669390400
transform 1 0 22512 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_197
timestamp 1669390400
transform 1 0 23408 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_215
timestamp 1669390400
transform 1 0 25424 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_224
timestamp 1669390400
transform 1 0 26432 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_232
timestamp 1669390400
transform 1 0 27328 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_236
timestamp 1669390400
transform 1 0 27776 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_274
timestamp 1669390400
transform 1 0 32032 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_278
timestamp 1669390400
transform 1 0 32480 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_282
timestamp 1669390400
transform 1 0 32928 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_51_286
timestamp 1669390400
transform 1 0 33376 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_294
timestamp 1669390400
transform 1 0 34272 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_298
timestamp 1669390400
transform 1 0 34720 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_302
timestamp 1669390400
transform 1 0 35168 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_306
timestamp 1669390400
transform 1 0 35616 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_342
timestamp 1669390400
transform 1 0 39648 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_354
timestamp 1669390400
transform 1 0 40992 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_357
timestamp 1669390400
transform 1 0 41328 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_364
timestamp 1669390400
transform 1 0 42112 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_376
timestamp 1669390400
transform 1 0 43456 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_380
timestamp 1669390400
transform 1 0 43904 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_394
timestamp 1669390400
transform 1 0 45472 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_406
timestamp 1669390400
transform 1 0 46816 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_408
timestamp 1669390400
transform 1 0 47040 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_415
timestamp 1669390400
transform 1 0 47824 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_419
timestamp 1669390400
transform 1 0 48272 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_423
timestamp 1669390400
transform 1 0 48720 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_425
timestamp 1669390400
transform 1 0 48944 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_428
timestamp 1669390400
transform 1 0 49280 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_442
timestamp 1669390400
transform 1 0 50848 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_455
timestamp 1669390400
transform 1 0 52304 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_457
timestamp 1669390400
transform 1 0 52528 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_460
timestamp 1669390400
transform 1 0 52864 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_464
timestamp 1669390400
transform 1 0 53312 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_475
timestamp 1669390400
transform 1 0 54544 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_491
timestamp 1669390400
transform 1 0 56336 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_495
timestamp 1669390400
transform 1 0 56784 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_499
timestamp 1669390400
transform 1 0 57232 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_502
timestamp 1669390400
transform 1 0 57568 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_506
timestamp 1669390400
transform 1 0 58016 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_508
timestamp 1669390400
transform 1 0 58240 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_2
timestamp 1669390400
transform 1 0 1568 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_18
timestamp 1669390400
transform 1 0 3360 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_26
timestamp 1669390400
transform 1 0 4256 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_30
timestamp 1669390400
transform 1 0 4704 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1669390400
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_37
timestamp 1669390400
transform 1 0 5488 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_44
timestamp 1669390400
transform 1 0 6272 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_52
timestamp 1669390400
transform 1 0 7168 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_60
timestamp 1669390400
transform 1 0 8064 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_68
timestamp 1669390400
transform 1 0 8960 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_76
timestamp 1669390400
transform 1 0 9856 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_84
timestamp 1669390400
transform 1 0 10752 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_92
timestamp 1669390400
transform 1 0 11648 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_96
timestamp 1669390400
transform 1 0 12096 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_100
timestamp 1669390400
transform 1 0 12544 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_104
timestamp 1669390400
transform 1 0 12992 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_108
timestamp 1669390400
transform 1 0 13440 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_112
timestamp 1669390400
transform 1 0 13888 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_114
timestamp 1669390400
transform 1 0 14112 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_117
timestamp 1669390400
transform 1 0 14448 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_129
timestamp 1669390400
transform 1 0 15792 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_131
timestamp 1669390400
transform 1 0 16016 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_140
timestamp 1669390400
transform 1 0 17024 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_144
timestamp 1669390400
transform 1 0 17472 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_154
timestamp 1669390400
transform 1 0 18592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_162
timestamp 1669390400
transform 1 0 19488 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1669390400
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_179
timestamp 1669390400
transform 1 0 21392 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_183
timestamp 1669390400
transform 1 0 21840 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_197
timestamp 1669390400
transform 1 0 23408 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_201
timestamp 1669390400
transform 1 0 23856 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_211
timestamp 1669390400
transform 1 0 24976 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_226
timestamp 1669390400
transform 1 0 26656 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_242
timestamp 1669390400
transform 1 0 28448 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_246
timestamp 1669390400
transform 1 0 28896 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_250
timestamp 1669390400
transform 1 0 29344 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_261
timestamp 1669390400
transform 1 0 30576 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_271
timestamp 1669390400
transform 1 0 31696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_277
timestamp 1669390400
transform 1 0 32368 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_287
timestamp 1669390400
transform 1 0 33488 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_295
timestamp 1669390400
transform 1 0 34384 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_299
timestamp 1669390400
transform 1 0 34832 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_302
timestamp 1669390400
transform 1 0 35168 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_306
timestamp 1669390400
transform 1 0 35616 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_315
timestamp 1669390400
transform 1 0 36624 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_321
timestamp 1669390400
transform 1 0 37296 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_324
timestamp 1669390400
transform 1 0 37632 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_328
timestamp 1669390400
transform 1 0 38080 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_332
timestamp 1669390400
transform 1 0 38528 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_341
timestamp 1669390400
transform 1 0 39536 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_345
timestamp 1669390400
transform 1 0 39984 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_349
timestamp 1669390400
transform 1 0 40432 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_353
timestamp 1669390400
transform 1 0 40880 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_357
timestamp 1669390400
transform 1 0 41328 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_361
timestamp 1669390400
transform 1 0 41776 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_372
timestamp 1669390400
transform 1 0 43008 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_378
timestamp 1669390400
transform 1 0 43680 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_382
timestamp 1669390400
transform 1 0 44128 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_386
timestamp 1669390400
transform 1 0 44576 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_392
timestamp 1669390400
transform 1 0 45248 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_403
timestamp 1669390400
transform 1 0 46480 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_417
timestamp 1669390400
transform 1 0 48048 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_427
timestamp 1669390400
transform 1 0 49168 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_433
timestamp 1669390400
transform 1 0 49840 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_448
timestamp 1669390400
transform 1 0 51520 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_452
timestamp 1669390400
transform 1 0 51968 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_456
timestamp 1669390400
transform 1 0 52416 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_460
timestamp 1669390400
transform 1 0 52864 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_463
timestamp 1669390400
transform 1 0 53200 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_474
timestamp 1669390400
transform 1 0 54432 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_478
timestamp 1669390400
transform 1 0 54880 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_491
timestamp 1669390400
transform 1 0 56336 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_495
timestamp 1669390400
transform 1 0 56784 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_503
timestamp 1669390400
transform 1 0 57680 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_507
timestamp 1669390400
transform 1 0 58128 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_2
timestamp 1669390400
transform 1 0 1568 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_6
timestamp 1669390400
transform 1 0 2016 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_14
timestamp 1669390400
transform 1 0 2912 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_18
timestamp 1669390400
transform 1 0 3360 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_34
timestamp 1669390400
transform 1 0 5152 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_69
timestamp 1669390400
transform 1 0 9072 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_73
timestamp 1669390400
transform 1 0 9520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_80
timestamp 1669390400
transform 1 0 10304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_86
timestamp 1669390400
transform 1 0 10976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_90
timestamp 1669390400
transform 1 0 11424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_93
timestamp 1669390400
transform 1 0 11760 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_97
timestamp 1669390400
transform 1 0 12208 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_107
timestamp 1669390400
transform 1 0 13328 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_111
timestamp 1669390400
transform 1 0 13776 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_115
timestamp 1669390400
transform 1 0 14224 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_125
timestamp 1669390400
transform 1 0 15344 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_139
timestamp 1669390400
transform 1 0 16912 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1669390400
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_144
timestamp 1669390400
transform 1 0 17472 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_147
timestamp 1669390400
transform 1 0 17808 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_151
timestamp 1669390400
transform 1 0 18256 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_155
timestamp 1669390400
transform 1 0 18704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_162
timestamp 1669390400
transform 1 0 19488 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_172
timestamp 1669390400
transform 1 0 20608 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_176
timestamp 1669390400
transform 1 0 21056 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_184
timestamp 1669390400
transform 1 0 21952 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_188
timestamp 1669390400
transform 1 0 22400 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_190
timestamp 1669390400
transform 1 0 22624 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_196
timestamp 1669390400
transform 1 0 23296 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1669390400
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_215
timestamp 1669390400
transform 1 0 25424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_222
timestamp 1669390400
transform 1 0 26208 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_228
timestamp 1669390400
transform 1 0 26880 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_244
timestamp 1669390400
transform 1 0 28672 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_260
timestamp 1669390400
transform 1 0 30464 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_268
timestamp 1669390400
transform 1 0 31360 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1669390400
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_286
timestamp 1669390400
transform 1 0 33376 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_321
timestamp 1669390400
transform 1 0 37296 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_325
timestamp 1669390400
transform 1 0 37744 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_329
timestamp 1669390400
transform 1 0 38192 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_332
timestamp 1669390400
transform 1 0 38528 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_336
timestamp 1669390400
transform 1 0 38976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_340
timestamp 1669390400
transform 1 0 39424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_343
timestamp 1669390400
transform 1 0 39760 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_353
timestamp 1669390400
transform 1 0 40880 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_357
timestamp 1669390400
transform 1 0 41328 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_360
timestamp 1669390400
transform 1 0 41664 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_364
timestamp 1669390400
transform 1 0 42112 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_389
timestamp 1669390400
transform 1 0 44912 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_409
timestamp 1669390400
transform 1 0 47152 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_421
timestamp 1669390400
transform 1 0 48496 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_425
timestamp 1669390400
transform 1 0 48944 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_428
timestamp 1669390400
transform 1 0 49280 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_464
timestamp 1669390400
transform 1 0 53312 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_477
timestamp 1669390400
transform 1 0 54768 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_481
timestamp 1669390400
transform 1 0 55216 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_485
timestamp 1669390400
transform 1 0 55664 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_489
timestamp 1669390400
transform 1 0 56112 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_493
timestamp 1669390400
transform 1 0 56560 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_499
timestamp 1669390400
transform 1 0 57232 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_506
timestamp 1669390400
transform 1 0 58016 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_508
timestamp 1669390400
transform 1 0 58240 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1669390400
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_17
timestamp 1669390400
transform 1 0 3248 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_33
timestamp 1669390400
transform 1 0 5040 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_37
timestamp 1669390400
transform 1 0 5488 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_43
timestamp 1669390400
transform 1 0 6160 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_47
timestamp 1669390400
transform 1 0 6608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_51
timestamp 1669390400
transform 1 0 7056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_54
timestamp 1669390400
transform 1 0 7392 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_58
timestamp 1669390400
transform 1 0 7840 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_62
timestamp 1669390400
transform 1 0 8288 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_80
timestamp 1669390400
transform 1 0 10304 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_84
timestamp 1669390400
transform 1 0 10752 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_88
timestamp 1669390400
transform 1 0 11200 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_92
timestamp 1669390400
transform 1 0 11648 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_95
timestamp 1669390400
transform 1 0 11984 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_105
timestamp 1669390400
transform 1 0 13104 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_108
timestamp 1669390400
transform 1 0 13440 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_117
timestamp 1669390400
transform 1 0 14448 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_54_121
timestamp 1669390400
transform 1 0 14896 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_153
timestamp 1669390400
transform 1 0 18480 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_157
timestamp 1669390400
transform 1 0 18928 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_164
timestamp 1669390400
transform 1 0 19712 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_168
timestamp 1669390400
transform 1 0 20160 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_176
timestamp 1669390400
transform 1 0 21056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_179
timestamp 1669390400
transform 1 0 21392 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_183
timestamp 1669390400
transform 1 0 21840 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_185
timestamp 1669390400
transform 1 0 22064 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_199
timestamp 1669390400
transform 1 0 23632 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_207
timestamp 1669390400
transform 1 0 24528 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_217
timestamp 1669390400
transform 1 0 25648 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_231
timestamp 1669390400
transform 1 0 27216 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1669390400
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_250
timestamp 1669390400
transform 1 0 29344 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_263
timestamp 1669390400
transform 1 0 30800 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_279
timestamp 1669390400
transform 1 0 32592 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_285
timestamp 1669390400
transform 1 0 33264 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_289
timestamp 1669390400
transform 1 0 33712 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_297
timestamp 1669390400
transform 1 0 34608 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_301
timestamp 1669390400
transform 1 0 35056 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_318
timestamp 1669390400
transform 1 0 36960 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_321
timestamp 1669390400
transform 1 0 37296 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_327
timestamp 1669390400
transform 1 0 37968 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_331
timestamp 1669390400
transform 1 0 38416 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_335
timestamp 1669390400
transform 1 0 38864 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_339
timestamp 1669390400
transform 1 0 39312 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_343
timestamp 1669390400
transform 1 0 39760 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_350
timestamp 1669390400
transform 1 0 40544 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_354
timestamp 1669390400
transform 1 0 40992 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_358
timestamp 1669390400
transform 1 0 41440 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_362
timestamp 1669390400
transform 1 0 41888 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_366
timestamp 1669390400
transform 1 0 42336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_382
timestamp 1669390400
transform 1 0 44128 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_386
timestamp 1669390400
transform 1 0 44576 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_392
timestamp 1669390400
transform 1 0 45248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_398
timestamp 1669390400
transform 1 0 45920 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_418
timestamp 1669390400
transform 1 0 48160 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_422
timestamp 1669390400
transform 1 0 48608 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_426
timestamp 1669390400
transform 1 0 49056 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_428
timestamp 1669390400
transform 1 0 49280 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_435
timestamp 1669390400
transform 1 0 50064 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_439
timestamp 1669390400
transform 1 0 50512 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_443
timestamp 1669390400
transform 1 0 50960 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_447
timestamp 1669390400
transform 1 0 51408 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_451
timestamp 1669390400
transform 1 0 51856 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_454
timestamp 1669390400
transform 1 0 52192 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_460
timestamp 1669390400
transform 1 0 52864 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_463
timestamp 1669390400
transform 1 0 53200 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_470
timestamp 1669390400
transform 1 0 53984 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_474
timestamp 1669390400
transform 1 0 54432 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_476
timestamp 1669390400
transform 1 0 54656 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_479
timestamp 1669390400
transform 1 0 54992 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_483
timestamp 1669390400
transform 1 0 55440 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_487
timestamp 1669390400
transform 1 0 55888 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_491
timestamp 1669390400
transform 1 0 56336 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_495
timestamp 1669390400
transform 1 0 56784 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_497
timestamp 1669390400
transform 1 0 57008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_500
timestamp 1669390400
transform 1 0 57344 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_504
timestamp 1669390400
transform 1 0 57792 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_508
timestamp 1669390400
transform 1 0 58240 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_55_2
timestamp 1669390400
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_66
timestamp 1669390400
transform 1 0 8736 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_70
timestamp 1669390400
transform 1 0 9184 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_73
timestamp 1669390400
transform 1 0 9520 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_86
timestamp 1669390400
transform 1 0 10976 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_94
timestamp 1669390400
transform 1 0 11872 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_98
timestamp 1669390400
transform 1 0 12320 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_100
timestamp 1669390400
transform 1 0 12544 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_103
timestamp 1669390400
transform 1 0 12880 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_107
timestamp 1669390400
transform 1 0 13328 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_109
timestamp 1669390400
transform 1 0 13552 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_118
timestamp 1669390400
transform 1 0 14560 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_134
timestamp 1669390400
transform 1 0 16352 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_141
timestamp 1669390400
transform 1 0 17136 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_144
timestamp 1669390400
transform 1 0 17472 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_148
timestamp 1669390400
transform 1 0 17920 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_150
timestamp 1669390400
transform 1 0 18144 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_156
timestamp 1669390400
transform 1 0 18816 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_55_171
timestamp 1669390400
transform 1 0 20496 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_187
timestamp 1669390400
transform 1 0 22288 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_193
timestamp 1669390400
transform 1 0 22960 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_197
timestamp 1669390400
transform 1 0 23408 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_201
timestamp 1669390400
transform 1 0 23856 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_203
timestamp 1669390400
transform 1 0 24080 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_212
timestamp 1669390400
transform 1 0 25088 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_215
timestamp 1669390400
transform 1 0 25424 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_239
timestamp 1669390400
transform 1 0 28112 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_247
timestamp 1669390400
transform 1 0 29008 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_262
timestamp 1669390400
transform 1 0 30688 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_283
timestamp 1669390400
transform 1 0 33040 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_286
timestamp 1669390400
transform 1 0 33376 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_293
timestamp 1669390400
transform 1 0 34160 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_297
timestamp 1669390400
transform 1 0 34608 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_55_301
timestamp 1669390400
transform 1 0 35056 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_309
timestamp 1669390400
transform 1 0 35952 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_313
timestamp 1669390400
transform 1 0 36400 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_315
timestamp 1669390400
transform 1 0 36624 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_328
timestamp 1669390400
transform 1 0 38080 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_332
timestamp 1669390400
transform 1 0 38528 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_336
timestamp 1669390400
transform 1 0 38976 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_343
timestamp 1669390400
transform 1 0 39760 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_354
timestamp 1669390400
transform 1 0 40992 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_357
timestamp 1669390400
transform 1 0 41328 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_360
timestamp 1669390400
transform 1 0 41664 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_366
timestamp 1669390400
transform 1 0 42336 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_378
timestamp 1669390400
transform 1 0 43680 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_388
timestamp 1669390400
transform 1 0 44800 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_392
timestamp 1669390400
transform 1 0 45248 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_396
timestamp 1669390400
transform 1 0 45696 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_400
timestamp 1669390400
transform 1 0 46144 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_414
timestamp 1669390400
transform 1 0 47712 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_422
timestamp 1669390400
transform 1 0 48608 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_428
timestamp 1669390400
transform 1 0 49280 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_435
timestamp 1669390400
transform 1 0 50064 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_439
timestamp 1669390400
transform 1 0 50512 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_443
timestamp 1669390400
transform 1 0 50960 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_55_447
timestamp 1669390400
transform 1 0 51408 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_463
timestamp 1669390400
transform 1 0 53200 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_471
timestamp 1669390400
transform 1 0 54096 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_479
timestamp 1669390400
transform 1 0 54992 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_483
timestamp 1669390400
transform 1 0 55440 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_487
timestamp 1669390400
transform 1 0 55888 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_491
timestamp 1669390400
transform 1 0 56336 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_495
timestamp 1669390400
transform 1 0 56784 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_499
timestamp 1669390400
transform 1 0 57232 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_502
timestamp 1669390400
transform 1 0 57568 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_55_506
timestamp 1669390400
transform 1 0 58016 0 -1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_55_508
timestamp 1669390400
transform 1 0 58240 0 -1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_56_2
timestamp 1669390400
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_34
timestamp 1669390400
transform 1 0 5152 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_37
timestamp 1669390400
transform 1 0 5488 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_53
timestamp 1669390400
transform 1 0 7280 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_61
timestamp 1669390400
transform 1 0 8176 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_73
timestamp 1669390400
transform 1 0 9520 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_87
timestamp 1669390400
transform 1 0 11088 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_95
timestamp 1669390400
transform 1 0 11984 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_105
timestamp 1669390400
transform 1 0 13104 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_108
timestamp 1669390400
transform 1 0 13440 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_119
timestamp 1669390400
transform 1 0 14672 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_123
timestamp 1669390400
transform 1 0 15120 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_127
timestamp 1669390400
transform 1 0 15568 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_129
timestamp 1669390400
transform 1 0 15792 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_143
timestamp 1669390400
transform 1 0 17360 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_145
timestamp 1669390400
transform 1 0 17584 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_154
timestamp 1669390400
transform 1 0 18592 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_169
timestamp 1669390400
transform 1 0 20272 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_179
timestamp 1669390400
transform 1 0 21392 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_183
timestamp 1669390400
transform 1 0 21840 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_185
timestamp 1669390400
transform 1 0 22064 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_194
timestamp 1669390400
transform 1 0 23072 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_201
timestamp 1669390400
transform 1 0 23856 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_56_205
timestamp 1669390400
transform 1 0 24304 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_213
timestamp 1669390400
transform 1 0 25200 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_226
timestamp 1669390400
transform 1 0 26656 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_242
timestamp 1669390400
transform 1 0 28448 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_246
timestamp 1669390400
transform 1 0 28896 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_250
timestamp 1669390400
transform 1 0 29344 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_254
timestamp 1669390400
transform 1 0 29792 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_56_268
timestamp 1669390400
transform 1 0 31360 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_292
timestamp 1669390400
transform 1 0 34048 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_296
timestamp 1669390400
transform 1 0 34496 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_300
timestamp 1669390400
transform 1 0 34944 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_304
timestamp 1669390400
transform 1 0 35392 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_308
timestamp 1669390400
transform 1 0 35840 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_314
timestamp 1669390400
transform 1 0 36512 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_318
timestamp 1669390400
transform 1 0 36960 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_321
timestamp 1669390400
transform 1 0 37296 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_345
timestamp 1669390400
transform 1 0 39984 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_358
timestamp 1669390400
transform 1 0 41440 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_362
timestamp 1669390400
transform 1 0 41888 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_366
timestamp 1669390400
transform 1 0 42336 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_387
timestamp 1669390400
transform 1 0 44688 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_389
timestamp 1669390400
transform 1 0 44912 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_392
timestamp 1669390400
transform 1 0 45248 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_56_395
timestamp 1669390400
transform 1 0 45584 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_439
timestamp 1669390400
transform 1 0 50512 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_455
timestamp 1669390400
transform 1 0 52304 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_459
timestamp 1669390400
transform 1 0 52752 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_56_463
timestamp 1669390400
transform 1 0 53200 0 1 47040
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_475
timestamp 1669390400
transform 1 0 54544 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_483
timestamp 1669390400
transform 1 0 55440 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_487
timestamp 1669390400
transform 1 0 55888 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_491
timestamp 1669390400
transform 1 0 56336 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_495
timestamp 1669390400
transform 1 0 56784 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_499
timestamp 1669390400
transform 1 0 57232 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_503
timestamp 1669390400
transform 1 0 57680 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_56_507
timestamp 1669390400
transform 1 0 58128 0 1 47040
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_2
timestamp 1669390400
transform 1 0 1568 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_6
timestamp 1669390400
transform 1 0 2016 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_14
timestamp 1669390400
transform 1 0 2912 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_57_18
timestamp 1669390400
transform 1 0 3360 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_57_50
timestamp 1669390400
transform 1 0 6944 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_66
timestamp 1669390400
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_70
timestamp 1669390400
transform 1 0 9184 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_73
timestamp 1669390400
transform 1 0 9520 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_83
timestamp 1669390400
transform 1 0 10640 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_96
timestamp 1669390400
transform 1 0 12096 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_121
timestamp 1669390400
transform 1 0 14896 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_125
timestamp 1669390400
transform 1 0 15344 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_141
timestamp 1669390400
transform 1 0 17136 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_144
timestamp 1669390400
transform 1 0 17472 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_153
timestamp 1669390400
transform 1 0 18480 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_168
timestamp 1669390400
transform 1 0 20160 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_176
timestamp 1669390400
transform 1 0 21056 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_179
timestamp 1669390400
transform 1 0 21392 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_186
timestamp 1669390400
transform 1 0 22176 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_201
timestamp 1669390400
transform 1 0 23856 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_208
timestamp 1669390400
transform 1 0 24640 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_212
timestamp 1669390400
transform 1 0 25088 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_215
timestamp 1669390400
transform 1 0 25424 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_219
timestamp 1669390400
transform 1 0 25872 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_222
timestamp 1669390400
transform 1 0 26208 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_57_235
timestamp 1669390400
transform 1 0 27664 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_243
timestamp 1669390400
transform 1 0 28560 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_247
timestamp 1669390400
transform 1 0 29008 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_257
timestamp 1669390400
transform 1 0 30128 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_265
timestamp 1669390400
transform 1 0 31024 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_269
timestamp 1669390400
transform 1 0 31472 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_273
timestamp 1669390400
transform 1 0 31920 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_283
timestamp 1669390400
transform 1 0 33040 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_286
timestamp 1669390400
transform 1 0 33376 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_297
timestamp 1669390400
transform 1 0 34608 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_301
timestamp 1669390400
transform 1 0 35056 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_303
timestamp 1669390400
transform 1 0 35280 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_315
timestamp 1669390400
transform 1 0 36624 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_323
timestamp 1669390400
transform 1 0 37520 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_327
timestamp 1669390400
transform 1 0 37968 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_330
timestamp 1669390400
transform 1 0 38304 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_334
timestamp 1669390400
transform 1 0 38752 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_336
timestamp 1669390400
transform 1 0 38976 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_343
timestamp 1669390400
transform 1 0 39760 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_354
timestamp 1669390400
transform 1 0 40992 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_357
timestamp 1669390400
transform 1 0 41328 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_360
timestamp 1669390400
transform 1 0 41664 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_364
timestamp 1669390400
transform 1 0 42112 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_368
timestamp 1669390400
transform 1 0 42560 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_380
timestamp 1669390400
transform 1 0 43904 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_384
timestamp 1669390400
transform 1 0 44352 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_388
timestamp 1669390400
transform 1 0 44800 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_392
timestamp 1669390400
transform 1 0 45248 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_396
timestamp 1669390400
transform 1 0 45696 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_400
timestamp 1669390400
transform 1 0 46144 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_413
timestamp 1669390400
transform 1 0 47600 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_420
timestamp 1669390400
transform 1 0 48384 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_424
timestamp 1669390400
transform 1 0 48832 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_428
timestamp 1669390400
transform 1 0 49280 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_442
timestamp 1669390400
transform 1 0 50848 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_452
timestamp 1669390400
transform 1 0 51968 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_456
timestamp 1669390400
transform 1 0 52416 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_470
timestamp 1669390400
transform 1 0 53984 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_474
timestamp 1669390400
transform 1 0 54432 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_478
timestamp 1669390400
transform 1 0 54880 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_482
timestamp 1669390400
transform 1 0 55328 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_486
timestamp 1669390400
transform 1 0 55776 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_490
timestamp 1669390400
transform 1 0 56224 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_494
timestamp 1669390400
transform 1 0 56672 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_496
timestamp 1669390400
transform 1 0 56896 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_499
timestamp 1669390400
transform 1 0 57232 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_57_502
timestamp 1669390400
transform 1 0 57568 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_57_506
timestamp 1669390400
transform 1 0 58016 0 -1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_57_508
timestamp 1669390400
transform 1 0 58240 0 -1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_2
timestamp 1669390400
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_34
timestamp 1669390400
transform 1 0 5152 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_58_37
timestamp 1669390400
transform 1 0 5488 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_69
timestamp 1669390400
transform 1 0 9072 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_73
timestamp 1669390400
transform 1 0 9520 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_82
timestamp 1669390400
transform 1 0 10528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_90
timestamp 1669390400
transform 1 0 11424 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_94
timestamp 1669390400
transform 1 0 11872 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_96
timestamp 1669390400
transform 1 0 12096 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_105
timestamp 1669390400
transform 1 0 13104 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_108
timestamp 1669390400
transform 1 0 13440 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_117
timestamp 1669390400
transform 1 0 14448 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_125
timestamp 1669390400
transform 1 0 15344 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_127
timestamp 1669390400
transform 1 0 15568 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_136
timestamp 1669390400
transform 1 0 16576 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_143
timestamp 1669390400
transform 1 0 17360 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_151
timestamp 1669390400
transform 1 0 18256 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_58_159
timestamp 1669390400
transform 1 0 19152 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_167
timestamp 1669390400
transform 1 0 20048 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_171
timestamp 1669390400
transform 1 0 20496 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_173
timestamp 1669390400
transform 1 0 20720 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_176
timestamp 1669390400
transform 1 0 21056 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_179
timestamp 1669390400
transform 1 0 21392 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_186
timestamp 1669390400
transform 1 0 22176 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_190
timestamp 1669390400
transform 1 0 22624 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_194
timestamp 1669390400
transform 1 0 23072 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_202
timestamp 1669390400
transform 1 0 23968 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_218
timestamp 1669390400
transform 1 0 25760 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_232
timestamp 1669390400
transform 1 0 27328 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_250
timestamp 1669390400
transform 1 0 29344 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_253
timestamp 1669390400
transform 1 0 29680 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_263
timestamp 1669390400
transform 1 0 30800 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_265
timestamp 1669390400
transform 1 0 31024 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_272
timestamp 1669390400
transform 1 0 31808 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_282
timestamp 1669390400
transform 1 0 32928 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_296
timestamp 1669390400
transform 1 0 34496 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_307
timestamp 1669390400
transform 1 0 35728 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_311
timestamp 1669390400
transform 1 0 36176 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_317
timestamp 1669390400
transform 1 0 36848 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_321
timestamp 1669390400
transform 1 0 37296 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_328
timestamp 1669390400
transform 1 0 38080 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_332
timestamp 1669390400
transform 1 0 38528 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_336
timestamp 1669390400
transform 1 0 38976 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_341
timestamp 1669390400
transform 1 0 39536 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_354
timestamp 1669390400
transform 1 0 40992 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_358
timestamp 1669390400
transform 1 0 41440 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_362
timestamp 1669390400
transform 1 0 41888 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_372
timestamp 1669390400
transform 1 0 43008 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_383
timestamp 1669390400
transform 1 0 44240 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_387
timestamp 1669390400
transform 1 0 44688 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_389
timestamp 1669390400
transform 1 0 44912 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_392
timestamp 1669390400
transform 1 0 45248 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_395
timestamp 1669390400
transform 1 0 45584 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_410
timestamp 1669390400
transform 1 0 47264 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_420
timestamp 1669390400
transform 1 0 48384 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_424
timestamp 1669390400
transform 1 0 48832 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_428
timestamp 1669390400
transform 1 0 49280 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_442
timestamp 1669390400
transform 1 0 50848 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_446
timestamp 1669390400
transform 1 0 51296 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_450
timestamp 1669390400
transform 1 0 51744 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_58_454
timestamp 1669390400
transform 1 0 52192 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_460
timestamp 1669390400
transform 1 0 52864 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_463
timestamp 1669390400
transform 1 0 53200 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_466
timestamp 1669390400
transform 1 0 53536 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_470
timestamp 1669390400
transform 1 0 53984 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_474
timestamp 1669390400
transform 1 0 54432 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_58_476
timestamp 1669390400
transform 1 0 54656 0 1 48608
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_58_491
timestamp 1669390400
transform 1 0 56336 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_58_507
timestamp 1669390400
transform 1 0 58128 0 1 48608
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_59_2
timestamp 1669390400
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_66
timestamp 1669390400
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_70
timestamp 1669390400
transform 1 0 9184 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_73
timestamp 1669390400
transform 1 0 9520 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_87
timestamp 1669390400
transform 1 0 11088 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_103
timestamp 1669390400
transform 1 0 12880 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_113
timestamp 1669390400
transform 1 0 14000 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_129
timestamp 1669390400
transform 1 0 15792 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_137
timestamp 1669390400
transform 1 0 16688 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_141
timestamp 1669390400
transform 1 0 17136 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_59_144
timestamp 1669390400
transform 1 0 17472 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_160
timestamp 1669390400
transform 1 0 19264 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_164
timestamp 1669390400
transform 1 0 19712 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_167
timestamp 1669390400
transform 1 0 20048 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_182
timestamp 1669390400
transform 1 0 21728 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_184
timestamp 1669390400
transform 1 0 21952 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_191
timestamp 1669390400
transform 1 0 22736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_206
timestamp 1669390400
transform 1 0 24416 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_210
timestamp 1669390400
transform 1 0 24864 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_212
timestamp 1669390400
transform 1 0 25088 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_215
timestamp 1669390400
transform 1 0 25424 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_233
timestamp 1669390400
transform 1 0 27440 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_243
timestamp 1669390400
transform 1 0 28560 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_247
timestamp 1669390400
transform 1 0 29008 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_272
timestamp 1669390400
transform 1 0 31808 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_276
timestamp 1669390400
transform 1 0 32256 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_280
timestamp 1669390400
transform 1 0 32704 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_286
timestamp 1669390400
transform 1 0 33376 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_295
timestamp 1669390400
transform 1 0 34384 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_303
timestamp 1669390400
transform 1 0 35280 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_315
timestamp 1669390400
transform 1 0 36624 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_319
timestamp 1669390400
transform 1 0 37072 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_323
timestamp 1669390400
transform 1 0 37520 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_331
timestamp 1669390400
transform 1 0 38416 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_333
timestamp 1669390400
transform 1 0 38640 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_336
timestamp 1669390400
transform 1 0 38976 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_340
timestamp 1669390400
transform 1 0 39424 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_354
timestamp 1669390400
transform 1 0 40992 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_357
timestamp 1669390400
transform 1 0 41328 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_360
timestamp 1669390400
transform 1 0 41664 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_368
timestamp 1669390400
transform 1 0 42560 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_372
timestamp 1669390400
transform 1 0 43008 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_384
timestamp 1669390400
transform 1 0 44352 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_388
timestamp 1669390400
transform 1 0 44800 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_392
timestamp 1669390400
transform 1 0 45248 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_396
timestamp 1669390400
transform 1 0 45696 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_408
timestamp 1669390400
transform 1 0 47040 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_414
timestamp 1669390400
transform 1 0 47712 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_418
timestamp 1669390400
transform 1 0 48160 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_420
timestamp 1669390400
transform 1 0 48384 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_423
timestamp 1669390400
transform 1 0 48720 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_425
timestamp 1669390400
transform 1 0 48944 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_59_428
timestamp 1669390400
transform 1 0 49280 0 -1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_431
timestamp 1669390400
transform 1 0 49616 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_435
timestamp 1669390400
transform 1 0 50064 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_439
timestamp 1669390400
transform 1 0 50512 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_443
timestamp 1669390400
transform 1 0 50960 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_447
timestamp 1669390400
transform 1 0 51408 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_453
timestamp 1669390400
transform 1 0 52080 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_457
timestamp 1669390400
transform 1 0 52528 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_461
timestamp 1669390400
transform 1 0 52976 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_465
timestamp 1669390400
transform 1 0 53424 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_469
timestamp 1669390400
transform 1 0 53872 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_473
timestamp 1669390400
transform 1 0 54320 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_477
timestamp 1669390400
transform 1 0 54768 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_481
timestamp 1669390400
transform 1 0 55216 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_485
timestamp 1669390400
transform 1 0 55664 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_59_493
timestamp 1669390400
transform 1 0 56560 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_59_499
timestamp 1669390400
transform 1 0 57232 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_59_507
timestamp 1669390400
transform 1 0 58128 0 -1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_2
timestamp 1669390400
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_34
timestamp 1669390400
transform 1 0 5152 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_37
timestamp 1669390400
transform 1 0 5488 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_53
timestamp 1669390400
transform 1 0 7280 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_61
timestamp 1669390400
transform 1 0 8176 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_65
timestamp 1669390400
transform 1 0 8624 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_72
timestamp 1669390400
transform 1 0 9408 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_104
timestamp 1669390400
transform 1 0 12992 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_60_108
timestamp 1669390400
transform 1 0 13440 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_172
timestamp 1669390400
transform 1 0 20608 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_176
timestamp 1669390400
transform 1 0 21056 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_179
timestamp 1669390400
transform 1 0 21392 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_193
timestamp 1669390400
transform 1 0 22960 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_197
timestamp 1669390400
transform 1 0 23408 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_199
timestamp 1669390400
transform 1 0 23632 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_213
timestamp 1669390400
transform 1 0 25200 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_217
timestamp 1669390400
transform 1 0 25648 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_231
timestamp 1669390400
transform 1 0 27216 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_235
timestamp 1669390400
transform 1 0 27664 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_243
timestamp 1669390400
transform 1 0 28560 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_247
timestamp 1669390400
transform 1 0 29008 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_60_250
timestamp 1669390400
transform 1 0 29344 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_266
timestamp 1669390400
transform 1 0 31136 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_270
timestamp 1669390400
transform 1 0 31584 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_274
timestamp 1669390400
transform 1 0 32032 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_284
timestamp 1669390400
transform 1 0 33152 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_288
timestamp 1669390400
transform 1 0 33600 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_296
timestamp 1669390400
transform 1 0 34496 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_300
timestamp 1669390400
transform 1 0 34944 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_304
timestamp 1669390400
transform 1 0 35392 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_318
timestamp 1669390400
transform 1 0 36960 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_321
timestamp 1669390400
transform 1 0 37296 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_324
timestamp 1669390400
transform 1 0 37632 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_328
timestamp 1669390400
transform 1 0 38080 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_332
timestamp 1669390400
transform 1 0 38528 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_340
timestamp 1669390400
transform 1 0 39424 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_348
timestamp 1669390400
transform 1 0 40320 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_356
timestamp 1669390400
transform 1 0 41216 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_360
timestamp 1669390400
transform 1 0 41664 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_364
timestamp 1669390400
transform 1 0 42112 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_389
timestamp 1669390400
transform 1 0 44912 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_392
timestamp 1669390400
transform 1 0 45248 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_398
timestamp 1669390400
transform 1 0 45920 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_402
timestamp 1669390400
transform 1 0 46368 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_404
timestamp 1669390400
transform 1 0 46592 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_411
timestamp 1669390400
transform 1 0 47376 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_413
timestamp 1669390400
transform 1 0 47600 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_416
timestamp 1669390400
transform 1 0 47936 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_420
timestamp 1669390400
transform 1 0 48384 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_424
timestamp 1669390400
transform 1 0 48832 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_434
timestamp 1669390400
transform 1 0 49952 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_440
timestamp 1669390400
transform 1 0 50624 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_444
timestamp 1669390400
transform 1 0 51072 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_448
timestamp 1669390400
transform 1 0 51520 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_454
timestamp 1669390400
transform 1 0 52192 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_458
timestamp 1669390400
transform 1 0 52640 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_60_460
timestamp 1669390400
transform 1 0 52864 0 1 50176
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_60_463
timestamp 1669390400
transform 1 0 53200 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_60_495
timestamp 1669390400
transform 1 0 56784 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_60_503
timestamp 1669390400
transform 1 0 57680 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_60_507
timestamp 1669390400
transform 1 0 58128 0 1 50176
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_2
timestamp 1669390400
transform 1 0 1568 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_66
timestamp 1669390400
transform 1 0 8736 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_70
timestamp 1669390400
transform 1 0 9184 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_61_73
timestamp 1669390400
transform 1 0 9520 0 -1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_137
timestamp 1669390400
transform 1 0 16688 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_141
timestamp 1669390400
transform 1 0 17136 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_144
timestamp 1669390400
transform 1 0 17472 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_176
timestamp 1669390400
transform 1 0 21056 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_180
timestamp 1669390400
transform 1 0 21504 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_184
timestamp 1669390400
transform 1 0 21952 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_192
timestamp 1669390400
transform 1 0 22848 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_204
timestamp 1669390400
transform 1 0 24192 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_211
timestamp 1669390400
transform 1 0 24976 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_215
timestamp 1669390400
transform 1 0 25424 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_219
timestamp 1669390400
transform 1 0 25872 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_226
timestamp 1669390400
transform 1 0 26656 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_240
timestamp 1669390400
transform 1 0 28224 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_256
timestamp 1669390400
transform 1 0 30016 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_264
timestamp 1669390400
transform 1 0 30912 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_268
timestamp 1669390400
transform 1 0 31360 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_283
timestamp 1669390400
transform 1 0 33040 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_286
timestamp 1669390400
transform 1 0 33376 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_299
timestamp 1669390400
transform 1 0 34832 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_301
timestamp 1669390400
transform 1 0 35056 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_326
timestamp 1669390400
transform 1 0 37856 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_336
timestamp 1669390400
transform 1 0 38976 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_340
timestamp 1669390400
transform 1 0 39424 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_344
timestamp 1669390400
transform 1 0 39872 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_351
timestamp 1669390400
transform 1 0 40656 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_357
timestamp 1669390400
transform 1 0 41328 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_360
timestamp 1669390400
transform 1 0 41664 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_364
timestamp 1669390400
transform 1 0 42112 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_370
timestamp 1669390400
transform 1 0 42784 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_383
timestamp 1669390400
transform 1 0 44240 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_389
timestamp 1669390400
transform 1 0 44912 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_393
timestamp 1669390400
transform 1 0 45360 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_397
timestamp 1669390400
transform 1 0 45808 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_401
timestamp 1669390400
transform 1 0 46256 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_405
timestamp 1669390400
transform 1 0 46704 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_420
timestamp 1669390400
transform 1 0 48384 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_424
timestamp 1669390400
transform 1 0 48832 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_428
timestamp 1669390400
transform 1 0 49280 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_437
timestamp 1669390400
transform 1 0 50288 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_439
timestamp 1669390400
transform 1 0 50512 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_61_442
timestamp 1669390400
transform 1 0 50848 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_61_474
timestamp 1669390400
transform 1 0 54432 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_61_490
timestamp 1669390400
transform 1 0 56224 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_494
timestamp 1669390400
transform 1 0 56672 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_61_496
timestamp 1669390400
transform 1 0 56896 0 -1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_61_499
timestamp 1669390400
transform 1 0 57232 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_61_507
timestamp 1669390400
transform 1 0 58128 0 -1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_2
timestamp 1669390400
transform 1 0 1568 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_17
timestamp 1669390400
transform 1 0 3248 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_33
timestamp 1669390400
transform 1 0 5040 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_37
timestamp 1669390400
transform 1 0 5488 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_101
timestamp 1669390400
transform 1 0 12656 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_105
timestamp 1669390400
transform 1 0 13104 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_62_108
timestamp 1669390400
transform 1 0 13440 0 1 51744
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_172
timestamp 1669390400
transform 1 0 20608 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_176
timestamp 1669390400
transform 1 0 21056 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_179
timestamp 1669390400
transform 1 0 21392 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_211
timestamp 1669390400
transform 1 0 24976 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_219
timestamp 1669390400
transform 1 0 25872 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_223
timestamp 1669390400
transform 1 0 26320 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_225
timestamp 1669390400
transform 1 0 26544 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_228
timestamp 1669390400
transform 1 0 26880 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_244
timestamp 1669390400
transform 1 0 28672 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_62_250
timestamp 1669390400
transform 1 0 29344 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_266
timestamp 1669390400
transform 1 0 31136 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_274
timestamp 1669390400
transform 1 0 32032 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_276
timestamp 1669390400
transform 1 0 32256 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_293
timestamp 1669390400
transform 1 0 34160 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_303
timestamp 1669390400
transform 1 0 35280 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_318
timestamp 1669390400
transform 1 0 36960 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_321
timestamp 1669390400
transform 1 0 37296 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_324
timestamp 1669390400
transform 1 0 37632 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_328
timestamp 1669390400
transform 1 0 38080 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_332
timestamp 1669390400
transform 1 0 38528 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_347
timestamp 1669390400
transform 1 0 40208 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_351
timestamp 1669390400
transform 1 0 40656 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_355
timestamp 1669390400
transform 1 0 41104 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_359
timestamp 1669390400
transform 1 0 41552 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_372
timestamp 1669390400
transform 1 0 43008 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_386
timestamp 1669390400
transform 1 0 44576 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_392
timestamp 1669390400
transform 1 0 45248 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_395
timestamp 1669390400
transform 1 0 45584 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_62_397
timestamp 1669390400
transform 1 0 45808 0 1 51744
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_405
timestamp 1669390400
transform 1 0 46704 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_417
timestamp 1669390400
transform 1 0 48048 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_421
timestamp 1669390400
transform 1 0 48496 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_425
timestamp 1669390400
transform 1 0 48944 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_429
timestamp 1669390400
transform 1 0 49392 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_62_463
timestamp 1669390400
transform 1 0 53200 0 1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_62_495
timestamp 1669390400
transform 1 0 56784 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_62_503
timestamp 1669390400
transform 1 0 57680 0 1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_62_507
timestamp 1669390400
transform 1 0 58128 0 1 51744
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_2
timestamp 1669390400
transform 1 0 1568 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_66
timestamp 1669390400
transform 1 0 8736 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_70
timestamp 1669390400
transform 1 0 9184 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_73
timestamp 1669390400
transform 1 0 9520 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_137
timestamp 1669390400
transform 1 0 16688 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_141
timestamp 1669390400
transform 1 0 17136 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_144
timestamp 1669390400
transform 1 0 17472 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_208
timestamp 1669390400
transform 1 0 24640 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_212
timestamp 1669390400
transform 1 0 25088 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_215
timestamp 1669390400
transform 1 0 25424 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_279
timestamp 1669390400
transform 1 0 32592 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_283
timestamp 1669390400
transform 1 0 33040 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_286
timestamp 1669390400
transform 1 0 33376 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_295
timestamp 1669390400
transform 1 0 34384 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_299
timestamp 1669390400
transform 1 0 34832 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_303
timestamp 1669390400
transform 1 0 35280 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_307
timestamp 1669390400
transform 1 0 35728 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_311
timestamp 1669390400
transform 1 0 36176 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_315
timestamp 1669390400
transform 1 0 36624 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_323
timestamp 1669390400
transform 1 0 37520 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_327
timestamp 1669390400
transform 1 0 37968 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_329
timestamp 1669390400
transform 1 0 38192 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_332
timestamp 1669390400
transform 1 0 38528 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_340
timestamp 1669390400
transform 1 0 39424 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_344
timestamp 1669390400
transform 1 0 39872 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_348
timestamp 1669390400
transform 1 0 40320 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_354
timestamp 1669390400
transform 1 0 40992 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_357
timestamp 1669390400
transform 1 0 41328 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_365
timestamp 1669390400
transform 1 0 42224 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_374
timestamp 1669390400
transform 1 0 43232 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_387
timestamp 1669390400
transform 1 0 44688 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_391
timestamp 1669390400
transform 1 0 45136 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_399
timestamp 1669390400
transform 1 0 46032 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_403
timestamp 1669390400
transform 1 0 46480 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_413
timestamp 1669390400
transform 1 0 47600 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_417
timestamp 1669390400
transform 1 0 48048 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_425
timestamp 1669390400
transform 1 0 48944 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_63_428
timestamp 1669390400
transform 1 0 49280 0 -1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_63_492
timestamp 1669390400
transform 1 0 56448 0 -1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_63_496
timestamp 1669390400
transform 1 0 56896 0 -1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_63_499
timestamp 1669390400
transform 1 0 57232 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_63_507
timestamp 1669390400
transform 1 0 58128 0 -1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_2
timestamp 1669390400
transform 1 0 1568 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_6
timestamp 1669390400
transform 1 0 2016 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_14
timestamp 1669390400
transform 1 0 2912 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_64_18
timestamp 1669390400
transform 1 0 3360 0 1 53312
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_34
timestamp 1669390400
transform 1 0 5152 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_37
timestamp 1669390400
transform 1 0 5488 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_101
timestamp 1669390400
transform 1 0 12656 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_105
timestamp 1669390400
transform 1 0 13104 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_108
timestamp 1669390400
transform 1 0 13440 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_172
timestamp 1669390400
transform 1 0 20608 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_176
timestamp 1669390400
transform 1 0 21056 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_179
timestamp 1669390400
transform 1 0 21392 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_243
timestamp 1669390400
transform 1 0 28560 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_247
timestamp 1669390400
transform 1 0 29008 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_250
timestamp 1669390400
transform 1 0 29344 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_314
timestamp 1669390400
transform 1 0 36512 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_318
timestamp 1669390400
transform 1 0 36960 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_321
timestamp 1669390400
transform 1 0 37296 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_329
timestamp 1669390400
transform 1 0 38192 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_333
timestamp 1669390400
transform 1 0 38640 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_340
timestamp 1669390400
transform 1 0 39424 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_344
timestamp 1669390400
transform 1 0 39872 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_363
timestamp 1669390400
transform 1 0 42000 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_365
timestamp 1669390400
transform 1 0 42224 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_368
timestamp 1669390400
transform 1 0 42560 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_377
timestamp 1669390400
transform 1 0 43568 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_381
timestamp 1669390400
transform 1 0 44016 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_385
timestamp 1669390400
transform 1 0 44464 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_389
timestamp 1669390400
transform 1 0 44912 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_64_392
timestamp 1669390400
transform 1 0 45248 0 1 53312
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_456
timestamp 1669390400
transform 1 0 52416 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_64_460
timestamp 1669390400
transform 1 0 52864 0 1 53312
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_64_463
timestamp 1669390400
transform 1 0 53200 0 1 53312
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_64_495
timestamp 1669390400
transform 1 0 56784 0 1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_64_503
timestamp 1669390400
transform 1 0 57680 0 1 53312
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_64_507
timestamp 1669390400
transform 1 0 58128 0 1 53312
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_2
timestamp 1669390400
transform 1 0 1568 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_66
timestamp 1669390400
transform 1 0 8736 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_70
timestamp 1669390400
transform 1 0 9184 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_73
timestamp 1669390400
transform 1 0 9520 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_137
timestamp 1669390400
transform 1 0 16688 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_141
timestamp 1669390400
transform 1 0 17136 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_144
timestamp 1669390400
transform 1 0 17472 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_208
timestamp 1669390400
transform 1 0 24640 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_212
timestamp 1669390400
transform 1 0 25088 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_215
timestamp 1669390400
transform 1 0 25424 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_279
timestamp 1669390400
transform 1 0 32592 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_283
timestamp 1669390400
transform 1 0 33040 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_286
timestamp 1669390400
transform 1 0 33376 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_318
timestamp 1669390400
transform 1 0 36960 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_334
timestamp 1669390400
transform 1 0 38752 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_344
timestamp 1669390400
transform 1 0 39872 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_354
timestamp 1669390400
transform 1 0 40992 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_357
timestamp 1669390400
transform 1 0 41328 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_361
timestamp 1669390400
transform 1 0 41776 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_371
timestamp 1669390400
transform 1 0 42896 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_65_383
timestamp 1669390400
transform 1 0 44240 0 -1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_415
timestamp 1669390400
transform 1 0 47824 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_423
timestamp 1669390400
transform 1 0 48720 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_425
timestamp 1669390400
transform 1 0 48944 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_65_428
timestamp 1669390400
transform 1 0 49280 0 -1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_65_492
timestamp 1669390400
transform 1 0 56448 0 -1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_65_496
timestamp 1669390400
transform 1 0 56896 0 -1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_65_499
timestamp 1669390400
transform 1 0 57232 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_65_507
timestamp 1669390400
transform 1 0 58128 0 -1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_2
timestamp 1669390400
transform 1 0 1568 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_17
timestamp 1669390400
transform 1 0 3248 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_21
timestamp 1669390400
transform 1 0 3696 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_29
timestamp 1669390400
transform 1 0 4592 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_33
timestamp 1669390400
transform 1 0 5040 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_37
timestamp 1669390400
transform 1 0 5488 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_101
timestamp 1669390400
transform 1 0 12656 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_105
timestamp 1669390400
transform 1 0 13104 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_66_108
timestamp 1669390400
transform 1 0 13440 0 1 54880
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_172
timestamp 1669390400
transform 1 0 20608 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_176
timestamp 1669390400
transform 1 0 21056 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_179
timestamp 1669390400
transform 1 0 21392 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_187
timestamp 1669390400
transform 1 0 22288 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_193
timestamp 1669390400
transform 1 0 22960 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_201
timestamp 1669390400
transform 1 0 23856 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_217
timestamp 1669390400
transform 1 0 25648 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_225
timestamp 1669390400
transform 1 0 26544 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_232
timestamp 1669390400
transform 1 0 27328 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_250
timestamp 1669390400
transform 1 0 29344 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_257
timestamp 1669390400
transform 1 0 30128 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_265
timestamp 1669390400
transform 1 0 31024 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_269
timestamp 1669390400
transform 1 0 31472 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_296
timestamp 1669390400
transform 1 0 34496 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_312
timestamp 1669390400
transform 1 0 36288 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_316
timestamp 1669390400
transform 1 0 36736 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_318
timestamp 1669390400
transform 1 0 36960 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_321
timestamp 1669390400
transform 1 0 37296 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_328
timestamp 1669390400
transform 1 0 38080 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_336
timestamp 1669390400
transform 1 0 38976 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_350
timestamp 1669390400
transform 1 0 40544 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_358
timestamp 1669390400
transform 1 0 41440 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_360
timestamp 1669390400
transform 1 0 41664 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_384
timestamp 1669390400
transform 1 0 44352 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_388
timestamp 1669390400
transform 1 0 44800 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_392
timestamp 1669390400
transform 1 0 45248 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_400
timestamp 1669390400
transform 1 0 46144 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_66_402
timestamp 1669390400
transform 1 0 46368 0 1 54880
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_66_409
timestamp 1669390400
transform 1 0 47152 0 1 54880
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_66_441
timestamp 1669390400
transform 1 0 50736 0 1 54880
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_457
timestamp 1669390400
transform 1 0 52528 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_463
timestamp 1669390400
transform 1 0 53200 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_471
timestamp 1669390400
transform 1 0 54096 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_475
timestamp 1669390400
transform 1 0 54544 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_491
timestamp 1669390400
transform 1 0 56336 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_66_495
timestamp 1669390400
transform 1 0 56784 0 1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_66_503
timestamp 1669390400
transform 1 0 57680 0 1 54880
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_66_507
timestamp 1669390400
transform 1 0 58128 0 1 54880
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_2
timestamp 1669390400
transform 1 0 1568 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_10
timestamp 1669390400
transform 1 0 2464 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_12
timestamp 1669390400
transform 1 0 2688 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_27
timestamp 1669390400
transform 1 0 4368 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_31
timestamp 1669390400
transform 1 0 4816 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_37
timestamp 1669390400
transform 1 0 5488 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_53
timestamp 1669390400
transform 1 0 7280 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_69
timestamp 1669390400
transform 1 0 9072 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_72
timestamp 1669390400
transform 1 0 9408 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_104
timestamp 1669390400
transform 1 0 12992 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_107
timestamp 1669390400
transform 1 0 13328 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_113
timestamp 1669390400
transform 1 0 14000 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_129
timestamp 1669390400
transform 1 0 15792 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_137
timestamp 1669390400
transform 1 0 16688 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_139
timestamp 1669390400
transform 1 0 16912 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_142
timestamp 1669390400
transform 1 0 17248 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_158
timestamp 1669390400
transform 1 0 19040 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_174
timestamp 1669390400
transform 1 0 20832 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_177
timestamp 1669390400
transform 1 0 21168 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_180
timestamp 1669390400
transform 1 0 21504 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_196
timestamp 1669390400
transform 1 0 23296 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_204
timestamp 1669390400
transform 1 0 24192 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_208
timestamp 1669390400
transform 1 0 24640 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_212
timestamp 1669390400
transform 1 0 25088 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_216
timestamp 1669390400
transform 1 0 25536 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_231
timestamp 1669390400
transform 1 0 27216 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_235
timestamp 1669390400
transform 1 0 27664 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_243
timestamp 1669390400
transform 1 0 28560 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_247
timestamp 1669390400
transform 1 0 29008 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_279
timestamp 1669390400
transform 1 0 32592 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_282
timestamp 1669390400
transform 1 0 32928 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_298
timestamp 1669390400
transform 1 0 34720 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_306
timestamp 1669390400
transform 1 0 35616 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_310
timestamp 1669390400
transform 1 0 36064 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_314
timestamp 1669390400
transform 1 0 36512 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_317
timestamp 1669390400
transform 1 0 36848 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_333
timestamp 1669390400
transform 1 0 38640 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_349
timestamp 1669390400
transform 1 0 40432 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_352
timestamp 1669390400
transform 1 0 40768 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_361
timestamp 1669390400
transform 1 0 41776 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_365
timestamp 1669390400
transform 1 0 42224 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_368
timestamp 1669390400
transform 1 0 42560 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_384
timestamp 1669390400
transform 1 0 44352 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_67_387
timestamp 1669390400
transform 1 0 44688 0 -1 56448
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_419
timestamp 1669390400
transform 1 0 48272 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_422
timestamp 1669390400
transform 1 0 48608 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_67_437
timestamp 1669390400
transform 1 0 50288 0 -1 56448
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_453
timestamp 1669390400
transform 1 0 52080 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_67_457
timestamp 1669390400
transform 1 0 52528 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_67_465
timestamp 1669390400
transform 1 0 53424 0 -1 56448
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_469
timestamp 1669390400
transform 1 0 53872 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_473
timestamp 1669390400
transform 1 0 54320 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_489
timestamp 1669390400
transform 1 0 56112 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_67_492
timestamp 1669390400
transform 1 0 56448 0 -1 56448
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_67_507
timestamp 1669390400
transform 1 0 58128 0 -1 56448
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1669390400
transform -1 0 58576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1669390400
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1669390400
transform -1 0 58576 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1669390400
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1669390400
transform -1 0 58576 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1669390400
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1669390400
transform -1 0 58576 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1669390400
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1669390400
transform -1 0 58576 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1669390400
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1669390400
transform -1 0 58576 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1669390400
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1669390400
transform -1 0 58576 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1669390400
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1669390400
transform -1 0 58576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1669390400
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1669390400
transform -1 0 58576 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1669390400
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1669390400
transform -1 0 58576 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1669390400
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1669390400
transform -1 0 58576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1669390400
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1669390400
transform -1 0 58576 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1669390400
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1669390400
transform -1 0 58576 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1669390400
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1669390400
transform -1 0 58576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1669390400
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1669390400
transform -1 0 58576 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1669390400
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1669390400
transform -1 0 58576 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1669390400
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1669390400
transform -1 0 58576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1669390400
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1669390400
transform -1 0 58576 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1669390400
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1669390400
transform -1 0 58576 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1669390400
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1669390400
transform -1 0 58576 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1669390400
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1669390400
transform -1 0 58576 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1669390400
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1669390400
transform -1 0 58576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1669390400
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1669390400
transform -1 0 58576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1669390400
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1669390400
transform -1 0 58576 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1669390400
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1669390400
transform -1 0 58576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1669390400
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1669390400
transform -1 0 58576 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1669390400
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1669390400
transform -1 0 58576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1669390400
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1669390400
transform -1 0 58576 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1669390400
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1669390400
transform -1 0 58576 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1669390400
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1669390400
transform -1 0 58576 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1669390400
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1669390400
transform -1 0 58576 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1669390400
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1669390400
transform -1 0 58576 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1669390400
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1669390400
transform -1 0 58576 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1669390400
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1669390400
transform -1 0 58576 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1669390400
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1669390400
transform -1 0 58576 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1669390400
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1669390400
transform -1 0 58576 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1669390400
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1669390400
transform -1 0 58576 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1669390400
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1669390400
transform -1 0 58576 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1669390400
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1669390400
transform -1 0 58576 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1669390400
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1669390400
transform -1 0 58576 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1669390400
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1669390400
transform -1 0 58576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1669390400
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1669390400
transform -1 0 58576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1669390400
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1669390400
transform -1 0 58576 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1669390400
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1669390400
transform -1 0 58576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1669390400
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1669390400
transform -1 0 58576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1669390400
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1669390400
transform -1 0 58576 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1669390400
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1669390400
transform -1 0 58576 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1669390400
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1669390400
transform -1 0 58576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1669390400
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1669390400
transform -1 0 58576 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1669390400
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1669390400
transform -1 0 58576 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1669390400
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1669390400
transform -1 0 58576 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1669390400
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1669390400
transform -1 0 58576 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1669390400
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1669390400
transform -1 0 58576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1669390400
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1669390400
transform -1 0 58576 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1669390400
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1669390400
transform -1 0 58576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_110
timestamp 1669390400
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_111
timestamp 1669390400
transform -1 0 58576 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_112
timestamp 1669390400
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_113
timestamp 1669390400
transform -1 0 58576 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_114
timestamp 1669390400
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_115
timestamp 1669390400
transform -1 0 58576 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_116
timestamp 1669390400
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_117
timestamp 1669390400
transform -1 0 58576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_118
timestamp 1669390400
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_119
timestamp 1669390400
transform -1 0 58576 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_120
timestamp 1669390400
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_121
timestamp 1669390400
transform -1 0 58576 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_122
timestamp 1669390400
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_123
timestamp 1669390400
transform -1 0 58576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_124
timestamp 1669390400
transform 1 0 1344 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_125
timestamp 1669390400
transform -1 0 58576 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_126
timestamp 1669390400
transform 1 0 1344 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_127
timestamp 1669390400
transform -1 0 58576 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_128
timestamp 1669390400
transform 1 0 1344 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_129
timestamp 1669390400
transform -1 0 58576 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_130
timestamp 1669390400
transform 1 0 1344 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_131
timestamp 1669390400
transform -1 0 58576 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_132
timestamp 1669390400
transform 1 0 1344 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_133
timestamp 1669390400
transform -1 0 58576 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_134
timestamp 1669390400
transform 1 0 1344 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_135
timestamp 1669390400
transform -1 0 58576 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1669390400
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1669390400
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1669390400
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1669390400
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1669390400
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1669390400
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1669390400
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1669390400
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1669390400
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1669390400
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1669390400
transform 1 0 48384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1669390400
transform 1 0 52304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1669390400
transform 1 0 56224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1669390400
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1669390400
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1669390400
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1669390400
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1669390400
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1669390400
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1669390400
transform 1 0 57008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1669390400
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1669390400
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1669390400
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1669390400
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1669390400
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1669390400
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1669390400
transform 1 0 52976 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1669390400
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1669390400
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1669390400
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1669390400
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1669390400
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1669390400
transform 1 0 49056 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1669390400
transform 1 0 57008 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1669390400
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1669390400
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1669390400
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1669390400
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1669390400
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1669390400
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1669390400
transform 1 0 52976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1669390400
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1669390400
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1669390400
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1669390400
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1669390400
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1669390400
transform 1 0 49056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1669390400
transform 1 0 57008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1669390400
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1669390400
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1669390400
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1669390400
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1669390400
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1669390400
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1669390400
transform 1 0 52976 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1669390400
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1669390400
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1669390400
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1669390400
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1669390400
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1669390400
transform 1 0 49056 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1669390400
transform 1 0 57008 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1669390400
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1669390400
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1669390400
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1669390400
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1669390400
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1669390400
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1669390400
transform 1 0 52976 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1669390400
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1669390400
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1669390400
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1669390400
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1669390400
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1669390400
transform 1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1669390400
transform 1 0 57008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1669390400
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1669390400
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1669390400
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1669390400
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1669390400
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1669390400
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1669390400
transform 1 0 52976 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1669390400
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1669390400
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1669390400
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1669390400
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1669390400
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1669390400
transform 1 0 49056 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1669390400
transform 1 0 57008 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1669390400
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1669390400
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1669390400
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1669390400
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1669390400
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1669390400
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1669390400
transform 1 0 52976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1669390400
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1669390400
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1669390400
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1669390400
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1669390400
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1669390400
transform 1 0 49056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1669390400
transform 1 0 57008 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1669390400
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1669390400
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1669390400
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1669390400
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1669390400
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1669390400
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1669390400
transform 1 0 52976 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1669390400
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1669390400
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1669390400
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1669390400
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1669390400
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1669390400
transform 1 0 49056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1669390400
transform 1 0 57008 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1669390400
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1669390400
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1669390400
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1669390400
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1669390400
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1669390400
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1669390400
transform 1 0 52976 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1669390400
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1669390400
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1669390400
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1669390400
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1669390400
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1669390400
transform 1 0 49056 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1669390400
transform 1 0 57008 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1669390400
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1669390400
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1669390400
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1669390400
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1669390400
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1669390400
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1669390400
transform 1 0 52976 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1669390400
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1669390400
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1669390400
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1669390400
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1669390400
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1669390400
transform 1 0 49056 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1669390400
transform 1 0 57008 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1669390400
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1669390400
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1669390400
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1669390400
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1669390400
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1669390400
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1669390400
transform 1 0 52976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1669390400
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1669390400
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1669390400
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1669390400
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1669390400
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1669390400
transform 1 0 49056 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1669390400
transform 1 0 57008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1669390400
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1669390400
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1669390400
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1669390400
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1669390400
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1669390400
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1669390400
transform 1 0 52976 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1669390400
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1669390400
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1669390400
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1669390400
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1669390400
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1669390400
transform 1 0 49056 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1669390400
transform 1 0 57008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1669390400
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1669390400
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1669390400
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1669390400
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1669390400
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1669390400
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1669390400
transform 1 0 52976 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1669390400
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1669390400
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1669390400
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1669390400
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1669390400
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1669390400
transform 1 0 49056 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1669390400
transform 1 0 57008 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1669390400
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1669390400
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1669390400
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1669390400
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1669390400
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1669390400
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1669390400
transform 1 0 52976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1669390400
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1669390400
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1669390400
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1669390400
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1669390400
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1669390400
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1669390400
transform 1 0 57008 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1669390400
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1669390400
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1669390400
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1669390400
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1669390400
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1669390400
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1669390400
transform 1 0 52976 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1669390400
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1669390400
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1669390400
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1669390400
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1669390400
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1669390400
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1669390400
transform 1 0 57008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1669390400
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1669390400
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1669390400
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1669390400
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1669390400
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1669390400
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1669390400
transform 1 0 52976 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1669390400
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1669390400
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1669390400
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1669390400
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1669390400
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1669390400
transform 1 0 49056 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1669390400
transform 1 0 57008 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1669390400
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1669390400
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1669390400
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1669390400
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1669390400
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1669390400
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1669390400
transform 1 0 52976 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1669390400
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1669390400
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1669390400
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1669390400
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1669390400
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1669390400
transform 1 0 49056 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1669390400
transform 1 0 57008 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1669390400
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1669390400
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1669390400
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1669390400
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1669390400
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1669390400
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1669390400
transform 1 0 52976 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1669390400
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1669390400
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1669390400
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1669390400
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1669390400
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1669390400
transform 1 0 49056 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1669390400
transform 1 0 57008 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1669390400
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1669390400
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1669390400
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1669390400
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1669390400
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1669390400
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1669390400
transform 1 0 52976 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1669390400
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1669390400
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1669390400
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1669390400
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1669390400
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1669390400
transform 1 0 49056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1669390400
transform 1 0 57008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1669390400
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1669390400
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1669390400
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1669390400
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1669390400
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1669390400
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1669390400
transform 1 0 52976 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1669390400
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1669390400
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1669390400
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1669390400
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1669390400
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1669390400
transform 1 0 49056 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1669390400
transform 1 0 57008 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_423
timestamp 1669390400
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_424
timestamp 1669390400
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_425
timestamp 1669390400
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_426
timestamp 1669390400
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_427
timestamp 1669390400
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_428
timestamp 1669390400
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_429
timestamp 1669390400
transform 1 0 52976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_430
timestamp 1669390400
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_431
timestamp 1669390400
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_432
timestamp 1669390400
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_433
timestamp 1669390400
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_434
timestamp 1669390400
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_435
timestamp 1669390400
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_436
timestamp 1669390400
transform 1 0 57008 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_437
timestamp 1669390400
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_438
timestamp 1669390400
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_439
timestamp 1669390400
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_440
timestamp 1669390400
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_441
timestamp 1669390400
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_442
timestamp 1669390400
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_443
timestamp 1669390400
transform 1 0 52976 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_444
timestamp 1669390400
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_445
timestamp 1669390400
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_446
timestamp 1669390400
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_447
timestamp 1669390400
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_448
timestamp 1669390400
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_449
timestamp 1669390400
transform 1 0 49056 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_450
timestamp 1669390400
transform 1 0 57008 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_451
timestamp 1669390400
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_452
timestamp 1669390400
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_453
timestamp 1669390400
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_454
timestamp 1669390400
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_455
timestamp 1669390400
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_456
timestamp 1669390400
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_457
timestamp 1669390400
transform 1 0 52976 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_458
timestamp 1669390400
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_459
timestamp 1669390400
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_460
timestamp 1669390400
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_461
timestamp 1669390400
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_462
timestamp 1669390400
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_463
timestamp 1669390400
transform 1 0 49056 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_464
timestamp 1669390400
transform 1 0 57008 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_465
timestamp 1669390400
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_466
timestamp 1669390400
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_467
timestamp 1669390400
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_468
timestamp 1669390400
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_469
timestamp 1669390400
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_470
timestamp 1669390400
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_471
timestamp 1669390400
transform 1 0 52976 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_472
timestamp 1669390400
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_473
timestamp 1669390400
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_474
timestamp 1669390400
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_475
timestamp 1669390400
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_476
timestamp 1669390400
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_477
timestamp 1669390400
transform 1 0 49056 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_478
timestamp 1669390400
transform 1 0 57008 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_479
timestamp 1669390400
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_480
timestamp 1669390400
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_481
timestamp 1669390400
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_482
timestamp 1669390400
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_483
timestamp 1669390400
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_484
timestamp 1669390400
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_485
timestamp 1669390400
transform 1 0 52976 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_486
timestamp 1669390400
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_487
timestamp 1669390400
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_488
timestamp 1669390400
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_489
timestamp 1669390400
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_490
timestamp 1669390400
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_491
timestamp 1669390400
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_492
timestamp 1669390400
transform 1 0 57008 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_493
timestamp 1669390400
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_494
timestamp 1669390400
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_495
timestamp 1669390400
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_496
timestamp 1669390400
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_497
timestamp 1669390400
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_498
timestamp 1669390400
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_499
timestamp 1669390400
transform 1 0 52976 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_500
timestamp 1669390400
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_501
timestamp 1669390400
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_502
timestamp 1669390400
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_503
timestamp 1669390400
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_504
timestamp 1669390400
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_505
timestamp 1669390400
transform 1 0 49056 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_506
timestamp 1669390400
transform 1 0 57008 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_507
timestamp 1669390400
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_508
timestamp 1669390400
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_509
timestamp 1669390400
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_510
timestamp 1669390400
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_511
timestamp 1669390400
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_512
timestamp 1669390400
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_513
timestamp 1669390400
transform 1 0 52976 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_514
timestamp 1669390400
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_515
timestamp 1669390400
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_516
timestamp 1669390400
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_517
timestamp 1669390400
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_518
timestamp 1669390400
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_519
timestamp 1669390400
transform 1 0 49056 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_520
timestamp 1669390400
transform 1 0 57008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_521
timestamp 1669390400
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_522
timestamp 1669390400
transform 1 0 13216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_523
timestamp 1669390400
transform 1 0 21168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_524
timestamp 1669390400
transform 1 0 29120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_525
timestamp 1669390400
transform 1 0 37072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_526
timestamp 1669390400
transform 1 0 45024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_527
timestamp 1669390400
transform 1 0 52976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_528
timestamp 1669390400
transform 1 0 9296 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_529
timestamp 1669390400
transform 1 0 17248 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_530
timestamp 1669390400
transform 1 0 25200 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_531
timestamp 1669390400
transform 1 0 33152 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_532
timestamp 1669390400
transform 1 0 41104 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_533
timestamp 1669390400
transform 1 0 49056 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_534
timestamp 1669390400
transform 1 0 57008 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_535
timestamp 1669390400
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_536
timestamp 1669390400
transform 1 0 13216 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_537
timestamp 1669390400
transform 1 0 21168 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_538
timestamp 1669390400
transform 1 0 29120 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_539
timestamp 1669390400
transform 1 0 37072 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_540
timestamp 1669390400
transform 1 0 45024 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_541
timestamp 1669390400
transform 1 0 52976 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_542
timestamp 1669390400
transform 1 0 9296 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_543
timestamp 1669390400
transform 1 0 17248 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_544
timestamp 1669390400
transform 1 0 25200 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_545
timestamp 1669390400
transform 1 0 33152 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_546
timestamp 1669390400
transform 1 0 41104 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_547
timestamp 1669390400
transform 1 0 49056 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_548
timestamp 1669390400
transform 1 0 57008 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_549
timestamp 1669390400
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_550
timestamp 1669390400
transform 1 0 13216 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_551
timestamp 1669390400
transform 1 0 21168 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_552
timestamp 1669390400
transform 1 0 29120 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_553
timestamp 1669390400
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_554
timestamp 1669390400
transform 1 0 45024 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_555
timestamp 1669390400
transform 1 0 52976 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_556
timestamp 1669390400
transform 1 0 9296 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_557
timestamp 1669390400
transform 1 0 17248 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_558
timestamp 1669390400
transform 1 0 25200 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_559
timestamp 1669390400
transform 1 0 33152 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_560
timestamp 1669390400
transform 1 0 41104 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_561
timestamp 1669390400
transform 1 0 49056 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_562
timestamp 1669390400
transform 1 0 57008 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_563
timestamp 1669390400
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_564
timestamp 1669390400
transform 1 0 13216 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_565
timestamp 1669390400
transform 1 0 21168 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_566
timestamp 1669390400
transform 1 0 29120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_567
timestamp 1669390400
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_568
timestamp 1669390400
transform 1 0 45024 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_569
timestamp 1669390400
transform 1 0 52976 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_570
timestamp 1669390400
transform 1 0 9296 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_571
timestamp 1669390400
transform 1 0 17248 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_572
timestamp 1669390400
transform 1 0 25200 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_573
timestamp 1669390400
transform 1 0 33152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_574
timestamp 1669390400
transform 1 0 41104 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_575
timestamp 1669390400
transform 1 0 49056 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_576
timestamp 1669390400
transform 1 0 57008 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_577
timestamp 1669390400
transform 1 0 5264 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_578
timestamp 1669390400
transform 1 0 13216 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_579
timestamp 1669390400
transform 1 0 21168 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_580
timestamp 1669390400
transform 1 0 29120 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_581
timestamp 1669390400
transform 1 0 37072 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_582
timestamp 1669390400
transform 1 0 45024 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_583
timestamp 1669390400
transform 1 0 52976 0 1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_584
timestamp 1669390400
transform 1 0 9296 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_585
timestamp 1669390400
transform 1 0 17248 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_586
timestamp 1669390400
transform 1 0 25200 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_587
timestamp 1669390400
transform 1 0 33152 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_588
timestamp 1669390400
transform 1 0 41104 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_589
timestamp 1669390400
transform 1 0 49056 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_590
timestamp 1669390400
transform 1 0 57008 0 -1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_591
timestamp 1669390400
transform 1 0 5264 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_592
timestamp 1669390400
transform 1 0 13216 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_593
timestamp 1669390400
transform 1 0 21168 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_594
timestamp 1669390400
transform 1 0 29120 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_595
timestamp 1669390400
transform 1 0 37072 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_596
timestamp 1669390400
transform 1 0 45024 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_597
timestamp 1669390400
transform 1 0 52976 0 1 53312
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_598
timestamp 1669390400
transform 1 0 9296 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_599
timestamp 1669390400
transform 1 0 17248 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_600
timestamp 1669390400
transform 1 0 25200 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_601
timestamp 1669390400
transform 1 0 33152 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_602
timestamp 1669390400
transform 1 0 41104 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_603
timestamp 1669390400
transform 1 0 49056 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_604
timestamp 1669390400
transform 1 0 57008 0 -1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_605
timestamp 1669390400
transform 1 0 5264 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_606
timestamp 1669390400
transform 1 0 13216 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_607
timestamp 1669390400
transform 1 0 21168 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_608
timestamp 1669390400
transform 1 0 29120 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_609
timestamp 1669390400
transform 1 0 37072 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_610
timestamp 1669390400
transform 1 0 45024 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_611
timestamp 1669390400
transform 1 0 52976 0 1 54880
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_612
timestamp 1669390400
transform 1 0 5264 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_613
timestamp 1669390400
transform 1 0 9184 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_614
timestamp 1669390400
transform 1 0 13104 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_615
timestamp 1669390400
transform 1 0 17024 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_616
timestamp 1669390400
transform 1 0 20944 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_617
timestamp 1669390400
transform 1 0 24864 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_618
timestamp 1669390400
transform 1 0 28784 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_619
timestamp 1669390400
transform 1 0 32704 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_620
timestamp 1669390400
transform 1 0 36624 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_621
timestamp 1669390400
transform 1 0 40544 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_622
timestamp 1669390400
transform 1 0 44464 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_623
timestamp 1669390400
transform 1 0 48384 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_624
timestamp 1669390400
transform 1 0 52304 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_625
timestamp 1669390400
transform 1 0 56224 0 -1 56448
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1444_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 51184 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1445_
timestamp 1669390400
transform -1 0 54656 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1446_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 54432 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1447_
timestamp 1669390400
transform 1 0 54208 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1448_
timestamp 1669390400
transform -1 0 56896 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1449_
timestamp 1669390400
transform -1 0 57680 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1450_
timestamp 1669390400
transform 1 0 45248 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1451_
timestamp 1669390400
transform -1 0 47152 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1452_
timestamp 1669390400
transform -1 0 58016 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1453_
timestamp 1669390400
transform -1 0 58016 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1454_
timestamp 1669390400
transform -1 0 58016 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1455_
timestamp 1669390400
transform -1 0 56448 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1456_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 54096 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1457_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 55328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1458_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 39760 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1459_
timestamp 1669390400
transform 1 0 38976 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1669390400
transform 1 0 21616 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1461_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 17136 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1462_
timestamp 1669390400
transform -1 0 12544 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1463_
timestamp 1669390400
transform -1 0 23520 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1464_
timestamp 1669390400
transform 1 0 25984 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1465_
timestamp 1669390400
transform -1 0 25424 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1466_
timestamp 1669390400
transform -1 0 22288 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1467_
timestamp 1669390400
transform 1 0 21392 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1468_
timestamp 1669390400
transform 1 0 22960 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1469_
timestamp 1669390400
transform 1 0 26880 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1470_
timestamp 1669390400
transform -1 0 24864 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1471_
timestamp 1669390400
transform -1 0 19936 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1472_
timestamp 1669390400
transform 1 0 19936 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1473_
timestamp 1669390400
transform 1 0 21840 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1474_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 23184 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1475_
timestamp 1669390400
transform -1 0 4032 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1476_
timestamp 1669390400
transform -1 0 28896 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1477_
timestamp 1669390400
transform -1 0 28784 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1478_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22960 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1479_
timestamp 1669390400
transform 1 0 23520 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1480_
timestamp 1669390400
transform -1 0 7952 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1669390400
transform -1 0 5152 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1482_
timestamp 1669390400
transform -1 0 18368 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1483_
timestamp 1669390400
transform 1 0 19488 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1484_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 5600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1485_
timestamp 1669390400
transform -1 0 19488 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1486_
timestamp 1669390400
transform -1 0 6384 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1487_
timestamp 1669390400
transform -1 0 30128 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1488_
timestamp 1669390400
transform 1 0 25648 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1489_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 23408 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1490_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22736 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1491_
timestamp 1669390400
transform -1 0 21056 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1492_
timestamp 1669390400
transform 1 0 10528 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1493_
timestamp 1669390400
transform 1 0 23632 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1494_
timestamp 1669390400
transform 1 0 23632 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1495_
timestamp 1669390400
transform -1 0 23968 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1496_
timestamp 1669390400
transform -1 0 10528 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1497_
timestamp 1669390400
transform 1 0 10192 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1498_
timestamp 1669390400
transform -1 0 30128 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1499_
timestamp 1669390400
transform -1 0 29680 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1500_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10416 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1501_
timestamp 1669390400
transform 1 0 22288 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1502_
timestamp 1669390400
transform -1 0 21056 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1503_
timestamp 1669390400
transform -1 0 21168 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1504_
timestamp 1669390400
transform 1 0 19040 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1505_
timestamp 1669390400
transform -1 0 23408 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1506_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22848 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1507_
timestamp 1669390400
transform 1 0 23408 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1508_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23184 0 -1 29792
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1509_
timestamp 1669390400
transform -1 0 24976 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1510_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22400 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1511_
timestamp 1669390400
transform -1 0 24080 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1512_
timestamp 1669390400
transform -1 0 50064 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1513_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 47824 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1514_
timestamp 1669390400
transform 1 0 43344 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1515_
timestamp 1669390400
transform 1 0 39424 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1516_
timestamp 1669390400
transform 1 0 33488 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1517_
timestamp 1669390400
transform -1 0 31696 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1518_
timestamp 1669390400
transform 1 0 31136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1519_
timestamp 1669390400
transform 1 0 31360 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1520_
timestamp 1669390400
transform 1 0 28336 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1521_
timestamp 1669390400
transform -1 0 32704 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1522_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 30576 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1523_
timestamp 1669390400
transform -1 0 30352 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1524_
timestamp 1669390400
transform -1 0 30912 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1525_
timestamp 1669390400
transform -1 0 17472 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1526_
timestamp 1669390400
transform 1 0 17584 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1527_
timestamp 1669390400
transform -1 0 20832 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1528_
timestamp 1669390400
transform -1 0 18256 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1529_
timestamp 1669390400
transform -1 0 14224 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1530_
timestamp 1669390400
transform -1 0 27888 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1531_
timestamp 1669390400
transform 1 0 26544 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1532_
timestamp 1669390400
transform -1 0 26320 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1533_
timestamp 1669390400
transform -1 0 26768 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1534_
timestamp 1669390400
transform 1 0 29568 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1535_
timestamp 1669390400
transform 1 0 30688 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1536_
timestamp 1669390400
transform 1 0 27216 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1669390400
transform -1 0 28112 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1538_
timestamp 1669390400
transform 1 0 27104 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1539_
timestamp 1669390400
transform -1 0 17024 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1540_
timestamp 1669390400
transform 1 0 22064 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1541_
timestamp 1669390400
transform 1 0 8400 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1542_
timestamp 1669390400
transform -1 0 7504 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1543_
timestamp 1669390400
transform -1 0 13328 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1544_
timestamp 1669390400
transform 1 0 11760 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1545_
timestamp 1669390400
transform -1 0 5712 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1546_
timestamp 1669390400
transform -1 0 15344 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1547_
timestamp 1669390400
transform 1 0 15008 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1548_
timestamp 1669390400
transform -1 0 4480 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1549_
timestamp 1669390400
transform -1 0 5264 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1550_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 13216 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1551_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 12320 0 -1 7840
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1552_
timestamp 1669390400
transform -1 0 26992 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1553_
timestamp 1669390400
transform -1 0 27664 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1554_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 19712 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1555_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 16240 0 1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1556_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7056 0 -1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1557_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 18704 0 1 7840
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1558_
timestamp 1669390400
transform -1 0 17136 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1559_
timestamp 1669390400
transform -1 0 29008 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1560_
timestamp 1669390400
transform -1 0 9184 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1561_
timestamp 1669390400
transform 1 0 16464 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1562_
timestamp 1669390400
transform 1 0 15456 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1563_
timestamp 1669390400
transform 1 0 2016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1564_
timestamp 1669390400
transform -1 0 2800 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1565_
timestamp 1669390400
transform -1 0 4144 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1566_
timestamp 1669390400
transform -1 0 3920 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1567_
timestamp 1669390400
transform -1 0 3584 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1568_
timestamp 1669390400
transform 1 0 24416 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1569_
timestamp 1669390400
transform -1 0 25200 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1570_
timestamp 1669390400
transform -1 0 14560 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1571_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7504 0 1 6272
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1572_
timestamp 1669390400
transform -1 0 5712 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1573_
timestamp 1669390400
transform -1 0 4928 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1574_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11424 0 1 14112
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1575_
timestamp 1669390400
transform 1 0 9632 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1576_
timestamp 1669390400
transform -1 0 14672 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1577_
timestamp 1669390400
transform -1 0 28672 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1578_
timestamp 1669390400
transform -1 0 28112 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1579_
timestamp 1669390400
transform -1 0 28448 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1580_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7840 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1581_
timestamp 1669390400
transform 1 0 8064 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1582_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 13104 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1583_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 12656 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1584_
timestamp 1669390400
transform -1 0 12432 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1585_
timestamp 1669390400
transform 1 0 8288 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1586_
timestamp 1669390400
transform 1 0 9520 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1587_
timestamp 1669390400
transform 1 0 4256 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1588_
timestamp 1669390400
transform -1 0 5152 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1589_
timestamp 1669390400
transform 1 0 27552 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1590_
timestamp 1669390400
transform -1 0 9856 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1591_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25312 0 1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1592_
timestamp 1669390400
transform -1 0 26768 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1593_
timestamp 1669390400
transform 1 0 8288 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1594_
timestamp 1669390400
transform 1 0 12096 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1595_
timestamp 1669390400
transform 1 0 12432 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1596_
timestamp 1669390400
transform -1 0 27776 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1597_
timestamp 1669390400
transform 1 0 19600 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1598_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10976 0 -1 21952
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1599_
timestamp 1669390400
transform 1 0 2688 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1600_
timestamp 1669390400
transform -1 0 7168 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1601_
timestamp 1669390400
transform 1 0 15792 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1602_
timestamp 1669390400
transform -1 0 10304 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1603_
timestamp 1669390400
transform 1 0 10528 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1604_
timestamp 1669390400
transform 1 0 15680 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1605_
timestamp 1669390400
transform -1 0 15568 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1606_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 14560 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1607_
timestamp 1669390400
transform 1 0 4256 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1608_
timestamp 1669390400
transform -1 0 9184 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1609_
timestamp 1669390400
transform -1 0 7616 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1610_
timestamp 1669390400
transform 1 0 5152 0 -1 17248
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1611_
timestamp 1669390400
transform 1 0 2800 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1612_
timestamp 1669390400
transform 1 0 2688 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1669390400
transform 1 0 3024 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1614_
timestamp 1669390400
transform 1 0 2912 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1615_
timestamp 1669390400
transform -1 0 14784 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1616_
timestamp 1669390400
transform 1 0 12208 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1617_
timestamp 1669390400
transform -1 0 10192 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1618_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 4144 0 -1 21952
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _1619_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 2576 0 -1 23520
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1620_
timestamp 1669390400
transform -1 0 26880 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1621_
timestamp 1669390400
transform 1 0 26320 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1622_
timestamp 1669390400
transform -1 0 25760 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1623_
timestamp 1669390400
transform 1 0 13552 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1624_
timestamp 1669390400
transform -1 0 9968 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1625_
timestamp 1669390400
transform -1 0 6832 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1626_
timestamp 1669390400
transform -1 0 7168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1627_
timestamp 1669390400
transform -1 0 27552 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1628_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 22288 0 -1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1629_
timestamp 1669390400
transform 1 0 25648 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1630_
timestamp 1669390400
transform -1 0 24528 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1631_
timestamp 1669390400
transform -1 0 23408 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1632_
timestamp 1669390400
transform -1 0 30016 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1633_
timestamp 1669390400
transform 1 0 26768 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1634_
timestamp 1669390400
transform -1 0 19264 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1635_
timestamp 1669390400
transform 1 0 23184 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1636_
timestamp 1669390400
transform -1 0 6048 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1637_
timestamp 1669390400
transform -1 0 5600 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1638_
timestamp 1669390400
transform -1 0 5152 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1639_
timestamp 1669390400
transform 1 0 11088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1640_
timestamp 1669390400
transform 1 0 5712 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1641_
timestamp 1669390400
transform -1 0 8064 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1642_
timestamp 1669390400
transform 1 0 6496 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1643_
timestamp 1669390400
transform 1 0 9184 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1644_
timestamp 1669390400
transform -1 0 28112 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1645_
timestamp 1669390400
transform -1 0 29232 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1669390400
transform -1 0 9520 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1647_
timestamp 1669390400
transform -1 0 13888 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1648_
timestamp 1669390400
transform -1 0 9184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1649_
timestamp 1669390400
transform 1 0 13216 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1650_
timestamp 1669390400
transform -1 0 10976 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1651_
timestamp 1669390400
transform 1 0 14448 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1652_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 15792 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1653_
timestamp 1669390400
transform -1 0 5824 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1654_
timestamp 1669390400
transform -1 0 5376 0 -1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1669390400
transform 1 0 2016 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1656_
timestamp 1669390400
transform 1 0 3472 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1657_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3808 0 -1 25088
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1658_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 10864 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1659_
timestamp 1669390400
transform 1 0 9968 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1660_
timestamp 1669390400
transform 1 0 11088 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1661_
timestamp 1669390400
transform 1 0 23184 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1662_
timestamp 1669390400
transform -1 0 11536 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1663_
timestamp 1669390400
transform -1 0 9184 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1664_
timestamp 1669390400
transform 1 0 19152 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1665_
timestamp 1669390400
transform -1 0 8736 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1666_
timestamp 1669390400
transform -1 0 7504 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1667_
timestamp 1669390400
transform -1 0 9184 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1668_
timestamp 1669390400
transform 1 0 10640 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1669_
timestamp 1669390400
transform 1 0 9968 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1670_
timestamp 1669390400
transform 1 0 6160 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1671_
timestamp 1669390400
transform -1 0 5936 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1672_
timestamp 1669390400
transform 1 0 6160 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1673_
timestamp 1669390400
transform -1 0 7840 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1674_
timestamp 1669390400
transform 1 0 10976 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1675_
timestamp 1669390400
transform -1 0 12432 0 -1 28224
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1676_
timestamp 1669390400
transform 1 0 13552 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1677_
timestamp 1669390400
transform 1 0 24080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1678_
timestamp 1669390400
transform 1 0 17696 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1679_
timestamp 1669390400
transform 1 0 24304 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1680_
timestamp 1669390400
transform -1 0 24528 0 -1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1681_
timestamp 1669390400
transform 1 0 28336 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1682_
timestamp 1669390400
transform 1 0 29456 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1683_
timestamp 1669390400
transform -1 0 30576 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1684_
timestamp 1669390400
transform 1 0 24080 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1685_
timestamp 1669390400
transform -1 0 18928 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1686_
timestamp 1669390400
transform 1 0 17136 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1687_
timestamp 1669390400
transform 1 0 3920 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1688_
timestamp 1669390400
transform -1 0 7728 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1689_
timestamp 1669390400
transform 1 0 6160 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1690_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 7056 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1691_
timestamp 1669390400
transform -1 0 7392 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1692_
timestamp 1669390400
transform -1 0 8176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1693_
timestamp 1669390400
transform 1 0 6048 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1694_
timestamp 1669390400
transform -1 0 5152 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1695_
timestamp 1669390400
transform 1 0 6608 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1696_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 12320 0 1 7840
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1697_
timestamp 1669390400
transform 1 0 7392 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1698_
timestamp 1669390400
transform -1 0 26768 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1699_
timestamp 1669390400
transform 1 0 24864 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1700_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 6496 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1701_
timestamp 1669390400
transform 1 0 5824 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1702_
timestamp 1669390400
transform 1 0 7056 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1703_
timestamp 1669390400
transform 1 0 17920 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1704_
timestamp 1669390400
transform -1 0 20720 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1705_
timestamp 1669390400
transform -1 0 30576 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1706_
timestamp 1669390400
transform 1 0 18368 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1707_
timestamp 1669390400
transform -1 0 17136 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _1708_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 8624 0 -1 20384
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1709_
timestamp 1669390400
transform 1 0 28784 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1710_
timestamp 1669390400
transform 1 0 5936 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _1711_
timestamp 1669390400
transform 1 0 7056 0 1 20384
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1712_
timestamp 1669390400
transform 1 0 19936 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1713_
timestamp 1669390400
transform 1 0 10752 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1714_
timestamp 1669390400
transform 1 0 11088 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1715_
timestamp 1669390400
transform -1 0 15008 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1716_
timestamp 1669390400
transform 1 0 23520 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_2  _1717_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 25424 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1718_
timestamp 1669390400
transform 1 0 29232 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1719_
timestamp 1669390400
transform 1 0 26880 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1720_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 24304 0 1 21952
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1721_
timestamp 1669390400
transform -1 0 11200 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1722_
timestamp 1669390400
transform 1 0 10864 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1723_
timestamp 1669390400
transform 1 0 8288 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1724_
timestamp 1669390400
transform -1 0 14336 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1725_
timestamp 1669390400
transform 1 0 9296 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1726_
timestamp 1669390400
transform -1 0 9072 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1727_
timestamp 1669390400
transform 1 0 7056 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1728_
timestamp 1669390400
transform -1 0 12656 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1729_
timestamp 1669390400
transform -1 0 22624 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1730_
timestamp 1669390400
transform -1 0 19152 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1731_
timestamp 1669390400
transform -1 0 12544 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1732_
timestamp 1669390400
transform 1 0 12432 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1733_
timestamp 1669390400
transform 1 0 12096 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1734_
timestamp 1669390400
transform -1 0 14112 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1735_
timestamp 1669390400
transform 1 0 14112 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _1736_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 11872 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1737_
timestamp 1669390400
transform 1 0 25088 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1738_
timestamp 1669390400
transform 1 0 26208 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1739_
timestamp 1669390400
transform 1 0 5600 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1740_
timestamp 1669390400
transform 1 0 12656 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1741_
timestamp 1669390400
transform -1 0 13104 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1742_
timestamp 1669390400
transform -1 0 12656 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1743_
timestamp 1669390400
transform 1 0 8064 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1744_
timestamp 1669390400
transform 1 0 10976 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1745_
timestamp 1669390400
transform 1 0 18928 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1746_
timestamp 1669390400
transform 1 0 9632 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1747_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 9968 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1748_
timestamp 1669390400
transform 1 0 8512 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1749_
timestamp 1669390400
transform 1 0 10192 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1750_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7728 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1751_
timestamp 1669390400
transform 1 0 7168 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1752_
timestamp 1669390400
transform 1 0 5936 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1753_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 6608 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1754_
timestamp 1669390400
transform 1 0 10192 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1755_
timestamp 1669390400
transform 1 0 23408 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _1756_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 27776 0 -1 14112
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1757_
timestamp 1669390400
transform -1 0 29120 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1758_
timestamp 1669390400
transform -1 0 14448 0 -1 14112
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1759_
timestamp 1669390400
transform -1 0 6832 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1760_
timestamp 1669390400
transform 1 0 7616 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1761_
timestamp 1669390400
transform -1 0 11984 0 1 10976
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1762_
timestamp 1669390400
transform -1 0 11424 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1763_
timestamp 1669390400
transform 1 0 5824 0 1 12544
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1764_
timestamp 1669390400
transform -1 0 5600 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1765_
timestamp 1669390400
transform -1 0 6384 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1766_
timestamp 1669390400
transform 1 0 4480 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1767_
timestamp 1669390400
transform -1 0 11088 0 1 18816
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1768_
timestamp 1669390400
transform 1 0 9632 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1769_
timestamp 1669390400
transform -1 0 6272 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1770_
timestamp 1669390400
transform 1 0 13552 0 1 14112
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1771_
timestamp 1669390400
transform -1 0 18144 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1772_
timestamp 1669390400
transform 1 0 18704 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1773_
timestamp 1669390400
transform 1 0 12992 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1774_
timestamp 1669390400
transform 1 0 15904 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1775_
timestamp 1669390400
transform -1 0 19376 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1776_
timestamp 1669390400
transform -1 0 18816 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1777_
timestamp 1669390400
transform 1 0 9520 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1778_
timestamp 1669390400
transform 1 0 24192 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1779_
timestamp 1669390400
transform 1 0 23408 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1780_
timestamp 1669390400
transform -1 0 10976 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1781_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 14112 0 -1 23520
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1782_
timestamp 1669390400
transform -1 0 24528 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1783_
timestamp 1669390400
transform -1 0 24080 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1784_
timestamp 1669390400
transform 1 0 21952 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1785_
timestamp 1669390400
transform -1 0 15008 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1786_
timestamp 1669390400
transform 1 0 17808 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1787_
timestamp 1669390400
transform 1 0 24976 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1788_
timestamp 1669390400
transform 1 0 19600 0 -1 20384
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1789_
timestamp 1669390400
transform -1 0 19376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1790_
timestamp 1669390400
transform 1 0 20496 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1791_
timestamp 1669390400
transform -1 0 30912 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1792_
timestamp 1669390400
transform -1 0 8960 0 -1 10976
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1793_
timestamp 1669390400
transform -1 0 21056 0 1 18816
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _1794_
timestamp 1669390400
transform 1 0 11424 0 -1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1795_
timestamp 1669390400
transform 1 0 11760 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1796_
timestamp 1669390400
transform -1 0 13104 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1797_
timestamp 1669390400
transform 1 0 19600 0 1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1798_
timestamp 1669390400
transform 1 0 19936 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1799_
timestamp 1669390400
transform -1 0 22512 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1800_
timestamp 1669390400
transform 1 0 21168 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1801_
timestamp 1669390400
transform 1 0 22960 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1802_
timestamp 1669390400
transform -1 0 23968 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1803_
timestamp 1669390400
transform 1 0 17584 0 -1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1804_
timestamp 1669390400
transform -1 0 24304 0 -1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1805_
timestamp 1669390400
transform -1 0 16800 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1806_
timestamp 1669390400
transform 1 0 22512 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1807_
timestamp 1669390400
transform 1 0 15904 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _1808_
timestamp 1669390400
transform -1 0 12656 0 1 28224
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1809_
timestamp 1669390400
transform -1 0 16016 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1810_
timestamp 1669390400
transform -1 0 5376 0 -1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1811_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 3920 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1812_
timestamp 1669390400
transform 1 0 13216 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1813_
timestamp 1669390400
transform 1 0 13664 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1814_
timestamp 1669390400
transform -1 0 15904 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1815_
timestamp 1669390400
transform -1 0 11200 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1816_
timestamp 1669390400
transform 1 0 14896 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1817_
timestamp 1669390400
transform 1 0 19600 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1818_
timestamp 1669390400
transform -1 0 20384 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1819_
timestamp 1669390400
transform -1 0 15680 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1820_
timestamp 1669390400
transform -1 0 15232 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1821_
timestamp 1669390400
transform 1 0 14560 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1822_
timestamp 1669390400
transform 1 0 15232 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1823_
timestamp 1669390400
transform 1 0 14784 0 1 17248
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1824_
timestamp 1669390400
transform -1 0 12992 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1825_
timestamp 1669390400
transform 1 0 5600 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1826_
timestamp 1669390400
transform 1 0 4480 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1827_
timestamp 1669390400
transform -1 0 6720 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1828_
timestamp 1669390400
transform 1 0 5264 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1829_
timestamp 1669390400
transform -1 0 4144 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1830_
timestamp 1669390400
transform 1 0 1904 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1831_
timestamp 1669390400
transform -1 0 2912 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1832_
timestamp 1669390400
transform -1 0 6608 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1833_
timestamp 1669390400
transform -1 0 5152 0 1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1834_
timestamp 1669390400
transform -1 0 6832 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1835_
timestamp 1669390400
transform 1 0 7056 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1836_
timestamp 1669390400
transform 1 0 5712 0 1 7840
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1837_
timestamp 1669390400
transform -1 0 10416 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1838_
timestamp 1669390400
transform 1 0 6832 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1839_
timestamp 1669390400
transform 1 0 14784 0 1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1840_
timestamp 1669390400
transform 1 0 13552 0 1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1841_
timestamp 1669390400
transform -1 0 18256 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1842_
timestamp 1669390400
transform 1 0 6048 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1843_
timestamp 1669390400
transform -1 0 21056 0 1 10976
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _1844_
timestamp 1669390400
transform -1 0 10976 0 1 10976
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1845_
timestamp 1669390400
transform -1 0 5824 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1846_
timestamp 1669390400
transform 1 0 3696 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1847_
timestamp 1669390400
transform 1 0 6944 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1848_
timestamp 1669390400
transform 1 0 8064 0 1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1849_
timestamp 1669390400
transform -1 0 22288 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1850_
timestamp 1669390400
transform 1 0 17584 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1851_
timestamp 1669390400
transform -1 0 22400 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1852_
timestamp 1669390400
transform -1 0 20272 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1853_
timestamp 1669390400
transform 1 0 18368 0 -1 12544
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1854_
timestamp 1669390400
transform -1 0 19376 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _1855_
timestamp 1669390400
transform 1 0 17696 0 -1 18816
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1856_
timestamp 1669390400
transform -1 0 17136 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1857_
timestamp 1669390400
transform 1 0 15344 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1858_
timestamp 1669390400
transform 1 0 15680 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1859_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 15120 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1860_
timestamp 1669390400
transform -1 0 11648 0 1 37632
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _1861_
timestamp 1669390400
transform 1 0 10416 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1862_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 10752 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1863_
timestamp 1669390400
transform 1 0 13552 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1864_
timestamp 1669390400
transform 1 0 14784 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1865_
timestamp 1669390400
transform -1 0 14224 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1866_
timestamp 1669390400
transform 1 0 13552 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _1867_
timestamp 1669390400
transform 1 0 10416 0 1 12544
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1868_
timestamp 1669390400
transform 1 0 19936 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1869_
timestamp 1669390400
transform -1 0 17136 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1870_
timestamp 1669390400
transform 1 0 15680 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1871_
timestamp 1669390400
transform 1 0 28336 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1872_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 20496 0 -1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1873_
timestamp 1669390400
transform -1 0 22848 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1874_
timestamp 1669390400
transform 1 0 14896 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1875_
timestamp 1669390400
transform -1 0 24080 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1876_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 23632 0 1 23520
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1877_
timestamp 1669390400
transform 1 0 21952 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1878_
timestamp 1669390400
transform -1 0 16464 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1879_
timestamp 1669390400
transform -1 0 11424 0 -1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1880_
timestamp 1669390400
transform 1 0 2800 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1881_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 4256 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1882_
timestamp 1669390400
transform 1 0 2240 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1883_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 12768 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1884_
timestamp 1669390400
transform -1 0 10752 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1885_
timestamp 1669390400
transform -1 0 14448 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1886_
timestamp 1669390400
transform 1 0 5600 0 1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1887_
timestamp 1669390400
transform -1 0 7280 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1888_
timestamp 1669390400
transform 1 0 14336 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1889_
timestamp 1669390400
transform -1 0 15792 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1890_
timestamp 1669390400
transform -1 0 14448 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1891_
timestamp 1669390400
transform -1 0 11984 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1892_
timestamp 1669390400
transform -1 0 11312 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1893_
timestamp 1669390400
transform 1 0 7952 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1894_
timestamp 1669390400
transform 1 0 8288 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1895_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 7616 0 1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1896_
timestamp 1669390400
transform 1 0 7392 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1897_
timestamp 1669390400
transform -1 0 8848 0 1 34496
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1898_
timestamp 1669390400
transform 1 0 12768 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1899_
timestamp 1669390400
transform 1 0 13664 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1900_
timestamp 1669390400
transform 1 0 29680 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1901_
timestamp 1669390400
transform 1 0 9968 0 -1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1902_
timestamp 1669390400
transform -1 0 22176 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1903_
timestamp 1669390400
transform -1 0 15008 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1904_
timestamp 1669390400
transform 1 0 16016 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1905_
timestamp 1669390400
transform 1 0 16240 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1906_
timestamp 1669390400
transform 1 0 16576 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1907_
timestamp 1669390400
transform 1 0 17584 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1908_
timestamp 1669390400
transform -1 0 14560 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1909_
timestamp 1669390400
transform -1 0 16352 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1910_
timestamp 1669390400
transform 1 0 13664 0 -1 36064
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1911_
timestamp 1669390400
transform -1 0 17136 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1912_
timestamp 1669390400
transform 1 0 14560 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1913_
timestamp 1669390400
transform -1 0 12656 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1914_
timestamp 1669390400
transform 1 0 7728 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1915_
timestamp 1669390400
transform -1 0 18368 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1916_
timestamp 1669390400
transform -1 0 12992 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1917_
timestamp 1669390400
transform -1 0 15008 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1918_
timestamp 1669390400
transform 1 0 13216 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _1919_
timestamp 1669390400
transform -1 0 15456 0 1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1920_
timestamp 1669390400
transform -1 0 14672 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _1921_
timestamp 1669390400
transform 1 0 11984 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1922_
timestamp 1669390400
transform 1 0 13552 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1923_
timestamp 1669390400
transform 1 0 16240 0 1 23520
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1924_
timestamp 1669390400
transform -1 0 17360 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1925_
timestamp 1669390400
transform 1 0 25536 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1926_
timestamp 1669390400
transform -1 0 21392 0 -1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1927_
timestamp 1669390400
transform -1 0 21056 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1928_
timestamp 1669390400
transform -1 0 22400 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1929_
timestamp 1669390400
transform -1 0 22288 0 1 25088
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1930_
timestamp 1669390400
transform -1 0 18256 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1931_
timestamp 1669390400
transform 1 0 16016 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1932_
timestamp 1669390400
transform -1 0 17024 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1933_
timestamp 1669390400
transform -1 0 13552 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1934_
timestamp 1669390400
transform -1 0 11088 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1935_
timestamp 1669390400
transform 1 0 4704 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1936_
timestamp 1669390400
transform 1 0 6832 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1937_
timestamp 1669390400
transform -1 0 8624 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1938_
timestamp 1669390400
transform 1 0 6384 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _1939_
timestamp 1669390400
transform 1 0 6160 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1940_
timestamp 1669390400
transform 1 0 8624 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1941_
timestamp 1669390400
transform 1 0 9632 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1942_
timestamp 1669390400
transform 1 0 26768 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1943_
timestamp 1669390400
transform 1 0 13552 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1944_
timestamp 1669390400
transform 1 0 13552 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1945_
timestamp 1669390400
transform 1 0 13776 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1946_
timestamp 1669390400
transform 1 0 6832 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1947_
timestamp 1669390400
transform -1 0 7504 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1948_
timestamp 1669390400
transform -1 0 27888 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1949_
timestamp 1669390400
transform -1 0 26768 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1950_
timestamp 1669390400
transform -1 0 27888 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1951_
timestamp 1669390400
transform -1 0 9184 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1952_
timestamp 1669390400
transform -1 0 6496 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1953_
timestamp 1669390400
transform 1 0 6944 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1954_
timestamp 1669390400
transform 1 0 7952 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1955_
timestamp 1669390400
transform 1 0 6832 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1956_
timestamp 1669390400
transform -1 0 10640 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1957_
timestamp 1669390400
transform 1 0 7840 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1958_
timestamp 1669390400
transform 1 0 9632 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1959_
timestamp 1669390400
transform -1 0 16576 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1960_
timestamp 1669390400
transform -1 0 17248 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1961_
timestamp 1669390400
transform 1 0 15120 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1962_
timestamp 1669390400
transform 1 0 16240 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1963_
timestamp 1669390400
transform -1 0 25088 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1964_
timestamp 1669390400
transform 1 0 15680 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1965_
timestamp 1669390400
transform 1 0 18928 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1966_
timestamp 1669390400
transform 1 0 19600 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _1967_
timestamp 1669390400
transform -1 0 21952 0 -1 15680
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _1968_
timestamp 1669390400
transform 1 0 16688 0 1 15680
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1969_
timestamp 1669390400
transform 1 0 17248 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1970_
timestamp 1669390400
transform -1 0 19040 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _1971_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 16912 0 1 34496
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1972_
timestamp 1669390400
transform 1 0 17584 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1973_
timestamp 1669390400
transform -1 0 17136 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1974_
timestamp 1669390400
transform 1 0 17584 0 -1 39200
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1975_
timestamp 1669390400
transform -1 0 13104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1976_
timestamp 1669390400
transform -1 0 13328 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1977_
timestamp 1669390400
transform 1 0 11536 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1978_
timestamp 1669390400
transform 1 0 27664 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1979_
timestamp 1669390400
transform 1 0 13328 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1980_
timestamp 1669390400
transform -1 0 18144 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _1981_
timestamp 1669390400
transform 1 0 18368 0 -1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1982_
timestamp 1669390400
transform -1 0 24192 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1983_
timestamp 1669390400
transform -1 0 14224 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1984_
timestamp 1669390400
transform -1 0 8176 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1985_
timestamp 1669390400
transform -1 0 11872 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1986_
timestamp 1669390400
transform -1 0 10192 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1987_
timestamp 1669390400
transform 1 0 18480 0 1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1988_
timestamp 1669390400
transform 1 0 20384 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1989_
timestamp 1669390400
transform -1 0 19712 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1990_
timestamp 1669390400
transform 1 0 19936 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1991_
timestamp 1669390400
transform -1 0 19936 0 -1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _1992_
timestamp 1669390400
transform -1 0 14896 0 -1 48608
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1993_
timestamp 1669390400
transform -1 0 11984 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1994_
timestamp 1669390400
transform 1 0 9632 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1995_
timestamp 1669390400
transform -1 0 11088 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1996_
timestamp 1669390400
transform -1 0 9408 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1997_
timestamp 1669390400
transform -1 0 14448 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1998_
timestamp 1669390400
transform 1 0 13552 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1999_
timestamp 1669390400
transform 1 0 13664 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2000_
timestamp 1669390400
transform 1 0 23184 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2001_
timestamp 1669390400
transform 1 0 20720 0 -1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _2002_
timestamp 1669390400
transform -1 0 28896 0 1 20384
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2003_
timestamp 1669390400
transform -1 0 28112 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2004_
timestamp 1669390400
transform -1 0 27216 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2005_
timestamp 1669390400
transform 1 0 27440 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2006_
timestamp 1669390400
transform 1 0 26768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2007_
timestamp 1669390400
transform -1 0 9520 0 1 31360
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2008_
timestamp 1669390400
transform -1 0 19152 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2009_
timestamp 1669390400
transform 1 0 17136 0 1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2010_
timestamp 1669390400
transform -1 0 15008 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2011_
timestamp 1669390400
transform 1 0 13888 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2012_
timestamp 1669390400
transform -1 0 13104 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2013_
timestamp 1669390400
transform 1 0 10080 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2014_
timestamp 1669390400
transform 1 0 11424 0 1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2015_
timestamp 1669390400
transform 1 0 11872 0 -1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2016_
timestamp 1669390400
transform 1 0 15008 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2017_
timestamp 1669390400
transform 1 0 15456 0 -1 42336
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2018_
timestamp 1669390400
transform 1 0 15120 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2019_
timestamp 1669390400
transform 1 0 14672 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2020_
timestamp 1669390400
transform 1 0 14896 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2021_
timestamp 1669390400
transform 1 0 19264 0 -1 31360
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2022_
timestamp 1669390400
transform 1 0 22960 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2023_
timestamp 1669390400
transform -1 0 17920 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2024_
timestamp 1669390400
transform -1 0 15568 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2025_
timestamp 1669390400
transform -1 0 16912 0 1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2026_
timestamp 1669390400
transform 1 0 15568 0 -1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2027_
timestamp 1669390400
transform 1 0 15904 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2028_
timestamp 1669390400
transform -1 0 10640 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2029_
timestamp 1669390400
transform 1 0 12208 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2030_
timestamp 1669390400
transform 1 0 13552 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2031_
timestamp 1669390400
transform 1 0 13104 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2032_
timestamp 1669390400
transform -1 0 13104 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2033_
timestamp 1669390400
transform 1 0 15680 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2034_
timestamp 1669390400
transform -1 0 17136 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2035_
timestamp 1669390400
transform -1 0 2912 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2036_
timestamp 1669390400
transform 1 0 16240 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2037_
timestamp 1669390400
transform 1 0 16128 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2038_
timestamp 1669390400
transform 1 0 17696 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2039_
timestamp 1669390400
transform 1 0 17584 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2040_
timestamp 1669390400
transform 1 0 13552 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2041_
timestamp 1669390400
transform -1 0 17136 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2042_
timestamp 1669390400
transform -1 0 23744 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2043_
timestamp 1669390400
transform 1 0 18480 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2044_
timestamp 1669390400
transform 1 0 18032 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2045_
timestamp 1669390400
transform 1 0 19376 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2046_
timestamp 1669390400
transform 1 0 21504 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2047_
timestamp 1669390400
transform -1 0 30352 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2048_
timestamp 1669390400
transform 1 0 21616 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2049_
timestamp 1669390400
transform 1 0 20048 0 -1 25088
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2050_
timestamp 1669390400
transform 1 0 19376 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2051_
timestamp 1669390400
transform 1 0 14224 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2052_
timestamp 1669390400
transform 1 0 21504 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2053_
timestamp 1669390400
transform -1 0 22176 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2054_
timestamp 1669390400
transform 1 0 19712 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2055_
timestamp 1669390400
transform 1 0 21504 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2056_
timestamp 1669390400
transform -1 0 21056 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2057_
timestamp 1669390400
transform 1 0 19712 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2058_
timestamp 1669390400
transform -1 0 20608 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2059_
timestamp 1669390400
transform 1 0 24192 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2060_
timestamp 1669390400
transform 1 0 26208 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2061_
timestamp 1669390400
transform 1 0 25872 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2062_
timestamp 1669390400
transform 1 0 25088 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2063_
timestamp 1669390400
transform -1 0 25088 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2064_
timestamp 1669390400
transform -1 0 21056 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2065_
timestamp 1669390400
transform 1 0 18816 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2066_
timestamp 1669390400
transform 1 0 16576 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2067_
timestamp 1669390400
transform 1 0 17584 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2068_
timestamp 1669390400
transform 1 0 19040 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2069_
timestamp 1669390400
transform 1 0 50064 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2070_
timestamp 1669390400
transform -1 0 20608 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2071_
timestamp 1669390400
transform 1 0 19936 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2072_
timestamp 1669390400
transform 1 0 19600 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2073_
timestamp 1669390400
transform 1 0 25536 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2074_
timestamp 1669390400
transform -1 0 20272 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2075_
timestamp 1669390400
transform 1 0 18928 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2076_
timestamp 1669390400
transform 1 0 18144 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2077_
timestamp 1669390400
transform 1 0 19264 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2078_
timestamp 1669390400
transform -1 0 21056 0 1 26656
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2079_
timestamp 1669390400
transform 1 0 19376 0 1 39200
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2080_
timestamp 1669390400
transform -1 0 19936 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2081_
timestamp 1669390400
transform 1 0 19712 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2082_
timestamp 1669390400
transform 1 0 23968 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2083_
timestamp 1669390400
transform -1 0 26544 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2084_
timestamp 1669390400
transform -1 0 25760 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2085_
timestamp 1669390400
transform 1 0 27776 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2086_
timestamp 1669390400
transform -1 0 28784 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2087_
timestamp 1669390400
transform -1 0 28224 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2088_
timestamp 1669390400
transform 1 0 25424 0 1 26656
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2089_
timestamp 1669390400
transform 1 0 24416 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2090_
timestamp 1669390400
transform -1 0 25312 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2091_
timestamp 1669390400
transform -1 0 25088 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2092_
timestamp 1669390400
transform -1 0 23744 0 1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2093_
timestamp 1669390400
transform -1 0 22176 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2094_
timestamp 1669390400
transform 1 0 19600 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2095_
timestamp 1669390400
transform -1 0 24640 0 -1 26656
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2096_
timestamp 1669390400
transform 1 0 21616 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2097_
timestamp 1669390400
transform 1 0 22176 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2098_
timestamp 1669390400
transform 1 0 21504 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2099_
timestamp 1669390400
transform 1 0 22064 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2100_
timestamp 1669390400
transform 1 0 22176 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2101_
timestamp 1669390400
transform 1 0 16800 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2102_
timestamp 1669390400
transform -1 0 19152 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2103_
timestamp 1669390400
transform -1 0 19712 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2104_
timestamp 1669390400
transform -1 0 18816 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2105_
timestamp 1669390400
transform -1 0 18592 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2106_
timestamp 1669390400
transform -1 0 20160 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2107_
timestamp 1669390400
transform 1 0 25312 0 1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2108_
timestamp 1669390400
transform 1 0 26656 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2109_
timestamp 1669390400
transform 1 0 23968 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2110_
timestamp 1669390400
transform -1 0 23408 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2111_
timestamp 1669390400
transform 1 0 25536 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2112_
timestamp 1669390400
transform 1 0 19264 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2113_
timestamp 1669390400
transform -1 0 26656 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2114_
timestamp 1669390400
transform -1 0 26432 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2115_
timestamp 1669390400
transform 1 0 20720 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2116_
timestamp 1669390400
transform 1 0 21392 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2117_
timestamp 1669390400
transform -1 0 22400 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2118_
timestamp 1669390400
transform -1 0 21056 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2119_
timestamp 1669390400
transform 1 0 20496 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2120_
timestamp 1669390400
transform -1 0 29680 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2121_
timestamp 1669390400
transform 1 0 27888 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2122_
timestamp 1669390400
transform -1 0 28000 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2123_
timestamp 1669390400
transform -1 0 26096 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2124_
timestamp 1669390400
transform -1 0 27552 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2125_
timestamp 1669390400
transform 1 0 24528 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2126_
timestamp 1669390400
transform -1 0 26432 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2127_
timestamp 1669390400
transform -1 0 25088 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2128_
timestamp 1669390400
transform -1 0 26432 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2129_
timestamp 1669390400
transform -1 0 26768 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2130_
timestamp 1669390400
transform 1 0 25200 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2131_
timestamp 1669390400
transform 1 0 22736 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2132_
timestamp 1669390400
transform -1 0 25088 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2133_
timestamp 1669390400
transform 1 0 25872 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2134_
timestamp 1669390400
transform -1 0 58016 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2135_
timestamp 1669390400
transform 1 0 9856 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2136_
timestamp 1669390400
transform 1 0 9744 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2137_
timestamp 1669390400
transform 1 0 17696 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2138_
timestamp 1669390400
transform -1 0 18704 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2139_
timestamp 1669390400
transform -1 0 27664 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2140_
timestamp 1669390400
transform -1 0 24640 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2141_
timestamp 1669390400
transform -1 0 27328 0 1 37632
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2142_
timestamp 1669390400
transform 1 0 20272 0 -1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2143_
timestamp 1669390400
transform -1 0 24864 0 1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2144_
timestamp 1669390400
transform 1 0 21504 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2145_
timestamp 1669390400
transform -1 0 27552 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2146_
timestamp 1669390400
transform -1 0 26208 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2147_
timestamp 1669390400
transform -1 0 26432 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2148_
timestamp 1669390400
transform 1 0 25872 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2149_
timestamp 1669390400
transform -1 0 26880 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2150_
timestamp 1669390400
transform 1 0 25536 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2151_
timestamp 1669390400
transform 1 0 24752 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2152_
timestamp 1669390400
transform -1 0 24976 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2153_
timestamp 1669390400
transform 1 0 25536 0 -1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2154_
timestamp 1669390400
transform 1 0 26880 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2155_
timestamp 1669390400
transform 1 0 29456 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2156_
timestamp 1669390400
transform -1 0 22176 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2157_
timestamp 1669390400
transform -1 0 22736 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2158_
timestamp 1669390400
transform 1 0 23296 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2159_
timestamp 1669390400
transform 1 0 21504 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2160_
timestamp 1669390400
transform -1 0 27552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2161_
timestamp 1669390400
transform -1 0 28448 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2162_
timestamp 1669390400
transform 1 0 20720 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2163_
timestamp 1669390400
transform 1 0 21616 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2164_
timestamp 1669390400
transform 1 0 22624 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2165_
timestamp 1669390400
transform -1 0 23072 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2166_
timestamp 1669390400
transform 1 0 22400 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2167_
timestamp 1669390400
transform -1 0 24640 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2168_
timestamp 1669390400
transform 1 0 22400 0 -1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2169_
timestamp 1669390400
transform 1 0 23744 0 1 50176
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2170_
timestamp 1669390400
transform -1 0 26656 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2171_
timestamp 1669390400
transform 1 0 27664 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2172_
timestamp 1669390400
transform -1 0 27328 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2173_
timestamp 1669390400
transform -1 0 2912 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2174_
timestamp 1669390400
transform 1 0 26320 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2175_
timestamp 1669390400
transform 1 0 23296 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2176_
timestamp 1669390400
transform -1 0 24416 0 -1 50176
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2177_
timestamp 1669390400
transform 1 0 24416 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2178_
timestamp 1669390400
transform -1 0 22176 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2179_
timestamp 1669390400
transform 1 0 23296 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2180_
timestamp 1669390400
transform 1 0 18928 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2181_
timestamp 1669390400
transform -1 0 27664 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2182_
timestamp 1669390400
transform 1 0 10192 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2183_
timestamp 1669390400
transform -1 0 10304 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2184_
timestamp 1669390400
transform -1 0 52080 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2185_
timestamp 1669390400
transform -1 0 46928 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2186_
timestamp 1669390400
transform -1 0 47152 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2187_
timestamp 1669390400
transform 1 0 45248 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2188_
timestamp 1669390400
transform 1 0 52304 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2189_
timestamp 1669390400
transform -1 0 57120 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2190_
timestamp 1669390400
transform -1 0 55104 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2191_
timestamp 1669390400
transform 1 0 45360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2192_
timestamp 1669390400
transform -1 0 45584 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2193_
timestamp 1669390400
transform 1 0 48496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2194_
timestamp 1669390400
transform 1 0 49392 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2195_
timestamp 1669390400
transform -1 0 47152 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2196_
timestamp 1669390400
transform -1 0 49056 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2197_
timestamp 1669390400
transform 1 0 47376 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2198_
timestamp 1669390400
transform 1 0 52192 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2199_
timestamp 1669390400
transform 1 0 52864 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2200_
timestamp 1669390400
transform -1 0 48608 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2201_
timestamp 1669390400
transform -1 0 46032 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2202_
timestamp 1669390400
transform -1 0 48496 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2203_
timestamp 1669390400
transform 1 0 43344 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2204_
timestamp 1669390400
transform -1 0 53088 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2205_
timestamp 1669390400
transform -1 0 58240 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2206_
timestamp 1669390400
transform -1 0 47152 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2207_
timestamp 1669390400
transform 1 0 41104 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2208_
timestamp 1669390400
transform 1 0 42112 0 1 21952
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2209_
timestamp 1669390400
transform 1 0 55216 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2210_
timestamp 1669390400
transform -1 0 52976 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2211_
timestamp 1669390400
transform 1 0 43008 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _2212_
timestamp 1669390400
transform 1 0 57344 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2213_
timestamp 1669390400
transform -1 0 58016 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2214_
timestamp 1669390400
transform 1 0 41440 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2215_
timestamp 1669390400
transform 1 0 56448 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2216_
timestamp 1669390400
transform -1 0 58016 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2217_
timestamp 1669390400
transform -1 0 51520 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2218_
timestamp 1669390400
transform -1 0 52080 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2219_
timestamp 1669390400
transform -1 0 44464 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2220_
timestamp 1669390400
transform -1 0 57568 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2221_
timestamp 1669390400
transform -1 0 58016 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2222_
timestamp 1669390400
transform 1 0 53312 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2223_
timestamp 1669390400
transform 1 0 44352 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2224_
timestamp 1669390400
transform -1 0 46704 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2225_
timestamp 1669390400
transform 1 0 45360 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2226_
timestamp 1669390400
transform -1 0 57456 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2227_
timestamp 1669390400
transform -1 0 56000 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2228_
timestamp 1669390400
transform 1 0 53984 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2229_
timestamp 1669390400
transform 1 0 56560 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2230_
timestamp 1669390400
transform -1 0 53648 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2231_
timestamp 1669390400
transform 1 0 52080 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2232_
timestamp 1669390400
transform -1 0 51968 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2233_
timestamp 1669390400
transform -1 0 49728 0 1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2234_
timestamp 1669390400
transform -1 0 46256 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2235_
timestamp 1669390400
transform 1 0 42448 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2236_
timestamp 1669390400
transform 1 0 49840 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2237_
timestamp 1669390400
transform -1 0 48272 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2238_
timestamp 1669390400
transform -1 0 35280 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2239_
timestamp 1669390400
transform -1 0 34608 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2240_
timestamp 1669390400
transform 1 0 39088 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2241_
timestamp 1669390400
transform -1 0 40320 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2242_
timestamp 1669390400
transform 1 0 38752 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2243_
timestamp 1669390400
transform -1 0 41216 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2244_
timestamp 1669390400
transform 1 0 45360 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2245_
timestamp 1669390400
transform -1 0 47376 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2246_
timestamp 1669390400
transform -1 0 57904 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2247_
timestamp 1669390400
transform -1 0 50064 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2248_
timestamp 1669390400
transform 1 0 45696 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2249_
timestamp 1669390400
transform 1 0 57344 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2250_
timestamp 1669390400
transform 1 0 51408 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2251_
timestamp 1669390400
transform -1 0 58128 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2252_
timestamp 1669390400
transform -1 0 54656 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2253_
timestamp 1669390400
transform -1 0 49392 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2254_
timestamp 1669390400
transform 1 0 53872 0 -1 12544
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2255_
timestamp 1669390400
transform 1 0 55776 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2256_
timestamp 1669390400
transform -1 0 56336 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2257_
timestamp 1669390400
transform 1 0 43568 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2258_
timestamp 1669390400
transform 1 0 53312 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2259_
timestamp 1669390400
transform 1 0 44016 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2260_
timestamp 1669390400
transform -1 0 43344 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2261_
timestamp 1669390400
transform -1 0 44240 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2262_
timestamp 1669390400
transform -1 0 43232 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2263_
timestamp 1669390400
transform 1 0 44016 0 -1 20384
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2264_
timestamp 1669390400
transform 1 0 42336 0 -1 21952
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2265_
timestamp 1669390400
transform -1 0 56896 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2266_
timestamp 1669390400
transform 1 0 52080 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2267_
timestamp 1669390400
transform 1 0 56896 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_2  _2268_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 55328 0 -1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2269_
timestamp 1669390400
transform -1 0 53984 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2270_
timestamp 1669390400
transform 1 0 55328 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2271_
timestamp 1669390400
transform 1 0 42448 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2272_
timestamp 1669390400
transform -1 0 51296 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2273_
timestamp 1669390400
transform -1 0 46368 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2274_
timestamp 1669390400
transform 1 0 45360 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2275_
timestamp 1669390400
transform -1 0 43344 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2276_
timestamp 1669390400
transform -1 0 56896 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2277_
timestamp 1669390400
transform 1 0 38976 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2278_
timestamp 1669390400
transform -1 0 58016 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2279_
timestamp 1669390400
transform 1 0 54656 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2280_
timestamp 1669390400
transform 1 0 41888 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2281_
timestamp 1669390400
transform 1 0 43456 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2282_
timestamp 1669390400
transform -1 0 46032 0 -1 34496
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2283_
timestamp 1669390400
transform -1 0 47040 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2284_
timestamp 1669390400
transform 1 0 54096 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2285_
timestamp 1669390400
transform 1 0 55552 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2286_
timestamp 1669390400
transform 1 0 55104 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2287_
timestamp 1669390400
transform 1 0 53312 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2288_
timestamp 1669390400
transform -1 0 56224 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2289_
timestamp 1669390400
transform -1 0 52640 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2290_
timestamp 1669390400
transform -1 0 52080 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2291_
timestamp 1669390400
transform -1 0 54432 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2292_
timestamp 1669390400
transform 1 0 53312 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2293_
timestamp 1669390400
transform 1 0 54208 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2294_
timestamp 1669390400
transform 1 0 55328 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2295_
timestamp 1669390400
transform -1 0 55440 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2296_
timestamp 1669390400
transform -1 0 55216 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _2297_
timestamp 1669390400
transform -1 0 57008 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2298_
timestamp 1669390400
transform -1 0 58240 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2299_
timestamp 1669390400
transform -1 0 57120 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2300_
timestamp 1669390400
transform 1 0 57232 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2301_
timestamp 1669390400
transform 1 0 54880 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2302_
timestamp 1669390400
transform 1 0 51968 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2303_
timestamp 1669390400
transform -1 0 54096 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2304_
timestamp 1669390400
transform -1 0 48384 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2305_
timestamp 1669390400
transform -1 0 38080 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2306_
timestamp 1669390400
transform -1 0 34160 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2307_
timestamp 1669390400
transform -1 0 33040 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2308_
timestamp 1669390400
transform -1 0 2912 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2309_
timestamp 1669390400
transform -1 0 38080 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2310_
timestamp 1669390400
transform 1 0 36848 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2311_
timestamp 1669390400
transform -1 0 57568 0 1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2312_
timestamp 1669390400
transform 1 0 48048 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2313_
timestamp 1669390400
transform 1 0 57344 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2314_
timestamp 1669390400
transform -1 0 50176 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2315_
timestamp 1669390400
transform -1 0 47040 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2316_
timestamp 1669390400
transform -1 0 42560 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2317_
timestamp 1669390400
transform 1 0 38640 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2318_
timestamp 1669390400
transform 1 0 40208 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2319_
timestamp 1669390400
transform -1 0 46704 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2320_
timestamp 1669390400
transform 1 0 48496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2321_
timestamp 1669390400
transform 1 0 49392 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2322_
timestamp 1669390400
transform 1 0 47712 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2323_
timestamp 1669390400
transform 1 0 41440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2324_
timestamp 1669390400
transform 1 0 47600 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2325_
timestamp 1669390400
transform -1 0 48944 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2326_
timestamp 1669390400
transform -1 0 40096 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2327_
timestamp 1669390400
transform 1 0 47376 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2328_
timestamp 1669390400
transform -1 0 50624 0 1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2329_
timestamp 1669390400
transform -1 0 47824 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2330_
timestamp 1669390400
transform 1 0 41440 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2331_
timestamp 1669390400
transform -1 0 53200 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2332_
timestamp 1669390400
transform -1 0 46928 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2333_
timestamp 1669390400
transform -1 0 43456 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _2334_
timestamp 1669390400
transform 1 0 42560 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _2335_
timestamp 1669390400
transform 1 0 37408 0 1 47040
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2336_
timestamp 1669390400
transform 1 0 47264 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2337_
timestamp 1669390400
transform 1 0 46704 0 1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2338_
timestamp 1669390400
transform 1 0 42112 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2339_
timestamp 1669390400
transform 1 0 42336 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2340_
timestamp 1669390400
transform 1 0 51184 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2341_
timestamp 1669390400
transform -1 0 46928 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2342_
timestamp 1669390400
transform -1 0 46592 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2343_
timestamp 1669390400
transform 1 0 53312 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2344_
timestamp 1669390400
transform 1 0 53312 0 1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2345_
timestamp 1669390400
transform -1 0 54544 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2346_
timestamp 1669390400
transform -1 0 50960 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2347_
timestamp 1669390400
transform 1 0 49392 0 -1 17248
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2348_
timestamp 1669390400
transform 1 0 49616 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2349_
timestamp 1669390400
transform 1 0 56112 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2350_
timestamp 1669390400
transform -1 0 57568 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2351_
timestamp 1669390400
transform 1 0 57344 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2352_
timestamp 1669390400
transform 1 0 57344 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2353_
timestamp 1669390400
transform -1 0 57904 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2354_
timestamp 1669390400
transform 1 0 55888 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2355_
timestamp 1669390400
transform -1 0 55776 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2356_
timestamp 1669390400
transform -1 0 54992 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2357_
timestamp 1669390400
transform -1 0 53984 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2358_
timestamp 1669390400
transform -1 0 44352 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2359_
timestamp 1669390400
transform 1 0 50176 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2360_
timestamp 1669390400
transform 1 0 50176 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2361_
timestamp 1669390400
transform -1 0 51184 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2362_
timestamp 1669390400
transform -1 0 46032 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2363_
timestamp 1669390400
transform 1 0 43792 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2364_
timestamp 1669390400
transform -1 0 52864 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2365_
timestamp 1669390400
transform 1 0 43008 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2366_
timestamp 1669390400
transform -1 0 44800 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2367_
timestamp 1669390400
transform 1 0 44240 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2368_
timestamp 1669390400
transform -1 0 45920 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2369_
timestamp 1669390400
transform -1 0 42224 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2370_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 46592 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2371_
timestamp 1669390400
transform -1 0 47488 0 -1 29792
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2372_
timestamp 1669390400
transform 1 0 57008 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2373_
timestamp 1669390400
transform -1 0 42112 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2374_
timestamp 1669390400
transform 1 0 54880 0 -1 14112
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2375_
timestamp 1669390400
transform -1 0 39312 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2376_
timestamp 1669390400
transform 1 0 54992 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2377_
timestamp 1669390400
transform -1 0 55664 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2378_
timestamp 1669390400
transform -1 0 53088 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2379_
timestamp 1669390400
transform 1 0 45360 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2380_
timestamp 1669390400
transform 1 0 39872 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2381_
timestamp 1669390400
transform 1 0 41440 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2382_
timestamp 1669390400
transform -1 0 43792 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2383_
timestamp 1669390400
transform 1 0 47600 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2384_
timestamp 1669390400
transform -1 0 42336 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2385_
timestamp 1669390400
transform -1 0 54768 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _2386_
timestamp 1669390400
transform 1 0 53312 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2387_
timestamp 1669390400
transform 1 0 45808 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2388_
timestamp 1669390400
transform -1 0 54096 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2389_
timestamp 1669390400
transform 1 0 51072 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2390_
timestamp 1669390400
transform 1 0 51968 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2391_
timestamp 1669390400
transform 1 0 43568 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2392_
timestamp 1669390400
transform 1 0 42000 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2393_
timestamp 1669390400
transform 1 0 41440 0 -1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2394_
timestamp 1669390400
transform -1 0 43568 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2395_
timestamp 1669390400
transform -1 0 43904 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2396_
timestamp 1669390400
transform 1 0 43232 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2397_
timestamp 1669390400
transform -1 0 44912 0 1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2398_
timestamp 1669390400
transform -1 0 45920 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2399_
timestamp 1669390400
transform 1 0 55104 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2400_
timestamp 1669390400
transform -1 0 48160 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2401_
timestamp 1669390400
transform -1 0 47712 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2402_
timestamp 1669390400
transform -1 0 48944 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2403_
timestamp 1669390400
transform -1 0 47488 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2404_
timestamp 1669390400
transform 1 0 50288 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2405_
timestamp 1669390400
transform -1 0 49616 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2406_
timestamp 1669390400
transform -1 0 52752 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2407_
timestamp 1669390400
transform 1 0 49952 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2408_
timestamp 1669390400
transform -1 0 50064 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2409_
timestamp 1669390400
transform 1 0 46368 0 -1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2410_
timestamp 1669390400
transform -1 0 30800 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2411_
timestamp 1669390400
transform -1 0 32592 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2412_
timestamp 1669390400
transform 1 0 32816 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2413_
timestamp 1669390400
transform -1 0 40208 0 1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2414_
timestamp 1669390400
transform 1 0 38976 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2415_
timestamp 1669390400
transform -1 0 45920 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2416_
timestamp 1669390400
transform -1 0 44240 0 -1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2417_
timestamp 1669390400
transform 1 0 52416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2418_
timestamp 1669390400
transform 1 0 54768 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2419_
timestamp 1669390400
transform -1 0 51968 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2420_
timestamp 1669390400
transform 1 0 48048 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2421_
timestamp 1669390400
transform 1 0 49504 0 1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2422_
timestamp 1669390400
transform 1 0 47936 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_2  _2423_
timestamp 1669390400
transform 1 0 49392 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2424_
timestamp 1669390400
transform -1 0 58016 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2425_
timestamp 1669390400
transform -1 0 56784 0 -1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2426_
timestamp 1669390400
transform -1 0 56448 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2427_
timestamp 1669390400
transform 1 0 52640 0 -1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2428_
timestamp 1669390400
transform -1 0 54432 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2429_
timestamp 1669390400
transform 1 0 49616 0 1 25088
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2430_
timestamp 1669390400
transform -1 0 50624 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2431_
timestamp 1669390400
transform -1 0 49952 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2432_
timestamp 1669390400
transform -1 0 50288 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_4  _2433_
timestamp 1669390400
transform 1 0 51968 0 -1 29792
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2434_
timestamp 1669390400
transform -1 0 58016 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2435_
timestamp 1669390400
transform 1 0 51520 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2436_
timestamp 1669390400
transform -1 0 51184 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2437_
timestamp 1669390400
transform -1 0 54208 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2438_
timestamp 1669390400
transform -1 0 55888 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2439_
timestamp 1669390400
transform 1 0 48272 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2440_
timestamp 1669390400
transform 1 0 49728 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2441_
timestamp 1669390400
transform -1 0 52864 0 1 29792
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _2442_
timestamp 1669390400
transform -1 0 54432 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2443_
timestamp 1669390400
transform 1 0 54208 0 1 31360
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2444_
timestamp 1669390400
transform 1 0 53312 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2445_
timestamp 1669390400
transform -1 0 55888 0 -1 31360
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2446_
timestamp 1669390400
transform -1 0 50064 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2447_
timestamp 1669390400
transform 1 0 32032 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2448_
timestamp 1669390400
transform 1 0 39984 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2449_
timestamp 1669390400
transform -1 0 48608 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2450_
timestamp 1669390400
transform -1 0 45136 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2451_
timestamp 1669390400
transform -1 0 48384 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2452_
timestamp 1669390400
transform -1 0 48048 0 1 51744
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2453_
timestamp 1669390400
transform 1 0 46704 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2454_
timestamp 1669390400
transform -1 0 35280 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2455_
timestamp 1669390400
transform 1 0 33488 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2456_
timestamp 1669390400
transform 1 0 49504 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2457_
timestamp 1669390400
transform 1 0 46928 0 -1 31360
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2458_
timestamp 1669390400
transform -1 0 53984 0 -1 23520
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2459_
timestamp 1669390400
transform 1 0 48160 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2460_
timestamp 1669390400
transform 1 0 39088 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2461_
timestamp 1669390400
transform -1 0 47936 0 1 28224
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _2462_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 49952 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2463_
timestamp 1669390400
transform 1 0 33488 0 -1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2464_
timestamp 1669390400
transform -1 0 44576 0 1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2465_
timestamp 1669390400
transform 1 0 43456 0 -1 53312
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2466_
timestamp 1669390400
transform -1 0 44240 0 -1 54880
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2467_
timestamp 1669390400
transform 1 0 42000 0 -1 54880
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2468_
timestamp 1669390400
transform 1 0 40320 0 -1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2469_
timestamp 1669390400
transform -1 0 40544 0 1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2470_
timestamp 1669390400
transform -1 0 2912 0 1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2471_
timestamp 1669390400
transform -1 0 39424 0 -1 53312
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2472_
timestamp 1669390400
transform -1 0 46704 0 1 51744
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2473_
timestamp 1669390400
transform -1 0 43008 0 1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2474_
timestamp 1669390400
transform 1 0 39088 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2475_
timestamp 1669390400
transform 1 0 48832 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2476_
timestamp 1669390400
transform 1 0 49392 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2477_
timestamp 1669390400
transform 1 0 49952 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2478_
timestamp 1669390400
transform 1 0 46368 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2479_
timestamp 1669390400
transform 1 0 47264 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2480_
timestamp 1669390400
transform -1 0 48272 0 -1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2481_
timestamp 1669390400
transform -1 0 47600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2482_
timestamp 1669390400
transform 1 0 47600 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2483_
timestamp 1669390400
transform 1 0 51408 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2484_
timestamp 1669390400
transform 1 0 51184 0 1 15680
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2485_
timestamp 1669390400
transform -1 0 53984 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2486_
timestamp 1669390400
transform 1 0 53312 0 1 25088
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2487_
timestamp 1669390400
transform 1 0 52640 0 -1 28224
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _2488_
timestamp 1669390400
transform -1 0 54768 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2489_
timestamp 1669390400
transform 1 0 53312 0 1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2490_
timestamp 1669390400
transform -1 0 53200 0 -1 47040
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2491_
timestamp 1669390400
transform -1 0 45920 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2492_
timestamp 1669390400
transform 1 0 42672 0 -1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2493_
timestamp 1669390400
transform 1 0 41328 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2494_
timestamp 1669390400
transform 1 0 53312 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2495_
timestamp 1669390400
transform 1 0 56000 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2496_
timestamp 1669390400
transform -1 0 56560 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2497_
timestamp 1669390400
transform -1 0 52640 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2498_
timestamp 1669390400
transform 1 0 51744 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2499_
timestamp 1669390400
transform 1 0 52304 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2500_
timestamp 1669390400
transform -1 0 50288 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2501_
timestamp 1669390400
transform 1 0 50512 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2502_
timestamp 1669390400
transform 1 0 51632 0 1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2503_
timestamp 1669390400
transform -1 0 52752 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2504_
timestamp 1669390400
transform -1 0 46480 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2505_
timestamp 1669390400
transform -1 0 44912 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2506_
timestamp 1669390400
transform 1 0 45136 0 -1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2507_
timestamp 1669390400
transform 1 0 47600 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2508_
timestamp 1669390400
transform -1 0 48496 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2509_
timestamp 1669390400
transform 1 0 46144 0 1 45472
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2510_
timestamp 1669390400
transform 1 0 39984 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2511_
timestamp 1669390400
transform -1 0 41440 0 1 47040
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2512_
timestamp 1669390400
transform 1 0 39872 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2513_
timestamp 1669390400
transform 1 0 39872 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2514_
timestamp 1669390400
transform 1 0 51184 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2515_
timestamp 1669390400
transform 1 0 39648 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2516_
timestamp 1669390400
transform -1 0 47152 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2517_
timestamp 1669390400
transform 1 0 39648 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2518_
timestamp 1669390400
transform 1 0 39984 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_2  _2519_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 40544 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2520_
timestamp 1669390400
transform -1 0 32816 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2521_
timestamp 1669390400
transform 1 0 33040 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2522_
timestamp 1669390400
transform 1 0 39648 0 -1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2523_
timestamp 1669390400
transform 1 0 39760 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2524_
timestamp 1669390400
transform 1 0 40432 0 -1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2525_
timestamp 1669390400
transform 1 0 40880 0 -1 56448
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2526_
timestamp 1669390400
transform 1 0 41776 0 1 54880
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2527_
timestamp 1669390400
transform 1 0 46480 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2528_
timestamp 1669390400
transform 1 0 39872 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2529_
timestamp 1669390400
transform 1 0 39984 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2530_
timestamp 1669390400
transform -1 0 40656 0 -1 51744
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2531_
timestamp 1669390400
transform -1 0 52304 0 1 47040
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2532_
timestamp 1669390400
transform 1 0 50064 0 1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2533_
timestamp 1669390400
transform 1 0 51296 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2534_
timestamp 1669390400
transform 1 0 43456 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2535_
timestamp 1669390400
transform 1 0 49504 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2536_
timestamp 1669390400
transform -1 0 52304 0 -1 36064
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2537_
timestamp 1669390400
transform -1 0 51632 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2538_
timestamp 1669390400
transform 1 0 49280 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2539_
timestamp 1669390400
transform -1 0 49168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2540_
timestamp 1669390400
transform -1 0 50400 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2541_
timestamp 1669390400
transform 1 0 50176 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2542_
timestamp 1669390400
transform 1 0 50176 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2543_
timestamp 1669390400
transform -1 0 44128 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2544_
timestamp 1669390400
transform 1 0 41440 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2545_
timestamp 1669390400
transform -1 0 47712 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2546_
timestamp 1669390400
transform -1 0 49504 0 1 18816
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2547_
timestamp 1669390400
transform -1 0 50176 0 -1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2548_
timestamp 1669390400
transform -1 0 47488 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2549_
timestamp 1669390400
transform 1 0 47824 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2550_
timestamp 1669390400
transform -1 0 55104 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2551_
timestamp 1669390400
transform 1 0 53872 0 1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2552_
timestamp 1669390400
transform 1 0 48048 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2553_
timestamp 1669390400
transform -1 0 48944 0 1 31360
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2554_
timestamp 1669390400
transform 1 0 47152 0 -1 37632
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2555_
timestamp 1669390400
transform -1 0 52864 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2556_
timestamp 1669390400
transform 1 0 46144 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2557_
timestamp 1669390400
transform -1 0 41776 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2558_
timestamp 1669390400
transform 1 0 42336 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2559_
timestamp 1669390400
transform 1 0 43680 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2560_
timestamp 1669390400
transform 1 0 40320 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2561_
timestamp 1669390400
transform 1 0 41440 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2562_
timestamp 1669390400
transform 1 0 45472 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2563_
timestamp 1669390400
transform -1 0 47040 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2564_
timestamp 1669390400
transform 1 0 43904 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2565_
timestamp 1669390400
transform 1 0 44688 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2566_
timestamp 1669390400
transform -1 0 45584 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2567_
timestamp 1669390400
transform -1 0 45360 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2568_
timestamp 1669390400
transform 1 0 43904 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2569_
timestamp 1669390400
transform -1 0 45584 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2570_
timestamp 1669390400
transform 1 0 43792 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2571_
timestamp 1669390400
transform -1 0 44912 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2572_
timestamp 1669390400
transform 1 0 49392 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2573_
timestamp 1669390400
transform 1 0 45024 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2574_
timestamp 1669390400
transform -1 0 46256 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2575_
timestamp 1669390400
transform -1 0 45472 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2576_
timestamp 1669390400
transform 1 0 42560 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2577_
timestamp 1669390400
transform -1 0 44688 0 1 47040
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2578_
timestamp 1669390400
transform 1 0 47152 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2579_
timestamp 1669390400
transform 1 0 48160 0 1 34496
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2580_
timestamp 1669390400
transform 1 0 47712 0 1 36064
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2581_
timestamp 1669390400
transform -1 0 49168 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2582_
timestamp 1669390400
transform -1 0 48048 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2583_
timestamp 1669390400
transform -1 0 44576 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2584_
timestamp 1669390400
transform -1 0 43008 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2585_
timestamp 1669390400
transform 1 0 43904 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2586_
timestamp 1669390400
transform 1 0 42336 0 -1 45472
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2587_
timestamp 1669390400
transform 1 0 38080 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2588_
timestamp 1669390400
transform -1 0 38080 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2589_
timestamp 1669390400
transform -1 0 40096 0 1 18816
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2590_
timestamp 1669390400
transform 1 0 34608 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2591_
timestamp 1669390400
transform 1 0 35728 0 1 18816
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2592_
timestamp 1669390400
transform 1 0 36624 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2593_
timestamp 1669390400
transform -1 0 43792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2594_
timestamp 1669390400
transform -1 0 38640 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2595_
timestamp 1669390400
transform 1 0 37520 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2596_
timestamp 1669390400
transform -1 0 33936 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2597_
timestamp 1669390400
transform -1 0 37632 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2598_
timestamp 1669390400
transform -1 0 36176 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2599_
timestamp 1669390400
transform 1 0 33488 0 -1 31360
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2600_
timestamp 1669390400
transform 1 0 33152 0 1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor3_1  _2601_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 37856 0 -1 51744
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2602_
timestamp 1669390400
transform 1 0 42448 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2603_
timestamp 1669390400
transform 1 0 38864 0 1 53312
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2604_
timestamp 1669390400
transform 1 0 41440 0 -1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2605_
timestamp 1669390400
transform -1 0 43568 0 1 53312
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _2606_
timestamp 1669390400
transform 1 0 39984 0 1 53312
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2607_
timestamp 1669390400
transform -1 0 35280 0 1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2608_
timestamp 1669390400
transform 1 0 33488 0 -1 51744
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2609_
timestamp 1669390400
transform 1 0 33712 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2610_
timestamp 1669390400
transform -1 0 43680 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2611_
timestamp 1669390400
transform 1 0 35392 0 -1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2612_
timestamp 1669390400
transform -1 0 39648 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2613_
timestamp 1669390400
transform -1 0 39984 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_4  _2614_
timestamp 1669390400
transform -1 0 40992 0 1 29792
box -86 -86 2774 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2615_
timestamp 1669390400
transform -1 0 43120 0 -1 34496
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2616_
timestamp 1669390400
transform -1 0 41104 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2617_
timestamp 1669390400
transform 1 0 38304 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2618_
timestamp 1669390400
transform 1 0 38976 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2619_
timestamp 1669390400
transform -1 0 38976 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2620_
timestamp 1669390400
transform -1 0 40992 0 -1 36064
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2621_
timestamp 1669390400
transform 1 0 39760 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _2622_
timestamp 1669390400
transform -1 0 40992 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_4  _2623_
timestamp 1669390400
transform -1 0 43568 0 1 34496
box -86 -86 3782 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2624_
timestamp 1669390400
transform 1 0 51744 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2625_
timestamp 1669390400
transform 1 0 53312 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2626_
timestamp 1669390400
transform 1 0 53536 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2627_
timestamp 1669390400
transform -1 0 50848 0 -1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2628_
timestamp 1669390400
transform -1 0 47824 0 -1 40768
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2629_
timestamp 1669390400
transform -1 0 47712 0 -1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2630_
timestamp 1669390400
transform 1 0 46032 0 1 47040
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2631_
timestamp 1669390400
transform -1 0 50848 0 1 48608
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2632_
timestamp 1669390400
transform 1 0 49392 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2633_
timestamp 1669390400
transform -1 0 48944 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2634_
timestamp 1669390400
transform 1 0 46592 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2635_
timestamp 1669390400
transform 1 0 39088 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2636_
timestamp 1669390400
transform 1 0 46032 0 1 48608
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2637_
timestamp 1669390400
transform -1 0 31808 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2638_
timestamp 1669390400
transform -1 0 38864 0 -1 28224
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2639_
timestamp 1669390400
transform 1 0 36176 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2640_
timestamp 1669390400
transform -1 0 38640 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2641_
timestamp 1669390400
transform -1 0 38528 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2642_
timestamp 1669390400
transform -1 0 36960 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2643_
timestamp 1669390400
transform 1 0 35840 0 -1 29792
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _2644_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 36960 0 1 29792
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2645_
timestamp 1669390400
transform -1 0 32032 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2646_
timestamp 1669390400
transform 1 0 29120 0 -1 31360
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2647_
timestamp 1669390400
transform 1 0 29232 0 -1 50176
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _2648_
timestamp 1669390400
transform -1 0 36960 0 1 50176
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2649_
timestamp 1669390400
transform 1 0 35728 0 1 51744
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2650_
timestamp 1669390400
transform -1 0 36624 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2651_
timestamp 1669390400
transform 1 0 33488 0 -1 53312
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2652_
timestamp 1669390400
transform 1 0 31584 0 -1 51744
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2653_
timestamp 1669390400
transform -1 0 57680 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2654_
timestamp 1669390400
transform 1 0 47488 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2655_
timestamp 1669390400
transform 1 0 29904 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2656_
timestamp 1669390400
transform -1 0 39536 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2657_
timestamp 1669390400
transform -1 0 50848 0 -1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2658_
timestamp 1669390400
transform -1 0 52304 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2659_
timestamp 1669390400
transform -1 0 33040 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2660_
timestamp 1669390400
transform 1 0 34384 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2661_
timestamp 1669390400
transform -1 0 36960 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2662_
timestamp 1669390400
transform 1 0 37408 0 1 25088
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2663_
timestamp 1669390400
transform -1 0 38080 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2664_
timestamp 1669390400
transform 1 0 36960 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2665_
timestamp 1669390400
transform -1 0 39536 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2666_
timestamp 1669390400
transform -1 0 33712 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2667_
timestamp 1669390400
transform -1 0 38416 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2668_
timestamp 1669390400
transform 1 0 38864 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2669_
timestamp 1669390400
transform -1 0 41552 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2670_
timestamp 1669390400
transform -1 0 40208 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2671_
timestamp 1669390400
transform 1 0 37632 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2672_
timestamp 1669390400
transform -1 0 51856 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2673_
timestamp 1669390400
transform 1 0 38528 0 1 40768
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2674_
timestamp 1669390400
transform -1 0 44240 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2675_
timestamp 1669390400
transform 1 0 40656 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2676_
timestamp 1669390400
transform -1 0 42672 0 -1 18816
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2677_
timestamp 1669390400
transform 1 0 41776 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2678_
timestamp 1669390400
transform 1 0 40208 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2679_
timestamp 1669390400
transform -1 0 40992 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2680_
timestamp 1669390400
transform 1 0 42336 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2681_
timestamp 1669390400
transform 1 0 41888 0 -1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2682_
timestamp 1669390400
transform 1 0 43344 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2683_
timestamp 1669390400
transform 1 0 45360 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2684_
timestamp 1669390400
transform 1 0 45696 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2685_
timestamp 1669390400
transform 1 0 45360 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2686_
timestamp 1669390400
transform 1 0 45920 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2687_
timestamp 1669390400
transform 1 0 45584 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2688_
timestamp 1669390400
transform -1 0 39536 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2689_
timestamp 1669390400
transform -1 0 40656 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2690_
timestamp 1669390400
transform -1 0 40432 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2691_
timestamp 1669390400
transform -1 0 47040 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2692_
timestamp 1669390400
transform 1 0 39872 0 -1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2693_
timestamp 1669390400
transform -1 0 39536 0 1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2694_
timestamp 1669390400
transform -1 0 31472 0 -1 29792
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2695_
timestamp 1669390400
transform -1 0 35840 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2696_
timestamp 1669390400
transform -1 0 36288 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2697_
timestamp 1669390400
transform 1 0 37408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2698_
timestamp 1669390400
transform -1 0 36400 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2699_
timestamp 1669390400
transform 1 0 34384 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2700_
timestamp 1669390400
transform -1 0 33040 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2701_
timestamp 1669390400
transform -1 0 32704 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2702_
timestamp 1669390400
transform 1 0 30688 0 -1 23520
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2703_
timestamp 1669390400
transform -1 0 33040 0 -1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2704_
timestamp 1669390400
transform -1 0 30688 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _2705_
timestamp 1669390400
transform -1 0 34160 0 1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2706_
timestamp 1669390400
transform 1 0 32032 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2707_
timestamp 1669390400
transform 1 0 30352 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2708_
timestamp 1669390400
transform 1 0 32368 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2709_
timestamp 1669390400
transform -1 0 34384 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2710_
timestamp 1669390400
transform 1 0 33488 0 -1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2711_
timestamp 1669390400
transform -1 0 34048 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2712_
timestamp 1669390400
transform 1 0 34720 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2713_
timestamp 1669390400
transform 1 0 33152 0 1 48608
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2714_
timestamp 1669390400
transform -1 0 30128 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2715_
timestamp 1669390400
transform 1 0 29456 0 1 45472
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2716_
timestamp 1669390400
transform -1 0 58016 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2717_
timestamp 1669390400
transform 1 0 32592 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2718_
timestamp 1669390400
transform -1 0 42224 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_2  _2719_
timestamp 1669390400
transform 1 0 39872 0 1 26656
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _2720_
timestamp 1669390400
transform 1 0 45696 0 -1 28224
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2721_
timestamp 1669390400
transform -1 0 43232 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2722_
timestamp 1669390400
transform -1 0 43456 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2723_
timestamp 1669390400
transform -1 0 42336 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2724_
timestamp 1669390400
transform -1 0 44464 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2725_
timestamp 1669390400
transform 1 0 42560 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2726_
timestamp 1669390400
transform -1 0 44912 0 1 28224
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2727_
timestamp 1669390400
transform -1 0 43120 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2728_
timestamp 1669390400
transform 1 0 41440 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2729_
timestamp 1669390400
transform -1 0 35280 0 -1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2730_
timestamp 1669390400
transform -1 0 38304 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2731_
timestamp 1669390400
transform -1 0 36512 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2732_
timestamp 1669390400
transform 1 0 35280 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2733_
timestamp 1669390400
transform -1 0 35056 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2734_
timestamp 1669390400
transform 1 0 37408 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2735_
timestamp 1669390400
transform -1 0 36960 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2736_
timestamp 1669390400
transform -1 0 38640 0 1 42336
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2737_
timestamp 1669390400
transform 1 0 36624 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2738_
timestamp 1669390400
transform 1 0 31136 0 -1 42336
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _2739_
timestamp 1669390400
transform -1 0 34944 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2740_
timestamp 1669390400
transform -1 0 34832 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2741_
timestamp 1669390400
transform -1 0 34048 0 1 23520
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2742_
timestamp 1669390400
transform -1 0 35392 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _2743_
timestamp 1669390400
transform -1 0 34048 0 1 20384
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2744_
timestamp 1669390400
transform -1 0 33040 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2745_
timestamp 1669390400
transform 1 0 30464 0 1 23520
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2746_
timestamp 1669390400
transform -1 0 32144 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2747_
timestamp 1669390400
transform 1 0 32368 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2748_
timestamp 1669390400
transform -1 0 30800 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2749_
timestamp 1669390400
transform 1 0 30800 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2750_
timestamp 1669390400
transform -1 0 30576 0 1 43904
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _2751_
timestamp 1669390400
transform 1 0 29568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2752_
timestamp 1669390400
transform 1 0 28112 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2753_
timestamp 1669390400
transform 1 0 27664 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2754_
timestamp 1669390400
transform -1 0 28560 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2755_
timestamp 1669390400
transform -1 0 32032 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2756_
timestamp 1669390400
transform 1 0 28448 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2757_
timestamp 1669390400
transform 1 0 39984 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2758_
timestamp 1669390400
transform 1 0 37408 0 1 20384
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _2759_
timestamp 1669390400
transform 1 0 35616 0 1 21952
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2760_
timestamp 1669390400
transform -1 0 42112 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2761_
timestamp 1669390400
transform 1 0 35728 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2762_
timestamp 1669390400
transform -1 0 35952 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2763_
timestamp 1669390400
transform -1 0 36624 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2764_
timestamp 1669390400
transform -1 0 45584 0 -1 42336
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2765_
timestamp 1669390400
transform -1 0 36624 0 1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2766_
timestamp 1669390400
transform -1 0 39760 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2767_
timestamp 1669390400
transform -1 0 38640 0 -1 34496
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2768_
timestamp 1669390400
transform -1 0 38640 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2769_
timestamp 1669390400
transform -1 0 37968 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2770_
timestamp 1669390400
transform 1 0 37968 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2771_
timestamp 1669390400
transform -1 0 34048 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2772_
timestamp 1669390400
transform -1 0 34160 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2773_
timestamp 1669390400
transform -1 0 36064 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2774_
timestamp 1669390400
transform -1 0 32816 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2775_
timestamp 1669390400
transform -1 0 34720 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2776_
timestamp 1669390400
transform -1 0 38080 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2777_
timestamp 1669390400
transform -1 0 34944 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _2778_
timestamp 1669390400
transform -1 0 32704 0 -1 26656
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2779_
timestamp 1669390400
transform -1 0 31584 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2780_
timestamp 1669390400
transform -1 0 29008 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _2781_
timestamp 1669390400
transform 1 0 35504 0 -1 31360
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2782_
timestamp 1669390400
transform -1 0 29792 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2783_
timestamp 1669390400
transform -1 0 31136 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2784_
timestamp 1669390400
transform 1 0 29456 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2785_
timestamp 1669390400
transform -1 0 31808 0 -1 40768
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2786_
timestamp 1669390400
transform -1 0 29568 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2787_
timestamp 1669390400
transform 1 0 29904 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2788_
timestamp 1669390400
transform -1 0 31360 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_4  _2789_
timestamp 1669390400
transform 1 0 28000 0 -1 43904
box -86 -86 4118 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2790_
timestamp 1669390400
transform -1 0 28000 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2791_
timestamp 1669390400
transform -1 0 2912 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2792_
timestamp 1669390400
transform -1 0 34608 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _2793_
timestamp 1669390400
transform -1 0 32480 0 1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2794_
timestamp 1669390400
transform -1 0 44240 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _2795_
timestamp 1669390400
transform -1 0 40208 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _2796_
timestamp 1669390400
transform 1 0 35280 0 -1 32928
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2797_
timestamp 1669390400
transform -1 0 35504 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2798_
timestamp 1669390400
transform 1 0 35504 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2799_
timestamp 1669390400
transform -1 0 35840 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2800_
timestamp 1669390400
transform -1 0 34496 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2801_
timestamp 1669390400
transform 1 0 35168 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2802_
timestamp 1669390400
transform -1 0 36512 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2803_
timestamp 1669390400
transform -1 0 36176 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2804_
timestamp 1669390400
transform 1 0 36624 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _2805_
timestamp 1669390400
transform -1 0 36400 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2806_
timestamp 1669390400
transform -1 0 35504 0 1 37632
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2807_
timestamp 1669390400
transform -1 0 34832 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2808_
timestamp 1669390400
transform -1 0 32480 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2809_
timestamp 1669390400
transform -1 0 31584 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2810_
timestamp 1669390400
transform 1 0 30016 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2811_
timestamp 1669390400
transform -1 0 31472 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2812_
timestamp 1669390400
transform -1 0 32256 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2813_
timestamp 1669390400
transform -1 0 30128 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2814_
timestamp 1669390400
transform 1 0 29456 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2815_
timestamp 1669390400
transform 1 0 29456 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2816_
timestamp 1669390400
transform -1 0 27776 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2817_
timestamp 1669390400
transform -1 0 28896 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2818_
timestamp 1669390400
transform -1 0 27328 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2819_
timestamp 1669390400
transform 1 0 40208 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2820_
timestamp 1669390400
transform 1 0 49392 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _2821_
timestamp 1669390400
transform -1 0 38528 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2822_
timestamp 1669390400
transform 1 0 38080 0 -1 36064
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2823_
timestamp 1669390400
transform 1 0 53088 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2824_
timestamp 1669390400
transform -1 0 54320 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2825_
timestamp 1669390400
transform -1 0 36624 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2826_
timestamp 1669390400
transform 1 0 35952 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _2827_
timestamp 1669390400
transform -1 0 36960 0 1 37632
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _2828_
timestamp 1669390400
transform 1 0 38416 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2829_
timestamp 1669390400
transform -1 0 56336 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2830_
timestamp 1669390400
transform 1 0 30800 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _2831_
timestamp 1669390400
transform 1 0 53872 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2832_
timestamp 1669390400
transform -1 0 57008 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2833_
timestamp 1669390400
transform 1 0 32480 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2834_
timestamp 1669390400
transform -1 0 34272 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _2835_
timestamp 1669390400
transform -1 0 56896 0 1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2836_
timestamp 1669390400
transform 1 0 56000 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2837_
timestamp 1669390400
transform -1 0 31248 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2838_
timestamp 1669390400
transform -1 0 32032 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2839_
timestamp 1669390400
transform -1 0 30352 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _2840_
timestamp 1669390400
transform -1 0 30800 0 -1 39200
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2841_
timestamp 1669390400
transform -1 0 57792 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2842_
timestamp 1669390400
transform -1 0 56448 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2843_
timestamp 1669390400
transform 1 0 53760 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2844_
timestamp 1669390400
transform -1 0 55440 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _2845_
timestamp 1669390400
transform 1 0 38416 0 1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2846_
timestamp 1669390400
transform 1 0 48048 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2847_
timestamp 1669390400
transform -1 0 48944 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2848_
timestamp 1669390400
transform 1 0 48832 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _2849_
timestamp 1669390400
transform -1 0 51184 0 -1 42336
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _2850_
timestamp 1669390400
transform 1 0 53312 0 1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2851_
timestamp 1669390400
transform 1 0 55552 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2852_
timestamp 1669390400
transform 1 0 55888 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2853_
timestamp 1669390400
transform -1 0 58240 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2854_
timestamp 1669390400
transform -1 0 58016 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2855_
timestamp 1669390400
transform -1 0 58016 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2856_
timestamp 1669390400
transform -1 0 55216 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2857_
timestamp 1669390400
transform -1 0 58016 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2858_
timestamp 1669390400
transform 1 0 54880 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2859_
timestamp 1669390400
transform -1 0 57904 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2860_
timestamp 1669390400
transform 1 0 55552 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2861_
timestamp 1669390400
transform 1 0 54768 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2862_
timestamp 1669390400
transform 1 0 55104 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2863_
timestamp 1669390400
transform 1 0 56112 0 1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2864_
timestamp 1669390400
transform 1 0 56000 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2865_
timestamp 1669390400
transform 1 0 56672 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2866_
timestamp 1669390400
transform -1 0 38752 0 -1 54880
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2867_
timestamp 1669390400
transform -1 0 38080 0 1 54880
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2868_
timestamp 1669390400
transform -1 0 40432 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2869_
timestamp 1669390400
transform 1 0 38528 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2870_
timestamp 1669390400
transform -1 0 35280 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2871_
timestamp 1669390400
transform 1 0 34496 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _2872_
timestamp 1669390400
transform -1 0 34272 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2873_
timestamp 1669390400
transform -1 0 33712 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2874_
timestamp 1669390400
transform 1 0 33712 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2875_
timestamp 1669390400
transform 1 0 33264 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2876_
timestamp 1669390400
transform 1 0 37408 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2877_
timestamp 1669390400
transform 1 0 41440 0 1 12544
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2878_
timestamp 1669390400
transform 1 0 43120 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2879_
timestamp 1669390400
transform 1 0 38864 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2880_
timestamp 1669390400
transform -1 0 41216 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2881_
timestamp 1669390400
transform -1 0 40992 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2882_
timestamp 1669390400
transform 1 0 36176 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _2883_
timestamp 1669390400
transform 1 0 37744 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2884_
timestamp 1669390400
transform -1 0 37520 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _2885_
timestamp 1669390400
transform 1 0 37520 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _2886_
timestamp 1669390400
transform 1 0 36064 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2887_
timestamp 1669390400
transform 1 0 37520 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2888_
timestamp 1669390400
transform -1 0 36624 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _2889_
timestamp 1669390400
transform 1 0 35504 0 1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2890_
timestamp 1669390400
transform -1 0 33152 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _2891_
timestamp 1669390400
transform 1 0 35168 0 -1 17248
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _2892_
timestamp 1669390400
transform 1 0 33376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _2893_
timestamp 1669390400
transform -1 0 34608 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2894_
timestamp 1669390400
transform -1 0 35840 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _2895_
timestamp 1669390400
transform 1 0 35168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2896_
timestamp 1669390400
transform -1 0 32256 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2897_
timestamp 1669390400
transform -1 0 34048 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _2898_
timestamp 1669390400
transform 1 0 32144 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2899_
timestamp 1669390400
transform 1 0 29904 0 1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2900_
timestamp 1669390400
transform 1 0 29344 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _2901_
timestamp 1669390400
transform -1 0 31024 0 -1 15680
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _2902_
timestamp 1669390400
transform -1 0 32928 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2903_
timestamp 1669390400
transform -1 0 31472 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2904_
timestamp 1669390400
transform -1 0 32816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _2905_
timestamp 1669390400
transform 1 0 32032 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _2906_
timestamp 1669390400
transform 1 0 30688 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2907_
timestamp 1669390400
transform -1 0 6272 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2908_
timestamp 1669390400
transform -1 0 6160 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2909_
timestamp 1669390400
transform 1 0 34384 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _2910_
timestamp 1669390400
transform 1 0 35504 0 -1 12544
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _2911_
timestamp 1669390400
transform 1 0 35616 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2912_
timestamp 1669390400
transform -1 0 37968 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _2913_
timestamp 1669390400
transform -1 0 36624 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2914_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 45584 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2915_
timestamp 1669390400
transform 1 0 37184 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2916_
timestamp 1669390400
transform 1 0 38080 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2917_
timestamp 1669390400
transform -1 0 53200 0 -1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2918_
timestamp 1669390400
transform 1 0 45360 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2919_
timestamp 1669390400
transform 1 0 45360 0 1 7840
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2920_
timestamp 1669390400
transform 1 0 45360 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2921_
timestamp 1669390400
transform 1 0 45360 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2922_
timestamp 1669390400
transform 1 0 49392 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2923_
timestamp 1669390400
transform 1 0 37408 0 1 4704
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2924_
timestamp 1669390400
transform 1 0 41440 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2925_
timestamp 1669390400
transform 1 0 37184 0 -1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2926_
timestamp 1669390400
transform 1 0 38192 0 1 6272
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2927_
timestamp 1669390400
transform 1 0 38080 0 1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2928_
timestamp 1669390400
transform 1 0 44800 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2929_
timestamp 1669390400
transform 1 0 2576 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2930_
timestamp 1669390400
transform 1 0 5264 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2931_
timestamp 1669390400
transform 1 0 49056 0 1 39200
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2932_ dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 29456 0 1 34496
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2933_
timestamp 1669390400
transform 1 0 49504 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2934_
timestamp 1669390400
transform 1 0 37968 0 1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2935_
timestamp 1669390400
transform 1 0 21168 0 -1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__latrnq_1  _2936_
timestamp 1669390400
transform 1 0 25872 0 1 31360
box -86 -86 2550 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2937_
timestamp 1669390400
transform -1 0 28112 0 1 34496
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2938_
timestamp 1669390400
transform 1 0 33488 0 -1 45472
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _2939_
timestamp 1669390400
transform 1 0 35840 0 -1 43904
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_CLK dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 47040 0 -1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_CLK
timestamp 1669390400
transform -1 0 39760 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_CLK
timestamp 1669390400
transform 1 0 41776 0 -1 4704
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout42
timestamp 1669390400
transform 1 0 40320 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout43 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 36960 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout44
timestamp 1669390400
transform -1 0 29120 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout45
timestamp 1669390400
transform 1 0 29344 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout46
timestamp 1669390400
transform 1 0 28000 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout47 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform 1 0 53536 0 -1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout48
timestamp 1669390400
transform -1 0 10304 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout49
timestamp 1669390400
transform 1 0 24192 0 1 32928
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout50
timestamp 1669390400
transform 1 0 8512 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout51
timestamp 1669390400
transform -1 0 45472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout52
timestamp 1669390400
transform -1 0 42672 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  fanout53
timestamp 1669390400
transform 1 0 45472 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout54
timestamp 1669390400
transform 1 0 47600 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout55
timestamp 1669390400
transform -1 0 52192 0 1 9408
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout56
timestamp 1669390400
transform 1 0 42224 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  fanout57
timestamp 1669390400
transform 1 0 31360 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  fanout58
timestamp 1669390400
transform 1 0 41552 0 1 4704
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  fanout59
timestamp 1669390400
transform 1 0 42336 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input1
timestamp 1669390400
transform 1 0 1680 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__dlyc_1  input2
timestamp 1669390400
transform 1 0 31696 0 1 54880
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__dlyb_1  input3
timestamp 1669390400
transform 1 0 5600 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output4 dependencies/pdks/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1669390400
transform -1 0 3248 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output5
timestamp 1669390400
transform -1 0 56112 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output6
timestamp 1669390400
transform -1 0 56336 0 -1 4704
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output7
timestamp 1669390400
transform -1 0 56560 0 -1 37632
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output8
timestamp 1669390400
transform -1 0 4368 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output9
timestamp 1669390400
transform -1 0 3248 0 1 51744
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output10
timestamp 1669390400
transform 1 0 48720 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output11
timestamp 1669390400
transform 1 0 34384 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output12
timestamp 1669390400
transform -1 0 56336 0 -1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output13
timestamp 1669390400
transform -1 0 56336 0 1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output14
timestamp 1669390400
transform -1 0 12992 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output15
timestamp 1669390400
transform -1 0 3248 0 -1 40768
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output16
timestamp 1669390400
transform -1 0 3248 0 1 28224
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output17
timestamp 1669390400
transform 1 0 37072 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output18
timestamp 1669390400
transform 1 0 54544 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output19
timestamp 1669390400
transform -1 0 3248 0 1 34496
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output20
timestamp 1669390400
transform 1 0 54768 0 1 48608
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output21
timestamp 1669390400
transform 1 0 14224 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output22
timestamp 1669390400
transform -1 0 3248 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output23
timestamp 1669390400
transform -1 0 3248 0 -1 12544
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output24
timestamp 1669390400
transform 1 0 54768 0 -1 32928
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output25
timestamp 1669390400
transform -1 0 9072 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output26
timestamp 1669390400
transform -1 0 3248 0 -1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output27
timestamp 1669390400
transform 1 0 52640 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output28
timestamp 1669390400
transform 1 0 42784 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output29
timestamp 1669390400
transform -1 0 56336 0 1 14112
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output30
timestamp 1669390400
transform -1 0 18928 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output31
timestamp 1669390400
transform -1 0 24528 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output32
timestamp 1669390400
transform 1 0 54768 0 1 20384
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output33
timestamp 1669390400
transform -1 0 30688 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output34
timestamp 1669390400
transform 1 0 54768 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output35
timestamp 1669390400
transform 1 0 56560 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output36
timestamp 1669390400
transform -1 0 20832 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output37
timestamp 1669390400
transform -1 0 27216 0 -1 56448
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output38
timestamp 1669390400
transform 1 0 38864 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output39
timestamp 1669390400
transform -1 0 3248 0 1 21952
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output40
timestamp 1669390400
transform -1 0 3248 0 1 54880
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  output41
timestamp 1669390400
transform 1 0 54768 0 -1 26656
box -86 -86 1654 870
<< labels >>
flabel metal3 s 200 16800 800 16912 0 FreeSans 448 0 0 0 BitIn
port 0 nsew signal input
flabel metal2 s 45696 200 45808 800 0 FreeSans 448 90 0 0 CLK
port 1 nsew signal input
flabel metal2 s 31584 59200 31696 59800 0 FreeSans 448 90 0 0 EN
port 2 nsew signal input
flabel metal3 s 200 45696 800 45808 0 FreeSans 448 0 0 0 I[0]
port 3 nsew signal tristate
flabel metal2 s 57120 200 57232 800 0 FreeSans 448 90 0 0 I[10]
port 4 nsew signal tristate
flabel metal3 s 59200 2688 59800 2800 0 FreeSans 448 0 0 0 I[11]
port 5 nsew signal tristate
flabel metal3 s 59200 36960 59800 37072 0 FreeSans 448 0 0 0 I[12]
port 6 nsew signal tristate
flabel metal2 s 2688 59200 2800 59800 0 FreeSans 448 90 0 0 I[1]
port 7 nsew signal tristate
flabel metal3 s 200 51744 800 51856 0 FreeSans 448 0 0 0 I[2]
port 8 nsew signal tristate
flabel metal2 s 48384 59200 48496 59800 0 FreeSans 448 90 0 0 I[3]
port 9 nsew signal tristate
flabel metal2 s 34272 200 34384 800 0 FreeSans 448 90 0 0 I[4]
port 10 nsew signal tristate
flabel metal3 s 59200 43008 59800 43120 0 FreeSans 448 0 0 0 I[5]
port 11 nsew signal tristate
flabel metal3 s 59200 8064 59800 8176 0 FreeSans 448 0 0 0 I[6]
port 12 nsew signal tristate
flabel metal2 s 11424 200 11536 800 0 FreeSans 448 90 0 0 I[7]
port 13 nsew signal tristate
flabel metal3 s 200 39648 800 39760 0 FreeSans 448 0 0 0 I[8]
port 14 nsew signal tristate
flabel metal3 s 200 28224 800 28336 0 FreeSans 448 0 0 0 I[9]
port 15 nsew signal tristate
flabel metal2 s 36960 59200 37072 59800 0 FreeSans 448 90 0 0 Q[0]
port 16 nsew signal tristate
flabel metal2 s 54432 59200 54544 59800 0 FreeSans 448 90 0 0 Q[10]
port 17 nsew signal tristate
flabel metal3 s 200 34272 800 34384 0 FreeSans 448 0 0 0 Q[11]
port 18 nsew signal tristate
flabel metal3 s 59200 48384 59800 48496 0 FreeSans 448 0 0 0 Q[12]
port 19 nsew signal tristate
flabel metal2 s 14112 59200 14224 59800 0 FreeSans 448 90 0 0 Q[1]
port 20 nsew signal tristate
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 Q[2]
port 21 nsew signal tristate
flabel metal3 s 200 11424 800 11536 0 FreeSans 448 0 0 0 Q[3]
port 22 nsew signal tristate
flabel metal3 s 59200 31584 59800 31696 0 FreeSans 448 0 0 0 Q[4]
port 23 nsew signal tristate
flabel metal2 s 8064 59200 8176 59800 0 FreeSans 448 90 0 0 Q[5]
port 24 nsew signal tristate
flabel metal3 s 200 5376 800 5488 0 FreeSans 448 0 0 0 Q[6]
port 25 nsew signal tristate
flabel metal2 s 51744 200 51856 800 0 FreeSans 448 90 0 0 Q[7]
port 26 nsew signal tristate
flabel metal2 s 43008 59200 43120 59800 0 FreeSans 448 90 0 0 Q[8]
port 27 nsew signal tristate
flabel metal3 s 59200 14112 59800 14224 0 FreeSans 448 0 0 0 Q[9]
port 28 nsew signal tristate
flabel metal2 s 5376 200 5488 800 0 FreeSans 448 90 0 0 RST
port 29 nsew signal input
flabel metal2 s 16800 200 16912 800 0 FreeSans 448 90 0 0 addI[0]
port 30 nsew signal tristate
flabel metal2 s 22848 200 22960 800 0 FreeSans 448 90 0 0 addI[1]
port 31 nsew signal tristate
flabel metal3 s 59200 20160 59800 20272 0 FreeSans 448 0 0 0 addI[2]
port 32 nsew signal tristate
flabel metal2 s 28224 200 28336 800 0 FreeSans 448 90 0 0 addI[3]
port 33 nsew signal tristate
flabel metal3 s 59200 54432 59800 54544 0 FreeSans 448 0 0 0 addI[4]
port 34 nsew signal tristate
flabel metal2 s 59808 59200 59920 59800 0 FreeSans 448 90 0 0 addI[5]
port 35 nsew signal tristate
flabel metal2 s 19488 59200 19600 59800 0 FreeSans 448 90 0 0 addQ[0]
port 36 nsew signal tristate
flabel metal2 s 25536 59200 25648 59800 0 FreeSans 448 90 0 0 addQ[1]
port 37 nsew signal tristate
flabel metal2 s 40320 200 40432 800 0 FreeSans 448 90 0 0 addQ[2]
port 38 nsew signal tristate
flabel metal3 s 200 22848 800 22960 0 FreeSans 448 0 0 0 addQ[3]
port 39 nsew signal tristate
flabel metal3 s 200 57120 800 57232 0 FreeSans 448 0 0 0 addQ[4]
port 40 nsew signal tristate
flabel metal3 s 59200 25536 59800 25648 0 FreeSans 448 0 0 0 addQ[5]
port 41 nsew signal tristate
flabel metal4 s 4448 3076 4768 56508 0 FreeSans 1280 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 35168 3076 35488 56508 0 FreeSans 1280 90 0 0 vdd
port 42 nsew power bidirectional
flabel metal4 s 19808 3076 20128 56508 0 FreeSans 1280 90 0 0 vss
port 43 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 56508 0 FreeSans 1280 90 0 0 vss
port 43 nsew ground bidirectional
rlabel metal1 29960 55664 29960 55664 0 vdd
rlabel metal1 29960 56448 29960 56448 0 vss
rlabel metal2 1960 8344 1960 8344 0 BitIn
rlabel metal2 45752 4102 45752 4102 0 CLK
rlabel metal2 31416 55412 31416 55412 0 EN
rlabel metal3 1358 45752 1358 45752 0 I[0]
rlabel metal3 56224 3640 56224 3640 0 I[10]
rlabel metal3 57330 2744 57330 2744 0 I[11]
rlabel metal2 55720 37072 55720 37072 0 I[12]
rlabel metal2 2912 56168 2912 56168 0 I[1]
rlabel metal3 1358 51800 1358 51800 0 I[2]
rlabel metal3 49000 55944 49000 55944 0 I[3]
rlabel metal2 34328 854 34328 854 0 I[4]
rlabel metal2 55384 43232 55384 43232 0 I[5]
rlabel metal2 55384 8232 55384 8232 0 I[6]
rlabel metal2 11480 2058 11480 2058 0 I[7]
rlabel metal3 1358 39704 1358 39704 0 I[8]
rlabel metal3 1358 28280 1358 28280 0 I[9]
rlabel metal2 37912 56280 37912 56280 0 Q[0]
rlabel metal2 54488 57610 54488 57610 0 Q[10]
rlabel metal3 1358 34328 1358 34328 0 Q[11]
rlabel metal3 57666 48440 57666 48440 0 Q[12]
rlabel metal2 15176 56000 15176 56000 0 Q[1]
rlabel metal2 56 1302 56 1302 0 Q[2]
rlabel metal3 1358 11480 1358 11480 0 Q[3]
rlabel metal2 56056 32032 56056 32032 0 Q[4]
rlabel metal2 8120 57610 8120 57610 0 Q[5]
rlabel metal3 1358 5432 1358 5432 0 Q[6]
rlabel metal3 52640 3416 52640 3416 0 Q[7]
rlabel metal2 43624 56504 43624 56504 0 Q[8]
rlabel metal2 55384 14392 55384 14392 0 Q[9]
rlabel metal3 5264 3416 5264 3416 0 RST
rlabel metal2 40936 10192 40936 10192 0 Reg_Delay_Q.In
rlabel metal3 23968 34104 23968 34104 0 Reg_Delay_Q.Out
rlabel metal2 30072 35056 30072 35056 0 _0000_
rlabel metal2 26488 32816 26488 32816 0 _0002_
rlabel metal3 38808 45696 38808 45696 0 _0004_
rlabel metal2 8176 45640 8176 45640 0 _0005_
rlabel metal2 40936 8064 40936 8064 0 _0006_
rlabel metal2 35000 9856 35000 9856 0 _0007_
rlabel metal2 38696 7952 38696 7952 0 _0008_
rlabel metal2 52584 4144 52584 4144 0 _0009_
rlabel metal3 40320 4536 40320 4536 0 _0010_
rlabel metal2 39592 7952 39592 7952 0 _0011_
rlabel metal2 47096 5152 47096 5152 0 _0012_
rlabel metal2 45976 9744 45976 9744 0 _0013_
rlabel metal2 50008 5936 50008 5936 0 _0014_
rlabel metal3 34440 5208 34440 5208 0 _0015_
rlabel metal2 42056 5824 42056 5824 0 _0016_
rlabel metal3 33376 6104 33376 6104 0 _0017_
rlabel metal2 38808 7000 38808 7000 0 _0018_
rlabel metal3 32648 17304 32648 17304 0 _0019_
rlabel metal2 44744 5320 44744 5320 0 _0020_
rlabel metal3 4424 45640 4424 45640 0 _0021_
rlabel metal2 6440 46144 6440 46144 0 _0022_
rlabel metal2 36120 10248 36120 10248 0 _0023_
rlabel metal3 35280 44520 35280 44520 0 _0024_
rlabel metal2 40712 45024 40712 45024 0 _0025_
rlabel metal3 43960 26768 43960 26768 0 _0026_
rlabel metal2 44072 28616 44072 28616 0 _0027_
rlabel metal3 44576 20888 44576 20888 0 _0028_
rlabel metal2 43400 28336 43400 28336 0 _0029_
rlabel metal4 40712 25368 40712 25368 0 _0030_
rlabel metal3 45192 26376 45192 26376 0 _0031_
rlabel metal3 45920 29960 45920 29960 0 _0032_
rlabel metal2 43232 26824 43232 26824 0 _0033_
rlabel metal2 46704 19992 46704 19992 0 _0034_
rlabel metal2 43400 37408 43400 37408 0 _0035_
rlabel metal2 1960 14840 1960 14840 0 _0036_
rlabel metal2 49112 20496 49112 20496 0 _0037_
rlabel metal2 40264 26656 40264 26656 0 _0038_
rlabel metal2 38920 18872 38920 18872 0 _0039_
rlabel metal2 40040 26208 40040 26208 0 _0040_
rlabel metal2 55328 22904 55328 22904 0 _0041_
rlabel metal3 41496 23912 41496 23912 0 _0042_
rlabel metal3 46368 15624 46368 15624 0 _0043_
rlabel metal3 43176 25592 43176 25592 0 _0044_
rlabel metal3 41104 26152 41104 26152 0 _0045_
rlabel metal2 43624 37408 43624 37408 0 _0046_
rlabel metal2 19880 18088 19880 18088 0 _0047_
rlabel metal2 43792 48104 43792 48104 0 _0048_
rlabel metal3 43848 40488 43848 40488 0 _0049_
rlabel metal3 41944 28056 41944 28056 0 _0050_
rlabel metal3 53144 23912 53144 23912 0 _0051_
rlabel metal2 53816 25032 53816 25032 0 _0052_
rlabel metal2 47208 19936 47208 19936 0 _0053_
rlabel metal2 44072 14056 44072 14056 0 _0054_
rlabel metal2 51688 19600 51688 19600 0 _0055_
rlabel metal2 48216 31080 48216 31080 0 _0056_
rlabel metal2 43848 31080 43848 31080 0 _0057_
rlabel metal2 25256 5712 25256 5712 0 _0058_
rlabel metal2 43064 40992 43064 40992 0 _0059_
rlabel metal2 42616 39144 42616 39144 0 _0060_
rlabel metal2 45192 50820 45192 50820 0 _0061_
rlabel metal2 44744 50512 44744 50512 0 _0062_
rlabel metal2 43400 50792 43400 50792 0 _0063_
rlabel metal2 42504 50792 42504 50792 0 _0064_
rlabel metal2 48048 21672 48048 21672 0 _0065_
rlabel metal3 47432 32536 47432 32536 0 _0066_
rlabel metal2 47544 22064 47544 22064 0 _0067_
rlabel metal2 46984 23576 46984 23576 0 _0068_
rlabel metal2 24920 7000 24920 7000 0 _0069_
rlabel metal2 48496 23688 48496 23688 0 _0070_
rlabel metal2 47264 24024 47264 24024 0 _0071_
rlabel metal2 50456 25788 50456 25788 0 _0072_
rlabel metal2 49672 24920 49672 24920 0 _0073_
rlabel metal3 49448 2800 49448 2800 0 _0074_
rlabel metal2 50064 23912 50064 23912 0 _0075_
rlabel metal2 47992 24416 47992 24416 0 _0076_
rlabel metal2 47208 28672 47208 28672 0 _0077_
rlabel metal3 29848 28504 29848 28504 0 _0078_
rlabel metal2 33096 28784 33096 28784 0 _0079_
rlabel metal2 21784 9520 21784 9520 0 _0080_
rlabel metal2 43960 53368 43960 53368 0 _0081_
rlabel metal3 38920 54376 38920 54376 0 _0082_
rlabel metal2 39760 55272 39760 55272 0 _0083_
rlabel metal3 44744 50568 44744 50568 0 _0084_
rlabel metal2 43960 54096 43960 54096 0 _0085_
rlabel metal3 53088 47320 53088 47320 0 _0086_
rlabel metal2 40264 44464 40264 44464 0 _0087_
rlabel metal2 49784 50904 49784 50904 0 _0088_
rlabel metal2 48552 24584 48552 24584 0 _0089_
rlabel metal3 43344 22904 43344 22904 0 _0090_
rlabel metal3 18760 7448 18760 7448 0 _0091_
rlabel metal3 49168 25256 49168 25256 0 _0092_
rlabel metal2 50848 25368 50848 25368 0 _0093_
rlabel metal2 42504 18648 42504 18648 0 _0094_
rlabel metal3 47768 2968 47768 2968 0 _0095_
rlabel metal3 54880 24920 54880 24920 0 _0096_
rlabel metal2 54152 22456 54152 22456 0 _0097_
rlabel metal3 52360 25480 52360 25480 0 _0098_
rlabel metal2 50456 50960 50456 50960 0 _0099_
rlabel metal2 50288 50792 50288 50792 0 _0100_
rlabel metal3 48496 52024 48496 52024 0 _0101_
rlabel metal2 23800 9128 23800 9128 0 _0102_
rlabel metal2 47656 51856 47656 51856 0 _0103_
rlabel metal3 44016 28616 44016 28616 0 _0104_
rlabel metal2 47432 25144 47432 25144 0 _0105_
rlabel metal2 51800 21392 51800 21392 0 _0106_
rlabel metal3 51296 30744 51296 30744 0 _0107_
rlabel metal3 48104 2632 48104 2632 0 _0108_
rlabel metal3 42672 18424 42672 18424 0 _0109_
rlabel metal2 48552 18928 48552 18928 0 _0110_
rlabel metal2 46424 19040 46424 19040 0 _0111_
rlabel metal3 53704 30408 53704 30408 0 _0112_
rlabel metal2 15288 6328 15288 6328 0 _0113_
rlabel metal3 53760 19432 53760 19432 0 _0114_
rlabel metal2 54264 32032 54264 32032 0 _0115_
rlabel metal2 53760 30968 53760 30968 0 _0116_
rlabel metal2 49784 47152 49784 47152 0 _0117_
rlabel metal2 46984 45696 46984 45696 0 _0118_
rlabel metal2 41048 39368 41048 39368 0 _0119_
rlabel metal2 50232 40880 50232 40880 0 _0120_
rlabel metal2 48104 51240 48104 51240 0 _0121_
rlabel metal2 47320 51408 47320 51408 0 _0122_
rlabel metal2 47544 51576 47544 51576 0 _0123_
rlabel metal2 19656 5712 19656 5712 0 _0124_
rlabel metal3 45640 52248 45640 52248 0 _0125_
rlabel metal2 44408 53032 44408 53032 0 _0126_
rlabel metal2 34216 29008 34216 29008 0 _0127_
rlabel metal2 33992 34384 33992 34384 0 _0128_
rlabel metal2 48552 30016 48552 30016 0 _0129_
rlabel metal2 47432 30464 47432 30464 0 _0130_
rlabel metal4 40376 19432 40376 19432 0 _0131_
rlabel metal2 49448 29512 49448 29512 0 _0132_
rlabel metal2 46144 26152 46144 26152 0 _0133_
rlabel metal3 48160 28840 48160 28840 0 _0134_
rlabel metal2 19320 8288 19320 8288 0 _0135_
rlabel metal3 39704 30352 39704 30352 0 _0136_
rlabel metal3 44912 53480 44912 53480 0 _0137_
rlabel metal2 43848 54432 43848 54432 0 _0138_
rlabel metal2 43736 53200 43736 53200 0 _0139_
rlabel metal3 42056 54488 42056 54488 0 _0140_
rlabel metal3 41384 54376 41384 54376 0 _0141_
rlabel metal2 40600 54992 40600 54992 0 _0142_
rlabel metal3 2968 53592 2968 53592 0 _0143_
rlabel metal2 36120 51968 36120 51968 0 _0144_
rlabel metal3 19768 10584 19768 10584 0 _0145_
rlabel metal2 43064 52696 43064 52696 0 _0146_
rlabel metal2 42056 54152 42056 54152 0 _0147_
rlabel metal2 40040 44800 40040 44800 0 _0148_
rlabel metal2 49616 13048 49616 13048 0 _0149_
rlabel metal2 50232 14448 50232 14448 0 _0150_
rlabel metal3 50960 15176 50960 15176 0 _0151_
rlabel metal3 47320 24920 47320 24920 0 _0152_
rlabel metal2 47824 21000 47824 21000 0 _0153_
rlabel metal2 38808 26236 38808 26236 0 _0154_
rlabel metal3 45360 27832 45360 27832 0 _0155_
rlabel metal2 23352 9576 23352 9576 0 _0156_
rlabel metal2 47544 34832 47544 34832 0 _0157_
rlabel metal3 52472 27272 52472 27272 0 _0158_
rlabel metal2 52472 25032 52472 25032 0 _0159_
rlabel metal3 47712 1624 47712 1624 0 _0160_
rlabel metal2 54600 26712 54600 26712 0 _0161_
rlabel metal2 52136 44632 52136 44632 0 _0162_
rlabel metal2 51576 42392 51576 42392 0 _0163_
rlabel metal2 53816 46984 53816 46984 0 _0164_
rlabel metal3 40712 46928 40712 46928 0 _0165_
rlabel metal2 45640 45360 45640 45360 0 _0166_
rlabel metal2 22456 21728 22456 21728 0 _0167_
rlabel metal2 45136 43624 45136 43624 0 _0168_
rlabel metal2 47880 45024 47880 45024 0 _0169_
rlabel metal2 53704 31920 53704 31920 0 _0170_
rlabel metal2 56448 29624 56448 29624 0 _0171_
rlabel metal3 54320 46872 54320 46872 0 _0172_
rlabel metal2 49560 49504 49560 49504 0 _0173_
rlabel metal2 52248 28168 52248 28168 0 _0174_
rlabel metal2 52584 26768 52584 26768 0 _0175_
rlabel metal2 50008 28952 50008 28952 0 _0176_
rlabel metal3 51352 28392 51352 28392 0 _0177_
rlabel metal2 23352 26992 23352 26992 0 _0178_
rlabel metal2 54096 48440 54096 48440 0 _0179_
rlabel metal2 49672 43456 49672 43456 0 _0180_
rlabel metal2 46256 44520 46256 44520 0 _0181_
rlabel metal2 46200 43736 46200 43736 0 _0182_
rlabel metal2 44184 47880 44184 47880 0 _0183_
rlabel via2 47432 40936 47432 40936 0 _0184_
rlabel metal2 47544 45584 47544 45584 0 _0185_
rlabel metal2 44632 48048 44632 48048 0 _0186_
rlabel metal2 40488 48496 40488 48496 0 _0187_
rlabel metal3 40488 49000 40488 49000 0 _0188_
rlabel metal2 28616 26208 28616 26208 0 _0189_
rlabel metal2 40152 22792 40152 22792 0 _0190_
rlabel metal2 40040 21784 40040 21784 0 _0191_
rlabel metal3 44296 23240 44296 23240 0 _0192_
rlabel metal2 40096 23352 40096 23352 0 _0193_
rlabel metal2 41048 25312 41048 25312 0 _0194_
rlabel metal2 41944 24528 41944 24528 0 _0195_
rlabel metal2 39928 24976 39928 24976 0 _0196_
rlabel metal2 39536 24920 39536 24920 0 _0197_
rlabel metal3 32928 33320 32928 33320 0 _0198_
rlabel metal3 39144 49672 39144 49672 0 _0199_
rlabel metal2 23576 28672 23576 28672 0 _0200_
rlabel metal2 40768 53032 40768 53032 0 _0201_
rlabel metal2 40488 52920 40488 52920 0 _0202_
rlabel metal2 42616 54152 42616 54152 0 _0203_
rlabel metal3 42448 55272 42448 55272 0 _0204_
rlabel metal3 45416 55160 45416 55160 0 _0205_
rlabel metal2 40376 45920 40376 45920 0 _0206_
rlabel metal2 40600 50568 40600 50568 0 _0207_
rlabel metal3 38808 51352 38808 51352 0 _0208_
rlabel metal2 51352 45752 51352 45752 0 _0209_
rlabel metal2 23800 16352 23800 16352 0 _0210_
rlabel metal2 45976 46032 45976 46032 0 _0211_
rlabel metal2 49896 33768 49896 33768 0 _0212_
rlabel metal3 46816 34216 46816 34216 0 _0213_
rlabel metal2 49784 35000 49784 35000 0 _0214_
rlabel metal3 51072 35784 51072 35784 0 _0215_
rlabel metal2 50512 33096 50512 33096 0 _0216_
rlabel metal3 48496 22232 48496 22232 0 _0217_
rlabel metal4 50232 30016 50232 30016 0 _0218_
rlabel metal2 50120 32928 50120 32928 0 _0219_
rlabel metal2 50680 35504 50680 35504 0 _0220_
rlabel metal3 24976 26824 24976 26824 0 _0221_
rlabel metal3 44632 46648 44632 46648 0 _0222_
rlabel metal2 42952 47096 42952 47096 0 _0223_
rlabel metal3 43568 42728 43568 42728 0 _0224_
rlabel metal2 47432 19656 47432 19656 0 _0225_
rlabel metal3 48832 34776 48832 34776 0 _0226_
rlabel metal2 49112 32200 49112 32200 0 _0227_
rlabel metal2 47152 32312 47152 32312 0 _0228_
rlabel metal2 48216 35280 48216 35280 0 _0229_
rlabel metal2 40600 33488 40600 33488 0 _0230_
rlabel metal2 48776 35280 48776 35280 0 _0231_
rlabel metal3 5600 9800 5600 9800 0 _0232_
rlabel metal2 48328 36624 48328 36624 0 _0233_
rlabel metal2 48104 34216 48104 34216 0 _0234_
rlabel metal2 46424 39984 46424 39984 0 _0235_
rlabel metal2 46872 40488 46872 40488 0 _0236_
rlabel metal3 44016 40936 44016 40936 0 _0237_
rlabel metal2 42504 43456 42504 43456 0 _0238_
rlabel metal2 43288 46704 43288 46704 0 _0239_
rlabel metal3 42392 36344 42392 36344 0 _0240_
rlabel metal2 41608 16184 41608 16184 0 _0241_
rlabel metal3 43680 19432 43680 19432 0 _0242_
rlabel metal2 2856 9296 2856 9296 0 _0243_
rlabel metal2 45416 34440 45416 34440 0 _0244_
rlabel metal3 42728 39368 42728 39368 0 _0245_
rlabel metal2 44632 30520 44632 30520 0 _0246_
rlabel metal3 45192 31192 45192 31192 0 _0247_
rlabel metal2 41832 18256 41832 18256 0 _0248_
rlabel metal2 45752 27888 45752 27888 0 _0249_
rlabel metal2 44688 31976 44688 31976 0 _0250_
rlabel metal3 45584 36456 45584 36456 0 _0251_
rlabel metal2 44240 37464 44240 37464 0 _0252_
rlabel metal2 42952 41608 42952 41608 0 _0253_
rlabel metal2 19208 8960 19208 8960 0 _0254_
rlabel metal2 48216 42672 48216 42672 0 _0255_
rlabel metal2 45920 35896 45920 35896 0 _0256_
rlabel metal2 44856 43344 44856 43344 0 _0257_
rlabel metal2 43064 43064 43064 43064 0 _0258_
rlabel metal2 43568 46648 43568 46648 0 _0259_
rlabel metal2 36624 50568 36624 50568 0 _0260_
rlabel metal2 47656 43848 47656 43848 0 _0261_
rlabel metal2 49672 35728 49672 35728 0 _0262_
rlabel metal2 47376 50792 47376 50792 0 _0263_
rlabel metal3 48048 44296 48048 44296 0 _0264_
rlabel metal3 19824 9240 19824 9240 0 _0265_
rlabel metal2 43848 44296 43848 44296 0 _0266_
rlabel metal2 42392 43960 42392 43960 0 _0267_
rlabel metal2 42728 44800 42728 44800 0 _0268_
rlabel metal2 43960 45416 43960 45416 0 _0269_
rlabel metal3 41328 52248 41328 52248 0 _0270_
rlabel metal3 37968 51576 37968 51576 0 _0271_
rlabel metal2 39816 23632 39816 23632 0 _0272_
rlabel metal2 39760 23912 39760 23912 0 _0273_
rlabel metal3 35392 19096 35392 19096 0 _0274_
rlabel metal2 35896 18704 35896 18704 0 _0275_
rlabel metal2 16296 9856 16296 9856 0 _0276_
rlabel metal2 37464 19208 37464 19208 0 _0277_
rlabel metal2 42392 15512 42392 15512 0 _0278_
rlabel metal2 37688 19936 37688 19936 0 _0279_
rlabel metal2 37128 18760 37128 18760 0 _0280_
rlabel metal2 40152 16772 40152 16772 0 _0281_
rlabel metal3 36680 18536 36680 18536 0 _0282_
rlabel metal2 35672 19208 35672 19208 0 _0283_
rlabel metal2 33992 31472 33992 31472 0 _0284_
rlabel metal3 35560 50456 35560 50456 0 _0285_
rlabel metal3 34776 51352 34776 51352 0 _0286_
rlabel metal2 18760 7168 18760 7168 0 _0287_
rlabel metal3 39200 52808 39200 52808 0 _0288_
rlabel metal3 39872 53704 39872 53704 0 _0289_
rlabel metal2 41720 53200 41720 53200 0 _0290_
rlabel metal2 41608 53760 41608 53760 0 _0291_
rlabel metal2 36008 53368 36008 53368 0 _0292_
rlabel metal2 33712 51352 33712 51352 0 _0293_
rlabel metal3 31864 51240 31864 51240 0 _0294_
rlabel metal2 42728 47264 42728 47264 0 _0295_
rlabel metal2 33768 49504 33768 49504 0 _0296_
rlabel metal2 2184 20160 2184 20160 0 _0297_
rlabel metal2 39088 22456 39088 22456 0 _0298_
rlabel metal2 46648 29456 46648 29456 0 _0299_
rlabel metal2 40264 31976 40264 31976 0 _0300_
rlabel metal2 42168 34608 42168 34608 0 _0301_
rlabel metal2 40600 31864 40600 31864 0 _0302_
rlabel metal2 38920 25872 38920 25872 0 _0303_
rlabel metal3 39032 23688 39032 23688 0 _0304_
rlabel metal3 39256 35672 39256 35672 0 _0305_
rlabel metal2 40712 35112 40712 35112 0 _0306_
rlabel metal2 40656 21000 40656 21000 0 _0307_
rlabel metal2 25760 10024 25760 10024 0 _0308_
rlabel metal2 40600 34608 40600 34608 0 _0309_
rlabel metal2 50904 51464 50904 51464 0 _0310_
rlabel metal2 53984 41832 53984 41832 0 _0311_
rlabel metal2 54320 44520 54320 44520 0 _0312_
rlabel metal2 50008 46648 50008 46648 0 _0313_
rlabel metal2 49672 47768 49672 47768 0 _0314_
rlabel metal2 46872 46256 46872 46256 0 _0315_
rlabel metal2 46648 47432 46648 47432 0 _0316_
rlabel metal2 46088 47376 46088 47376 0 _0317_
rlabel metal3 48720 49000 48720 49000 0 _0318_
rlabel metal2 16856 4816 16856 4816 0 _0319_
rlabel metal2 48776 50820 48776 50820 0 _0320_
rlabel metal3 48104 51800 48104 51800 0 _0321_
rlabel metal3 47376 49112 47376 49112 0 _0322_
rlabel metal2 46424 51240 46424 51240 0 _0323_
rlabel metal2 35168 47544 35168 47544 0 _0324_
rlabel metal2 30296 49392 30296 49392 0 _0325_
rlabel metal2 36904 28560 36904 28560 0 _0326_
rlabel metal2 36512 35448 36512 35448 0 _0327_
rlabel metal2 39032 29568 39032 29568 0 _0328_
rlabel metal2 36792 28616 36792 28616 0 _0329_
rlabel metal3 21448 18200 21448 18200 0 _0330_
rlabel metal2 36400 28616 36400 28616 0 _0331_
rlabel metal2 31752 29232 31752 29232 0 _0332_
rlabel metal2 31864 30016 31864 30016 0 _0333_
rlabel metal3 30856 30408 30856 30408 0 _0334_
rlabel metal2 30520 45360 30520 45360 0 _0335_
rlabel metal2 32480 51352 32480 51352 0 _0336_
rlabel metal2 35616 50344 35616 50344 0 _0337_
rlabel metal2 36232 51212 36232 51212 0 _0338_
rlabel metal2 34160 52360 34160 52360 0 _0339_
rlabel metal3 33040 52808 33040 52808 0 _0340_
rlabel metal2 23800 22288 23800 22288 0 _0341_
rlabel metal2 32760 50960 32760 50960 0 _0342_
rlabel metal2 31472 48440 31472 48440 0 _0343_
rlabel metal2 30296 47712 30296 47712 0 _0344_
rlabel metal3 40152 42504 40152 42504 0 _0345_
rlabel metal2 50344 39648 50344 39648 0 _0346_
rlabel metal2 43736 43232 43736 43232 0 _0347_
rlabel metal2 32088 22064 32088 22064 0 _0348_
rlabel metal2 39032 39032 39032 39032 0 _0349_
rlabel metal2 36400 25480 36400 25480 0 _0350_
rlabel metal2 19320 4816 19320 4816 0 _0351_
rlabel metal2 38696 26320 38696 26320 0 _0352_
rlabel metal2 39424 20552 39424 20552 0 _0353_
rlabel metal2 37688 24360 37688 24360 0 _0354_
rlabel metal2 39256 26096 39256 26096 0 _0355_
rlabel metal2 37464 25144 37464 25144 0 _0356_
rlabel metal2 40040 39872 40040 39872 0 _0357_
rlabel metal3 39592 42728 39592 42728 0 _0358_
rlabel metal3 40096 42168 40096 42168 0 _0359_
rlabel metal3 39928 41048 39928 41048 0 _0360_
rlabel metal2 38920 41552 38920 41552 0 _0361_
rlabel metal2 10808 15736 10808 15736 0 _0362_
rlabel metal3 45976 42840 45976 42840 0 _0363_
rlabel metal2 39144 41608 39144 41608 0 _0364_
rlabel metal3 41664 15288 41664 15288 0 _0365_
rlabel metal2 41328 17416 41328 17416 0 _0366_
rlabel metal2 42224 17752 42224 17752 0 _0367_
rlabel metal2 42560 17864 42560 17864 0 _0368_
rlabel metal2 41048 18032 41048 18032 0 _0369_
rlabel metal2 45528 38668 45528 38668 0 _0370_
rlabel metal3 43344 15288 43344 15288 0 _0371_
rlabel metal3 43512 15176 43512 15176 0 _0372_
rlabel metal2 22400 5096 22400 5096 0 _0373_
rlabel metal2 46592 38920 46592 38920 0 _0374_
rlabel metal2 46088 43288 46088 43288 0 _0375_
rlabel metal2 46368 42952 46368 42952 0 _0376_
rlabel metal2 46088 39088 46088 39088 0 _0377_
rlabel metal2 46312 41720 46312 41720 0 _0378_
rlabel metal3 42728 42616 42728 42616 0 _0379_
rlabel metal2 39200 44072 39200 44072 0 _0380_
rlabel metal2 40208 42168 40208 42168 0 _0381_
rlabel metal2 40040 43176 40040 43176 0 _0382_
rlabel metal3 43176 41944 43176 41944 0 _0383_
rlabel metal2 1960 13104 1960 13104 0 _0384_
rlabel metal2 39368 43792 39368 43792 0 _0385_
rlabel metal2 38808 44016 38808 44016 0 _0386_
rlabel metal2 30968 24360 30968 24360 0 _0387_
rlabel metal2 34776 22848 34776 22848 0 _0388_
rlabel metal2 37800 21168 37800 21168 0 _0389_
rlabel metal3 37072 22344 37072 22344 0 _0390_
rlabel metal2 35112 22848 35112 22848 0 _0391_
rlabel metal2 32312 22680 32312 22680 0 _0392_
rlabel metal2 33768 17976 33768 17976 0 _0393_
rlabel metal2 31976 22512 31976 22512 0 _0394_
rlabel metal2 23464 5544 23464 5544 0 _0395_
rlabel metal2 31864 23632 31864 23632 0 _0396_
rlabel metal3 30856 45080 30856 45080 0 _0397_
rlabel metal2 29960 46928 29960 46928 0 _0398_
rlabel metal3 31808 47320 31808 47320 0 _0399_
rlabel metal3 33488 49224 33488 49224 0 _0400_
rlabel metal2 34048 47992 34048 47992 0 _0401_
rlabel metal2 32872 48552 32872 48552 0 _0402_
rlabel metal2 33320 49392 33320 49392 0 _0403_
rlabel metal2 34552 48720 34552 48720 0 _0404_
rlabel metal2 33768 47656 33768 47656 0 _0405_
rlabel metal2 10360 8680 10360 8680 0 _0406_
rlabel metal3 34608 48776 34608 48776 0 _0407_
rlabel metal2 31192 47824 31192 47824 0 _0408_
rlabel metal2 29848 46088 29848 46088 0 _0409_
rlabel metal2 39144 8120 39144 8120 0 _0410_
rlabel metal2 31528 44128 31528 44128 0 _0411_
rlabel metal2 40152 39256 40152 39256 0 _0412_
rlabel metal2 40712 27944 40712 27944 0 _0413_
rlabel metal2 44744 28112 44744 28112 0 _0414_
rlabel metal2 42728 19712 42728 19712 0 _0415_
rlabel metal2 10920 10920 10920 10920 0 _0416_
rlabel metal2 42728 27104 42728 27104 0 _0417_
rlabel metal3 43008 26376 43008 26376 0 _0418_
rlabel metal3 43512 26824 43512 26824 0 _0419_
rlabel metal2 42840 28336 42840 28336 0 _0420_
rlabel metal2 41608 39928 41608 39928 0 _0421_
rlabel metal2 42168 41496 42168 41496 0 _0422_
rlabel metal2 41720 41216 41720 41216 0 _0423_
rlabel metal2 31864 42000 31864 42000 0 _0424_
rlabel metal3 37464 41944 37464 41944 0 _0425_
rlabel metal2 37912 31304 37912 31304 0 _0426_
rlabel metal2 29512 16296 29512 16296 0 _0427_
rlabel metal3 36624 31752 36624 31752 0 _0428_
rlabel metal2 38136 30800 38136 30800 0 _0429_
rlabel metal3 37016 31528 37016 31528 0 _0430_
rlabel metal2 36792 40600 36792 40600 0 _0431_
rlabel metal2 37352 42280 37352 42280 0 _0432_
rlabel metal2 31640 42000 31640 42000 0 _0433_
rlabel metal3 32144 42728 32144 42728 0 _0434_
rlabel metal3 33656 24920 33656 24920 0 _0435_
rlabel metal3 33936 23800 33936 23800 0 _0436_
rlabel metal3 32872 23352 32872 23352 0 _0437_
rlabel metal2 2632 15568 2632 15568 0 _0438_
rlabel metal2 34888 18088 34888 18088 0 _0439_
rlabel metal2 33040 23128 33040 23128 0 _0440_
rlabel metal2 32312 23632 32312 23632 0 _0441_
rlabel metal3 30520 24136 30520 24136 0 _0442_
rlabel metal2 31136 42952 31136 42952 0 _0443_
rlabel metal3 31472 42616 31472 42616 0 _0444_
rlabel metal2 29904 44296 29904 44296 0 _0445_
rlabel metal2 31192 44464 31192 44464 0 _0446_
rlabel metal2 29624 43848 29624 43848 0 _0447_
rlabel metal3 29624 45304 29624 45304 0 _0448_
rlabel metal3 22008 29288 22008 29288 0 _0449_
rlabel metal2 28392 44912 28392 44912 0 _0450_
rlabel metal3 30520 25256 30520 25256 0 _0451_
rlabel metal3 30744 41048 30744 41048 0 _0452_
rlabel metal2 28952 40656 28952 40656 0 _0453_
rlabel metal2 39928 23464 39928 23464 0 _0454_
rlabel metal3 36792 21000 36792 21000 0 _0455_
rlabel metal2 36568 22736 36568 22736 0 _0456_
rlabel metal2 41608 23072 41608 23072 0 _0457_
rlabel metal3 35448 26768 35448 26768 0 _0458_
rlabel metal3 23464 29288 23464 29288 0 _0459_
rlabel metal2 35728 39816 35728 39816 0 _0460_
rlabel metal2 36344 40880 36344 40880 0 _0461_
rlabel metal2 50232 42000 50232 42000 0 _0462_
rlabel metal2 33656 39984 33656 39984 0 _0463_
rlabel metal2 39368 29680 39368 29680 0 _0464_
rlabel metal2 38024 39592 38024 39592 0 _0465_
rlabel metal3 38080 38024 38080 38024 0 _0466_
rlabel metal2 34216 38752 34216 38752 0 _0467_
rlabel metal3 36064 40488 36064 40488 0 _0468_
rlabel metal2 33544 40040 33544 40040 0 _0469_
rlabel metal2 2408 7952 2408 7952 0 _0470_
rlabel metal3 32256 39480 32256 39480 0 _0471_
rlabel metal3 31808 26264 31808 26264 0 _0472_
rlabel metal3 31864 26152 31864 26152 0 _0473_
rlabel metal3 34216 21560 34216 21560 0 _0474_
rlabel metal2 39032 34608 39032 34608 0 _0475_
rlabel metal3 33264 25368 33264 25368 0 _0476_
rlabel metal2 31472 28504 31472 28504 0 _0477_
rlabel metal3 30520 28840 30520 28840 0 _0478_
rlabel metal3 29624 29960 29624 29960 0 _0479_
rlabel metal2 38920 33264 38920 33264 0 _0480_
rlabel metal2 21560 14000 21560 14000 0 _0481_
rlabel metal3 30016 29624 30016 29624 0 _0482_
rlabel metal3 30240 30072 30240 30072 0 _0483_
rlabel metal2 30632 39312 30632 39312 0 _0484_
rlabel metal3 29848 40376 29848 40376 0 _0485_
rlabel metal3 27944 40376 27944 40376 0 _0486_
rlabel metal2 28504 44632 28504 44632 0 _0487_
rlabel metal2 31080 45024 31080 45024 0 _0488_
rlabel metal3 28392 40264 28392 40264 0 _0489_
rlabel metal2 3192 40152 3192 40152 0 _0490_
rlabel metal2 24024 10360 24024 10360 0 _0491_
rlabel metal3 32984 39032 32984 39032 0 _0492_
rlabel metal2 30856 37520 30856 37520 0 _0493_
rlabel metal2 43960 26152 43960 26152 0 _0494_
rlabel metal2 36904 32872 36904 32872 0 _0495_
rlabel metal3 35448 33544 35448 33544 0 _0496_
rlabel metal2 34776 40768 34776 40768 0 _0497_
rlabel metal2 34328 41440 34328 41440 0 _0498_
rlabel metal3 34720 41048 34720 41048 0 _0499_
rlabel metal2 33936 39816 33936 39816 0 _0500_
rlabel metal2 36008 36456 36008 36456 0 _0501_
rlabel metal2 23464 13944 23464 13944 0 _0502_
rlabel metal2 36456 24528 36456 24528 0 _0503_
rlabel metal2 38808 37072 38808 37072 0 _0504_
rlabel metal2 36904 37632 36904 37632 0 _0505_
rlabel metal2 35336 37688 35336 37688 0 _0506_
rlabel metal2 34104 38080 34104 38080 0 _0507_
rlabel metal2 32760 37296 32760 37296 0 _0508_
rlabel metal2 31024 25368 31024 25368 0 _0509_
rlabel metal2 31304 25592 31304 25592 0 _0510_
rlabel metal2 30576 27048 30576 27048 0 _0511_
rlabel metal2 31192 36344 31192 36344 0 _0512_
rlabel metal3 22792 28728 22792 28728 0 _0513_
rlabel metal3 30296 37128 30296 37128 0 _0514_
rlabel metal3 28616 38024 28616 38024 0 _0515_
rlabel metal2 29904 39816 29904 39816 0 _0516_
rlabel metal3 28840 39368 28840 39368 0 _0517_
rlabel metal2 27496 37520 27496 37520 0 _0518_
rlabel metal2 27160 37184 27160 37184 0 _0519_
rlabel metal3 55608 38808 55608 38808 0 _0520_
rlabel metal3 37800 35672 37800 35672 0 _0521_
rlabel metal3 24024 29400 24024 29400 0 _0522_
rlabel metal2 44408 37744 44408 37744 0 _0523_
rlabel metal2 54208 42616 54208 42616 0 _0524_
rlabel metal2 54040 43624 54040 43624 0 _0525_
rlabel metal2 36064 38024 36064 38024 0 _0526_
rlabel metal3 36512 38248 36512 38248 0 _0527_
rlabel metal3 37632 39704 37632 39704 0 _0528_
rlabel metal2 39368 39816 39368 39816 0 _0529_
rlabel metal2 55104 42728 55104 42728 0 _0530_
rlabel metal3 41720 55496 41720 55496 0 _0531_
rlabel metal3 55384 40936 55384 40936 0 _0532_
rlabel metal3 24360 31752 24360 31752 0 _0533_
rlabel metal2 56056 39368 56056 39368 0 _0534_
rlabel metal3 33264 37464 33264 37464 0 _0535_
rlabel metal3 55608 46536 55608 46536 0 _0536_
rlabel metal2 56168 37408 56168 37408 0 _0537_
rlabel metal3 57008 35672 57008 35672 0 _0538_
rlabel metal3 30464 38024 30464 38024 0 _0539_
rlabel metal3 30632 37800 30632 37800 0 _0540_
rlabel metal3 30240 38808 30240 38808 0 _0541_
rlabel metal2 49560 38808 49560 38808 0 _0542_
rlabel metal4 49448 2744 49448 2744 0 _0543_
rlabel metal2 22008 32256 22008 32256 0 _0544_
rlabel metal2 54544 42728 54544 42728 0 _0545_
rlabel metal2 56168 40768 56168 40768 0 _0546_
rlabel metal3 48496 40600 48496 40600 0 _0547_
rlabel metal2 48496 39032 48496 39032 0 _0548_
rlabel metal2 48664 40824 48664 40824 0 _0549_
rlabel metal2 49336 41608 49336 41608 0 _0550_
rlabel metal3 53200 41944 53200 41944 0 _0551_
rlabel metal3 55440 40376 55440 40376 0 _0552_
rlabel metal2 56840 40264 56840 40264 0 _0553_
rlabel metal2 23912 33880 23912 33880 0 _0554_
rlabel metal2 56616 39312 56616 39312 0 _0555_
rlabel metal2 57792 35896 57792 35896 0 _0556_
rlabel metal3 58016 3304 58016 3304 0 _0557_
rlabel metal3 56280 38024 56280 38024 0 _0558_
rlabel metal2 57288 38920 57288 38920 0 _0559_
rlabel metal2 55720 40040 55720 40040 0 _0560_
rlabel metal3 56224 39032 56224 39032 0 _0561_
rlabel metal3 55384 39480 55384 39480 0 _0562_
rlabel metal2 57064 39536 57064 39536 0 _0563_
rlabel metal3 55888 42056 55888 42056 0 _0564_
rlabel metal2 56616 41552 56616 41552 0 _0565_
rlabel metal2 56840 39928 56840 39928 0 _0566_
rlabel metal2 37632 54600 37632 54600 0 _0567_
rlabel metal2 39928 13328 39928 13328 0 _0568_
rlabel metal2 34776 11256 34776 11256 0 _0569_
rlabel metal3 47320 41048 47320 41048 0 _0570_
rlabel metal2 33544 18704 33544 18704 0 _0571_
rlabel metal2 32760 17528 32760 17528 0 _0572_
rlabel metal2 34104 12152 34104 12152 0 _0573_
rlabel metal3 41384 12824 41384 12824 0 _0574_
rlabel metal2 42952 12824 42952 12824 0 _0575_
rlabel metal2 39368 14224 39368 14224 0 _0576_
rlabel metal2 40880 13160 40880 13160 0 _0577_
rlabel metal2 47544 40544 47544 40544 0 _0578_
rlabel metal3 37184 15960 37184 15960 0 _0579_
rlabel metal3 36904 15288 36904 15288 0 _0580_
rlabel metal2 37016 15792 37016 15792 0 _0581_
rlabel metal2 37800 13272 37800 13272 0 _0582_
rlabel metal2 36176 14728 36176 14728 0 _0583_
rlabel metal2 33544 16408 33544 16408 0 _0584_
rlabel metal2 36344 17360 36344 17360 0 _0585_
rlabel metal3 43064 39480 43064 39480 0 _0586_
rlabel metal2 33768 16296 33768 16296 0 _0587_
rlabel metal2 35560 18144 35560 18144 0 _0588_
rlabel metal2 35560 16464 35560 16464 0 _0589_
rlabel metal3 29792 14504 29792 14504 0 _0590_
rlabel metal3 33264 15288 33264 15288 0 _0591_
rlabel metal2 40376 39004 40376 39004 0 _0592_
rlabel metal3 31752 17080 31752 17080 0 _0593_
rlabel metal2 31192 18480 31192 18480 0 _0594_
rlabel metal2 32648 18536 32648 18536 0 _0595_
rlabel metal2 5992 45136 5992 45136 0 _0596_
rlabel metal3 35616 12264 35616 12264 0 _0597_
rlabel metal2 35896 11256 35896 11256 0 _0598_
rlabel metal3 32032 23576 32032 23576 0 _0599_
rlabel metal2 36512 44296 36512 44296 0 _0600_
rlabel metal2 31080 29008 31080 29008 0 _0601_
rlabel metal2 31416 31304 31416 31304 0 _0602_
rlabel metal2 38920 13104 38920 13104 0 _0603_
rlabel metal3 30240 33432 30240 33432 0 _0604_
rlabel metal2 32368 35112 32368 35112 0 _0605_
rlabel metal3 30520 34104 30520 34104 0 _0606_
rlabel metal2 29848 35000 29848 35000 0 _0607_
rlabel metal2 16968 36064 16968 36064 0 _0608_
rlabel metal2 16072 39088 16072 39088 0 _0609_
rlabel metal3 22176 32536 22176 32536 0 _0610_
rlabel metal3 17192 33096 17192 33096 0 _0611_
rlabel metal2 26152 25676 26152 25676 0 _0612_
rlabel metal2 24248 32592 24248 32592 0 _0613_
rlabel metal3 26488 32536 26488 32536 0 _0614_
rlabel metal2 25872 32760 25872 32760 0 _0615_
rlabel metal3 30576 33096 30576 33096 0 _0616_
rlabel metal2 27944 33824 27944 33824 0 _0617_
rlabel metal2 15512 25200 15512 25200 0 _0618_
rlabel metal3 12656 27832 12656 27832 0 _0619_
rlabel metal3 22288 8008 22288 8008 0 _0620_
rlabel metal2 7560 16184 7560 16184 0 _0621_
rlabel metal2 19880 21784 19880 21784 0 _0622_
rlabel metal3 13328 6664 13328 6664 0 _0623_
rlabel metal2 12264 8008 12264 8008 0 _0624_
rlabel metal3 4312 18424 4312 18424 0 _0625_
rlabel metal2 15064 7280 15064 7280 0 _0626_
rlabel metal2 16184 3920 16184 3920 0 _0627_
rlabel metal2 6888 17864 6888 17864 0 _0628_
rlabel metal2 7392 19992 7392 19992 0 _0629_
rlabel metal2 18088 9408 18088 9408 0 _0630_
rlabel metal2 4200 6944 4200 6944 0 _0631_
rlabel metal2 26488 8568 26488 8568 0 _0632_
rlabel metal3 2856 14448 2856 14448 0 _0633_
rlabel metal2 18984 6496 18984 6496 0 _0634_
rlabel metal2 2184 17808 2184 17808 0 _0635_
rlabel metal3 8176 21784 8176 21784 0 _0636_
rlabel metal2 16856 11760 16856 11760 0 _0637_
rlabel metal2 22344 20384 22344 20384 0 _0638_
rlabel metal2 18984 11424 18984 11424 0 _0639_
rlabel metal2 2296 27328 2296 27328 0 _0640_
rlabel metal3 16632 28056 16632 28056 0 _0641_
rlabel metal2 15736 28168 15736 28168 0 _0642_
rlabel metal2 2856 11032 2856 11032 0 _0643_
rlabel metal2 1960 6776 1960 6776 0 _0644_
rlabel metal2 2520 7840 2520 7840 0 _0645_
rlabel metal3 3976 19992 3976 19992 0 _0646_
rlabel metal2 3080 20272 3080 20272 0 _0647_
rlabel metal3 25368 9016 25368 9016 0 _0648_
rlabel metal2 24696 11312 24696 11312 0 _0649_
rlabel metal2 12488 18032 12488 18032 0 _0650_
rlabel metal2 6776 7168 6776 7168 0 _0651_
rlabel metal2 3192 7784 3192 7784 0 _0652_
rlabel metal2 14952 17080 14952 17080 0 _0653_
rlabel metal2 12768 16856 12768 16856 0 _0654_
rlabel metal2 3304 13608 3304 13608 0 _0655_
rlabel metal2 16968 29848 16968 29848 0 _0656_
rlabel metal3 28224 14280 28224 14280 0 _0657_
rlabel metal2 7224 15344 7224 15344 0 _0658_
rlabel metal2 25144 17584 25144 17584 0 _0659_
rlabel metal2 9016 3920 9016 3920 0 _0660_
rlabel metal2 12376 27720 12376 27720 0 _0661_
rlabel metal3 13104 27384 13104 27384 0 _0662_
rlabel metal3 12656 30968 12656 30968 0 _0663_
rlabel metal3 12208 33208 12208 33208 0 _0664_
rlabel metal3 14560 44296 14560 44296 0 _0665_
rlabel metal2 24024 38080 24024 38080 0 _0666_
rlabel metal2 3192 22960 3192 22960 0 _0667_
rlabel metal3 6048 23352 6048 23352 0 _0668_
rlabel metal3 19656 4592 19656 4592 0 _0669_
rlabel metal2 1960 18816 1960 18816 0 _0670_
rlabel metal2 26712 17528 26712 17528 0 _0671_
rlabel metal2 3192 27048 3192 27048 0 _0672_
rlabel metal2 2464 30184 2464 30184 0 _0673_
rlabel metal2 13944 9352 13944 9352 0 _0674_
rlabel metal2 16464 8400 16464 8400 0 _0675_
rlabel metal2 20776 20496 20776 20496 0 _0676_
rlabel metal2 17752 23072 17752 23072 0 _0677_
rlabel metal2 3080 24360 3080 24360 0 _0678_
rlabel metal3 6216 23688 6216 23688 0 _0679_
rlabel metal3 15736 19432 15736 19432 0 _0680_
rlabel metal2 16072 22904 16072 22904 0 _0681_
rlabel metal3 9072 15960 9072 15960 0 _0682_
rlabel metal2 2856 18872 2856 18872 0 _0683_
rlabel metal4 16520 22680 16520 22680 0 _0684_
rlabel metal2 22680 25648 22680 25648 0 _0685_
rlabel metal2 4424 23184 4424 23184 0 _0686_
rlabel metal2 2856 30800 2856 30800 0 _0687_
rlabel metal2 7448 9352 7448 9352 0 _0688_
rlabel metal2 6104 16408 6104 16408 0 _0689_
rlabel metal2 6888 6104 6888 6104 0 _0690_
rlabel metal3 4312 23688 4312 23688 0 _0691_
rlabel metal2 3192 10920 3192 10920 0 _0692_
rlabel metal3 2912 15288 2912 15288 0 _0693_
rlabel metal3 2240 21672 2240 21672 0 _0694_
rlabel metal2 3304 7532 3304 7532 0 _0695_
rlabel metal2 16184 8456 16184 8456 0 _0696_
rlabel metal2 3304 23184 3304 23184 0 _0697_
rlabel metal2 3864 21896 3864 21896 0 _0698_
rlabel metal2 5712 23352 5712 23352 0 _0699_
rlabel metal2 26432 16072 26432 16072 0 _0700_
rlabel metal2 1400 6860 1400 6860 0 _0701_
rlabel metal2 22792 7392 22792 7392 0 _0702_
rlabel metal3 15512 2744 15512 2744 0 _0703_
rlabel metal2 7112 14392 7112 14392 0 _0704_
rlabel metal3 6496 12152 6496 12152 0 _0705_
rlabel metal3 6608 28392 6608 28392 0 _0706_
rlabel metal2 23912 18144 23912 18144 0 _0707_
rlabel metal2 23464 7280 23464 7280 0 _0708_
rlabel metal2 24584 20160 24584 20160 0 _0709_
rlabel metal4 23688 16968 23688 16968 0 _0710_
rlabel metal3 23072 17864 23072 17864 0 _0711_
rlabel metal2 24024 19040 24024 19040 0 _0712_
rlabel metal2 26824 19712 26824 19712 0 _0713_
rlabel metal2 19712 16856 19712 16856 0 _0714_
rlabel metal2 24136 20272 24136 20272 0 _0715_
rlabel metal2 5320 30296 5320 30296 0 _0716_
rlabel metal2 5432 32480 5432 32480 0 _0717_
rlabel metal2 8904 35448 8904 35448 0 _0718_
rlabel metal2 20328 35392 20328 35392 0 _0719_
rlabel metal2 6216 36232 6216 36232 0 _0720_
rlabel metal2 7504 43960 7504 43960 0 _0721_
rlabel metal3 7588 44072 7588 44072 0 _0722_
rlabel metal3 19264 45080 19264 45080 0 _0723_
rlabel metal3 18648 18424 18648 18424 0 _0724_
rlabel metal2 2296 18088 2296 18088 0 _0725_
rlabel metal2 9240 23632 9240 23632 0 _0726_
rlabel metal3 10416 8120 10416 8120 0 _0727_
rlabel metal2 8680 7448 8680 7448 0 _0728_
rlabel metal2 19040 12264 19040 12264 0 _0729_
rlabel metal2 12712 19712 12712 19712 0 _0730_
rlabel metal2 17808 24696 17808 24696 0 _0731_
rlabel metal2 3472 16856 3472 16856 0 _0732_
rlabel metal2 5544 23240 5544 23240 0 _0733_
rlabel metal2 4256 22120 4256 22120 0 _0734_
rlabel metal2 2520 24304 2520 24304 0 _0735_
rlabel metal3 4816 22456 4816 22456 0 _0736_
rlabel metal3 8568 35560 8568 35560 0 _0737_
rlabel metal2 10248 35112 10248 35112 0 _0738_
rlabel metal3 11032 34888 11032 34888 0 _0739_
rlabel metal2 23352 55104 23352 55104 0 _0740_
rlabel metal3 10024 34328 10024 34328 0 _0741_
rlabel metal2 9688 40320 9688 40320 0 _0742_
rlabel metal2 7560 40600 7560 40600 0 _0743_
rlabel metal2 7392 39704 7392 39704 0 _0744_
rlabel metal2 8456 33936 8456 33936 0 _0745_
rlabel metal3 3080 23800 3080 23800 0 _0746_
rlabel metal3 11928 12376 11928 12376 0 _0747_
rlabel metal3 8904 22120 8904 22120 0 _0748_
rlabel metal2 3528 44772 3528 44772 0 _0749_
rlabel metal2 2968 11424 2968 11424 0 _0750_
rlabel metal3 6832 22344 6832 22344 0 _0751_
rlabel metal2 7616 22456 7616 22456 0 _0752_
rlabel metal2 17864 26600 17864 26600 0 _0753_
rlabel metal2 1736 24304 1736 24304 0 _0754_
rlabel metal3 22512 12824 22512 12824 0 _0755_
rlabel metal2 26488 21336 26488 21336 0 _0756_
rlabel metal2 23464 25928 23464 25928 0 _0757_
rlabel metal2 24528 25480 24528 25480 0 _0758_
rlabel metal2 23352 15792 23352 15792 0 _0759_
rlabel metal2 21896 18424 21896 18424 0 _0760_
rlabel metal2 30296 21168 30296 21168 0 _0761_
rlabel metal2 24808 26180 24808 26180 0 _0762_
rlabel metal2 24360 25816 24360 25816 0 _0763_
rlabel metal2 18088 29792 18088 29792 0 _0764_
rlabel metal2 10248 28336 10248 28336 0 _0765_
rlabel metal2 15736 6160 15736 6160 0 _0766_
rlabel metal2 6832 20216 6832 20216 0 _0767_
rlabel metal3 7056 27832 7056 27832 0 _0768_
rlabel metal2 6104 34384 6104 34384 0 _0769_
rlabel metal2 7448 38724 7448 38724 0 _0770_
rlabel metal2 7896 33712 7896 33712 0 _0771_
rlabel metal2 6552 33432 6552 33432 0 _0772_
rlabel metal2 1848 26992 1848 26992 0 _0773_
rlabel metal2 6888 25816 6888 25816 0 _0774_
rlabel metal2 13496 13832 13496 13832 0 _0775_
rlabel metal2 8456 25424 8456 25424 0 _0776_
rlabel metal2 25032 19376 25032 19376 0 _0777_
rlabel metal3 7952 40040 7952 40040 0 _0778_
rlabel metal3 6384 30296 6384 30296 0 _0779_
rlabel metal2 7336 37072 7336 37072 0 _0780_
rlabel metal2 7784 38304 7784 38304 0 _0781_
rlabel metal2 20104 25368 20104 25368 0 _0782_
rlabel metal2 18872 27272 18872 27272 0 _0783_
rlabel metal2 11592 20496 11592 20496 0 _0784_
rlabel metal2 1848 18256 1848 18256 0 _0785_
rlabel metal2 2968 18200 2968 18200 0 _0786_
rlabel metal2 7672 20328 7672 20328 0 _0787_
rlabel metal2 2296 14336 2296 14336 0 _0788_
rlabel metal3 7840 20776 7840 20776 0 _0789_
rlabel metal2 8288 25704 8288 25704 0 _0790_
rlabel metal2 25704 22176 25704 22176 0 _0791_
rlabel metal2 11256 18984 11256 18984 0 _0792_
rlabel metal2 25592 22624 25592 22624 0 _0793_
rlabel metal2 23688 22568 23688 22568 0 _0794_
rlabel metal3 25312 23016 25312 23016 0 _0795_
rlabel metal2 20552 18704 20552 18704 0 _0796_
rlabel metal3 21000 24472 21000 24472 0 _0797_
rlabel metal2 27496 22680 27496 22680 0 _0798_
rlabel metal2 26768 22568 26768 22568 0 _0799_
rlabel metal3 11032 29400 11032 29400 0 _0800_
rlabel metal2 10024 28616 10024 28616 0 _0801_
rlabel metal2 8568 29792 8568 29792 0 _0802_
rlabel metal2 11928 36848 11928 36848 0 _0803_
rlabel metal2 9184 36568 9184 36568 0 _0804_
rlabel metal2 7448 37688 7448 37688 0 _0805_
rlabel metal3 9128 39816 9128 39816 0 _0806_
rlabel metal2 12152 32424 12152 32424 0 _0807_
rlabel metal2 22232 15148 22232 15148 0 _0808_
rlabel metal2 1960 15624 1960 15624 0 _0809_
rlabel metal2 2520 15008 2520 15008 0 _0810_
rlabel metal3 12544 15176 12544 15176 0 _0811_
rlabel metal2 17864 5544 17864 5544 0 _0812_
rlabel metal2 13608 15624 13608 15624 0 _0813_
rlabel metal2 15288 14280 15288 14280 0 _0814_
rlabel metal2 13048 15792 13048 15792 0 _0815_
rlabel metal3 25424 15288 25424 15288 0 _0816_
rlabel metal2 15512 13216 15512 13216 0 _0817_
rlabel metal2 2912 20888 2912 20888 0 _0818_
rlabel metal3 12712 26488 12712 26488 0 _0819_
rlabel metal3 13664 31864 13664 31864 0 _0820_
rlabel metal2 11480 33488 11480 33488 0 _0821_
rlabel metal3 10136 41048 10136 41048 0 _0822_
rlabel metal3 18648 44184 18648 44184 0 _0823_
rlabel metal2 4984 40712 4984 40712 0 _0824_
rlabel metal3 9016 41160 9016 41160 0 _0825_
rlabel metal2 3304 41888 3304 41888 0 _0826_
rlabel metal3 10304 38696 10304 38696 0 _0827_
rlabel metal3 5544 44072 5544 44072 0 _0828_
rlabel metal2 7168 40152 7168 40152 0 _0829_
rlabel metal2 6552 40824 6552 40824 0 _0830_
rlabel metal2 4984 35336 4984 35336 0 _0831_
rlabel metal2 6104 12656 6104 12656 0 _0832_
rlabel metal3 21728 17416 21728 17416 0 _0833_
rlabel metal2 27944 9576 27944 9576 0 _0834_
rlabel metal2 19208 11312 19208 11312 0 _0835_
rlabel metal2 15400 4088 15400 4088 0 _0836_
rlabel metal2 8792 13160 8792 13160 0 _0837_
rlabel metal2 2912 8344 2912 8344 0 _0838_
rlabel metal2 16408 24528 16408 24528 0 _0839_
rlabel metal3 10584 12152 10584 12152 0 _0840_
rlabel metal3 9408 12936 9408 12936 0 _0841_
rlabel metal3 7000 30408 7000 30408 0 _0842_
rlabel metal3 5152 37912 5152 37912 0 _0843_
rlabel metal2 10360 19768 10360 19768 0 _0844_
rlabel metal3 15232 19096 15232 19096 0 _0845_
rlabel metal2 9688 21952 9688 21952 0 _0846_
rlabel metal2 10528 23128 10528 23128 0 _0847_
rlabel metal2 3304 16576 3304 16576 0 _0848_
rlabel metal2 16072 16240 16072 16240 0 _0849_
rlabel metal3 17864 17080 17864 17080 0 _0850_
rlabel metal2 2408 13944 2408 13944 0 _0851_
rlabel metal2 7336 13048 7336 13048 0 _0852_
rlabel metal3 17360 15288 17360 15288 0 _0853_
rlabel metal2 18704 10696 18704 10696 0 _0854_
rlabel metal2 3192 14728 3192 14728 0 _0855_
rlabel metal2 10192 17864 10192 17864 0 _0856_
rlabel metal2 22792 18312 22792 18312 0 _0857_
rlabel metal3 19320 23240 19320 23240 0 _0858_
rlabel metal3 11144 23688 11144 23688 0 _0859_
rlabel metal3 12264 33992 12264 33992 0 _0860_
rlabel metal2 23464 32648 23464 32648 0 _0861_
rlabel metal2 16856 39144 16856 39144 0 _0862_
rlabel metal2 22792 39984 22792 39984 0 _0863_
rlabel metal2 14728 11088 14728 11088 0 _0864_
rlabel metal2 18256 10808 18256 10808 0 _0865_
rlabel metal2 21000 19600 21000 19600 0 _0866_
rlabel metal2 20216 21000 20216 21000 0 _0867_
rlabel metal2 21672 16632 21672 16632 0 _0868_
rlabel metal2 20776 18984 20776 18984 0 _0869_
rlabel metal2 19320 18088 19320 18088 0 _0870_
rlabel metal2 19488 16632 19488 16632 0 _0871_
rlabel metal2 15736 29288 15736 29288 0 _0872_
rlabel metal2 15512 39368 15512 39368 0 _0873_
rlabel metal2 22008 39088 22008 39088 0 _0874_
rlabel metal3 9296 37800 9296 37800 0 _0875_
rlabel metal2 3920 16744 3920 16744 0 _0876_
rlabel metal3 21448 15624 21448 15624 0 _0877_
rlabel metal2 22120 16352 22120 16352 0 _0878_
rlabel metal3 21448 16800 21448 16800 0 _0879_
rlabel metal3 24864 19208 24864 19208 0 _0880_
rlabel metal2 23184 16184 23184 16184 0 _0881_
rlabel metal3 18872 16744 18872 16744 0 _0882_
rlabel metal2 18872 34552 18872 34552 0 _0883_
rlabel metal2 16072 37128 16072 37128 0 _0884_
rlabel metal3 15624 40376 15624 40376 0 _0885_
rlabel metal3 17080 40376 17080 40376 0 _0886_
rlabel metal2 14336 38808 14336 38808 0 _0887_
rlabel metal3 10304 37128 10304 37128 0 _0888_
rlabel metal2 4424 39144 4424 39144 0 _0889_
rlabel metal2 5544 38808 5544 38808 0 _0890_
rlabel metal3 12992 32536 12992 32536 0 _0891_
rlabel metal3 14784 17640 14784 17640 0 _0892_
rlabel metal2 15288 25928 15288 25928 0 _0893_
rlabel metal3 24976 24808 24976 24808 0 _0894_
rlabel metal2 15512 18256 15512 18256 0 _0895_
rlabel metal2 20216 17248 20216 17248 0 _0896_
rlabel metal2 16520 17080 16520 17080 0 _0897_
rlabel metal3 20776 2968 20776 2968 0 _0898_
rlabel metal3 14672 9800 14672 9800 0 _0899_
rlabel metal2 11704 17920 11704 17920 0 _0900_
rlabel metal2 16184 17976 16184 17976 0 _0901_
rlabel metal2 16240 21896 16240 21896 0 _0902_
rlabel metal2 11816 33152 11816 33152 0 _0903_
rlabel metal3 6608 41048 6608 41048 0 _0904_
rlabel metal2 6216 40600 6216 40600 0 _0905_
rlabel metal3 3640 41048 3640 41048 0 _0906_
rlabel metal2 5544 41888 5544 41888 0 _0907_
rlabel metal2 2968 41888 2968 41888 0 _0908_
rlabel metal3 1904 4424 1904 4424 0 _0909_
rlabel metal3 5320 38136 5320 38136 0 _0910_
rlabel metal2 3752 41776 3752 41776 0 _0911_
rlabel metal2 6496 7672 6496 7672 0 _0912_
rlabel metal3 7056 7672 7056 7672 0 _0913_
rlabel metal2 6888 8372 6888 8372 0 _0914_
rlabel metal2 8792 17360 8792 17360 0 _0915_
rlabel metal2 10696 11424 10696 11424 0 _0916_
rlabel metal2 15400 7448 15400 7448 0 _0917_
rlabel metal2 13832 11424 13832 11424 0 _0918_
rlabel metal2 17192 23968 17192 23968 0 _0919_
rlabel metal2 1960 9968 1960 9968 0 _0920_
rlabel metal2 16968 11536 16968 11536 0 _0921_
rlabel metal2 8568 33936 8568 33936 0 _0922_
rlabel metal2 4760 33040 4760 33040 0 _0923_
rlabel metal2 9128 37744 9128 37744 0 _0924_
rlabel metal3 8232 17528 8232 17528 0 _0925_
rlabel metal2 18088 18256 18088 18256 0 _0926_
rlabel metal2 18312 18928 18312 18928 0 _0927_
rlabel metal2 18256 17864 18256 17864 0 _0928_
rlabel metal2 19544 5824 19544 5824 0 _0929_
rlabel metal3 19656 12376 19656 12376 0 _0930_
rlabel metal2 18872 12488 18872 12488 0 _0931_
rlabel metal2 18648 13608 18648 13608 0 _0932_
rlabel metal3 16016 38696 16016 38696 0 _0933_
rlabel metal2 16184 37856 16184 37856 0 _0934_
rlabel metal2 16072 38248 16072 38248 0 _0935_
rlabel metal3 15540 37800 15540 37800 0 _0936_
rlabel metal2 11368 38752 11368 38752 0 _0937_
rlabel metal2 11144 42000 11144 42000 0 _0938_
rlabel metal3 11256 42728 11256 42728 0 _0939_
rlabel metal2 10920 43008 10920 43008 0 _0940_
rlabel metal2 16408 32816 16408 32816 0 _0941_
rlabel metal2 15288 32368 15288 32368 0 _0942_
rlabel metal2 25592 18536 25592 18536 0 _0943_
rlabel metal2 2632 19824 2632 19824 0 _0944_
rlabel metal2 18816 24584 18816 24584 0 _0945_
rlabel metal3 21672 20888 21672 20888 0 _0946_
rlabel metal2 16632 22512 16632 22512 0 _0947_
rlabel metal3 19992 21560 19992 21560 0 _0948_
rlabel metal2 17976 19432 17976 19432 0 _0949_
rlabel metal3 21896 21672 21896 21672 0 _0950_
rlabel metal2 22624 21784 22624 21784 0 _0951_
rlabel metal2 23128 25256 23128 25256 0 _0952_
rlabel metal3 23688 23800 23688 23800 0 _0953_
rlabel metal3 23688 23912 23688 23912 0 _0954_
rlabel metal2 18088 31864 18088 31864 0 _0955_
rlabel metal2 12936 43876 12936 43876 0 _0956_
rlabel metal3 5096 42728 5096 42728 0 _0957_
rlabel metal2 2520 42392 2520 42392 0 _0958_
rlabel metal3 2128 5208 2128 5208 0 _0959_
rlabel metal3 11200 43624 11200 43624 0 _0960_
rlabel metal2 10472 45920 10472 45920 0 _0961_
rlabel metal2 19544 42448 19544 42448 0 _0962_
rlabel metal3 7224 31640 7224 31640 0 _0963_
rlabel metal2 8120 28784 8120 28784 0 _0964_
rlabel metal2 15624 26600 15624 26600 0 _0965_
rlabel metal2 10920 26152 10920 26152 0 _0966_
rlabel metal2 11816 16380 11816 16380 0 _0967_
rlabel metal2 11032 21952 11032 21952 0 _0968_
rlabel metal2 10864 31528 10864 31528 0 _0969_
rlabel metal2 8680 31836 8680 31836 0 _0970_
rlabel metal3 9856 39368 9856 39368 0 _0971_
rlabel metal2 8008 33488 8008 33488 0 _0972_
rlabel metal2 7672 33824 7672 33824 0 _0973_
rlabel metal2 11592 40264 11592 40264 0 _0974_
rlabel metal2 14336 35672 14336 35672 0 _0975_
rlabel metal2 14280 18424 14280 18424 0 _0976_
rlabel metal3 9464 20664 9464 20664 0 _0977_
rlabel metal3 12600 20776 12600 20776 0 _0978_
rlabel metal2 21672 19992 21672 19992 0 _0979_
rlabel metal2 14280 21112 14280 21112 0 _0980_
rlabel metal2 16632 19824 16632 19824 0 _0981_
rlabel metal3 17136 20888 17136 20888 0 _0982_
rlabel metal3 17584 21672 17584 21672 0 _0983_
rlabel metal2 18088 25032 18088 25032 0 _0984_
rlabel metal2 15960 34048 15960 34048 0 _0985_
rlabel metal2 15400 35392 15400 35392 0 _0986_
rlabel metal2 13944 40040 13944 40040 0 _0987_
rlabel metal2 20552 39760 20552 39760 0 _0988_
rlabel metal2 12264 20216 12264 20216 0 _0989_
rlabel metal2 12376 20384 12376 20384 0 _0990_
rlabel metal3 10584 20552 10584 20552 0 _0991_
rlabel metal2 18088 19824 18088 19824 0 _0992_
rlabel metal2 12488 22176 12488 22176 0 _0993_
rlabel metal2 18200 37072 18200 37072 0 _0994_
rlabel metal2 14000 37464 14000 37464 0 _0995_
rlabel metal2 14560 39592 14560 39592 0 _0996_
rlabel metal2 13888 41384 13888 41384 0 _0997_
rlabel metal2 13272 41664 13272 41664 0 _0998_
rlabel metal2 12936 42392 12936 42392 0 _0999_
rlabel metal2 16632 25256 16632 25256 0 _1000_
rlabel metal2 16856 27888 16856 27888 0 _1001_
rlabel metal3 23240 16688 23240 16688 0 _1002_
rlabel metal2 20888 24304 20888 24304 0 _1003_
rlabel metal2 20552 24584 20552 24584 0 _1004_
rlabel metal2 22120 24192 22120 24192 0 _1005_
rlabel metal2 18200 28672 18200 28672 0 _1006_
rlabel metal2 18536 31584 18536 31584 0 _1007_
rlabel metal2 16296 32760 16296 32760 0 _1008_
rlabel metal2 14952 40488 14952 40488 0 _1009_
rlabel metal2 11816 46704 11816 46704 0 _1010_
rlabel metal2 9912 47264 9912 47264 0 _1011_
rlabel metal3 6776 42952 6776 42952 0 _1012_
rlabel metal2 7224 45556 7224 45556 0 _1013_
rlabel metal2 7896 42056 7896 42056 0 _1014_
rlabel metal2 6832 42504 6832 42504 0 _1015_
rlabel metal2 7224 42952 7224 42952 0 _1016_
rlabel metal3 9856 47208 9856 47208 0 _1017_
rlabel metal3 25704 42840 25704 42840 0 _1018_
rlabel metal2 14280 41664 14280 41664 0 _1019_
rlabel metal2 14504 41216 14504 41216 0 _1020_
rlabel metal2 14168 48664 14168 48664 0 _1021_
rlabel metal3 7112 16968 7112 16968 0 _1022_
rlabel metal2 7112 29064 7112 29064 0 _1023_
rlabel metal3 29680 23688 29680 23688 0 _1024_
rlabel metal3 26040 25256 26040 25256 0 _1025_
rlabel metal3 20104 29008 20104 29008 0 _1026_
rlabel metal3 7224 28560 7224 28560 0 _1027_
rlabel metal3 6608 29400 6608 29400 0 _1028_
rlabel metal2 8568 30800 8568 30800 0 _1029_
rlabel metal2 10024 33320 10024 33320 0 _1030_
rlabel metal2 7784 30128 7784 30128 0 _1031_
rlabel metal3 9464 31864 9464 31864 0 _1032_
rlabel metal3 9240 33432 9240 33432 0 _1033_
rlabel metal3 11144 44968 11144 44968 0 _1034_
rlabel metal2 16184 15848 16184 15848 0 _1035_
rlabel metal2 16576 13720 16576 13720 0 _1036_
rlabel metal2 16128 13720 16128 13720 0 _1037_
rlabel metal2 17528 15848 17528 15848 0 _1038_
rlabel metal3 24696 15512 24696 15512 0 _1039_
rlabel metal3 17136 15960 17136 15960 0 _1040_
rlabel metal2 19208 15736 19208 15736 0 _1041_
rlabel metal2 21840 10024 21840 10024 0 _1042_
rlabel metal2 18312 16128 18312 16128 0 _1043_
rlabel metal2 17472 39368 17472 39368 0 _1044_
rlabel metal2 17976 37744 17976 37744 0 _1045_
rlabel metal2 18536 38416 18536 38416 0 _1046_
rlabel metal2 17864 40432 17864 40432 0 _1047_
rlabel metal2 21112 39088 21112 39088 0 _1048_
rlabel metal3 17192 38808 17192 38808 0 _1049_
rlabel metal2 14728 45192 14728 45192 0 _1050_
rlabel metal2 12712 47488 12712 47488 0 _1051_
rlabel metal3 11984 47432 11984 47432 0 _1052_
rlabel metal3 12936 48216 12936 48216 0 _1053_
rlabel metal2 24248 26152 24248 26152 0 _1054_
rlabel metal3 19376 26040 19376 26040 0 _1055_
rlabel metal3 18536 26264 18536 26264 0 _1056_
rlabel metal2 19376 26488 19376 26488 0 _1057_
rlabel metal2 18144 20776 18144 20776 0 _1058_
rlabel metal2 11816 24696 11816 24696 0 _1059_
rlabel metal2 1904 24920 1904 24920 0 _1060_
rlabel metal2 11592 25704 11592 25704 0 _1061_
rlabel metal2 16072 28336 16072 28336 0 _1062_
rlabel metal2 19768 29960 19768 29960 0 _1063_
rlabel metal2 22008 30184 22008 30184 0 _1064_
rlabel metal2 19432 31304 19432 31304 0 _1065_
rlabel metal3 19824 31864 19824 31864 0 _1066_
rlabel metal2 14952 47152 14952 47152 0 _1067_
rlabel metal2 10472 49056 10472 49056 0 _1068_
rlabel metal2 11480 48272 11480 48272 0 _1069_
rlabel metal2 10024 49224 10024 49224 0 _1070_
rlabel metal2 9240 50176 9240 50176 0 _1071_
rlabel metal2 13776 46088 13776 46088 0 _1072_
rlabel metal2 13944 49280 13944 49280 0 _1073_
rlabel metal2 16296 47152 16296 47152 0 _1074_
rlabel metal3 25200 21672 25200 21672 0 _1075_
rlabel metal2 18424 24080 18424 24080 0 _1076_
rlabel metal2 27608 21224 27608 21224 0 _1077_
rlabel metal2 27048 19656 27048 19656 0 _1078_
rlabel metal3 27496 21448 27496 21448 0 _1079_
rlabel metal2 27384 23240 27384 23240 0 _1080_
rlabel metal3 21112 33096 21112 33096 0 _1081_
rlabel metal2 17640 33600 17640 33600 0 _1082_
rlabel metal2 15064 44632 15064 44632 0 _1083_
rlabel metal3 18648 44296 18648 44296 0 _1084_
rlabel metal2 13832 29456 13832 29456 0 _1085_
rlabel metal3 14672 30072 14672 30072 0 _1086_
rlabel metal2 12432 23688 12432 23688 0 _1087_
rlabel metal2 12264 23240 12264 23240 0 _1088_
rlabel metal2 12432 24024 12432 24024 0 _1089_
rlabel metal2 15400 30464 15400 30464 0 _1090_
rlabel metal3 16240 41944 16240 41944 0 _1091_
rlabel metal3 15736 43512 15736 43512 0 _1092_
rlabel metal2 15344 42840 15344 42840 0 _1093_
rlabel metal2 15568 43512 15568 43512 0 _1094_
rlabel metal2 16408 44296 16408 44296 0 _1095_
rlabel metal2 23464 40376 23464 40376 0 _1096_
rlabel metal3 20496 25368 20496 25368 0 _1097_
rlabel metal2 17696 25592 17696 25592 0 _1098_
rlabel metal3 14952 40936 14952 40936 0 _1099_
rlabel metal2 16128 43960 16128 43960 0 _1100_
rlabel metal2 16744 47152 16744 47152 0 _1101_
rlabel metal3 18368 48440 18368 48440 0 _1102_
rlabel metal2 15848 49168 15848 49168 0 _1103_
rlabel metal2 13720 49056 13720 49056 0 _1104_
rlabel metal3 13384 48776 13384 48776 0 _1105_
rlabel metal2 12488 49056 12488 49056 0 _1106_
rlabel metal3 14448 49000 14448 49000 0 _1107_
rlabel via2 16296 48440 16296 48440 0 _1108_
rlabel metal3 1904 6664 1904 6664 0 _1109_
rlabel metal2 16968 44016 16968 44016 0 _1110_
rlabel metal2 19320 45584 19320 45584 0 _1111_
rlabel metal2 18312 23464 18312 23464 0 _1112_
rlabel metal2 17752 23352 17752 23352 0 _1113_
rlabel metal2 16296 25928 16296 25928 0 _1114_
rlabel metal2 16968 26488 16968 26488 0 _1115_
rlabel metal2 23072 25592 23072 25592 0 _1116_
rlabel metal2 18704 39368 18704 39368 0 _1117_
rlabel metal3 19544 37240 19544 37240 0 _1118_
rlabel metal2 19880 37408 19880 37408 0 _1119_
rlabel metal2 24024 20664 24024 20664 0 _1120_
rlabel metal2 29624 22400 29624 22400 0 _1121_
rlabel metal3 21392 22456 21392 22456 0 _1122_
rlabel metal2 20944 33096 20944 33096 0 _1123_
rlabel metal2 20664 35728 20664 35728 0 _1124_
rlabel metal3 21056 36344 21056 36344 0 _1125_
rlabel metal3 20608 40376 20608 40376 0 _1126_
rlabel metal2 20272 44632 20272 44632 0 _1127_
rlabel metal2 20104 35784 20104 35784 0 _1128_
rlabel metal2 23744 38696 23744 38696 0 _1129_
rlabel metal2 19880 35336 19880 35336 0 _1130_
rlabel metal3 20608 44968 20608 44968 0 _1131_
rlabel metal2 20384 45304 20384 45304 0 _1132_
rlabel metal2 25144 20720 25144 20720 0 _1133_
rlabel metal3 26544 16072 26544 16072 0 _1134_
rlabel metal2 26152 18424 26152 18424 0 _1135_
rlabel metal3 25536 39368 25536 39368 0 _1136_
rlabel metal2 20776 44408 20776 44408 0 _1137_
rlabel metal2 19544 45024 19544 45024 0 _1138_
rlabel metal2 19656 48272 19656 48272 0 _1139_
rlabel metal3 17640 47208 17640 47208 0 _1140_
rlabel metal3 18816 46536 18816 46536 0 _1141_
rlabel metal4 20216 25536 20216 25536 0 _1142_
rlabel metal2 20104 43120 20104 43120 0 _1143_
rlabel metal3 22008 45192 22008 45192 0 _1144_
rlabel metal2 24976 26152 24976 26152 0 _1145_
rlabel metal3 25312 27048 25312 27048 0 _1146_
rlabel metal2 19432 24528 19432 24528 0 _1147_
rlabel metal2 19208 21952 19208 21952 0 _1148_
rlabel metal2 19320 22792 19320 22792 0 _1149_
rlabel metal2 19824 26824 19824 26824 0 _1150_
rlabel metal2 19096 39200 19096 39200 0 _1151_
rlabel metal2 19712 39816 19712 39816 0 _1152_
rlabel metal2 19544 41272 19544 41272 0 _1153_
rlabel metal2 22904 42448 22904 42448 0 _1154_
rlabel metal2 24696 37632 24696 37632 0 _1155_
rlabel metal3 25816 25368 25816 25368 0 _1156_
rlabel metal3 26040 26936 26040 26936 0 _1157_
rlabel metal3 26376 29400 26376 29400 0 _1158_
rlabel metal2 28168 22232 28168 22232 0 _1159_
rlabel metal2 27664 25368 27664 25368 0 _1160_
rlabel metal3 26376 36232 26376 36232 0 _1161_
rlabel metal2 24976 28056 24976 28056 0 _1162_
rlabel metal2 24360 36624 24360 36624 0 _1163_
rlabel metal3 23744 42840 23744 42840 0 _1164_
rlabel metal2 22848 44296 22848 44296 0 _1165_
rlabel metal2 21672 32200 21672 32200 0 _1166_
rlabel metal2 20104 30576 20104 30576 0 _1167_
rlabel metal2 22288 27832 22288 27832 0 _1168_
rlabel metal2 22120 30464 22120 30464 0 _1169_
rlabel metal2 22456 31472 22456 31472 0 _1170_
rlabel metal3 23408 44296 23408 44296 0 _1171_
rlabel metal2 22904 45584 22904 45584 0 _1172_
rlabel metal3 24024 46648 24024 46648 0 _1173_
rlabel metal3 18144 48328 18144 48328 0 _1174_
rlabel metal2 18872 48496 18872 48496 0 _1175_
rlabel metal2 19208 46200 19208 46200 0 _1176_
rlabel metal2 18200 46872 18200 46872 0 _1177_
rlabel metal3 19040 47544 19040 47544 0 _1178_
rlabel metal2 24920 47320 24920 47320 0 _1179_
rlabel metal2 26488 48944 26488 48944 0 _1180_
rlabel metal2 25928 44464 25928 44464 0 _1181_
rlabel metal3 23856 43512 23856 43512 0 _1182_
rlabel metal2 26040 44576 26040 44576 0 _1183_
rlabel metal2 26264 21672 26264 21672 0 _1184_
rlabel metal2 25704 23352 25704 23352 0 _1185_
rlabel metal3 21784 39368 21784 39368 0 _1186_
rlabel metal2 21672 39872 21672 39872 0 _1187_
rlabel metal3 21560 39704 21560 39704 0 _1188_
rlabel metal2 20664 41272 20664 41272 0 _1189_
rlabel metal2 25928 41384 25928 41384 0 _1190_
rlabel metal3 28728 24696 28728 24696 0 _1191_
rlabel metal2 28168 25144 28168 25144 0 _1192_
rlabel metal2 25928 37408 25928 37408 0 _1193_
rlabel metal2 25592 37632 25592 37632 0 _1194_
rlabel metal2 26040 39424 26040 39424 0 _1195_
rlabel metal2 24808 29456 24808 29456 0 _1196_
rlabel metal3 25592 31080 25592 31080 0 _1197_
rlabel metal3 25088 30968 25088 30968 0 _1198_
rlabel metal2 26544 41944 26544 41944 0 _1199_
rlabel metal3 25144 44408 25144 44408 0 _1200_
rlabel metal2 26712 44632 26712 44632 0 _1201_
rlabel metal3 24080 45864 24080 45864 0 _1202_
rlabel metal3 25480 45976 25480 45976 0 _1203_
rlabel metal2 57848 45584 57848 45584 0 _1204_
rlabel metal2 10136 26208 10136 26208 0 _1205_
rlabel metal2 3304 36372 3304 36372 0 _1206_
rlabel metal2 18088 43904 18088 43904 0 _1207_
rlabel metal2 20664 49728 20664 49728 0 _1208_
rlabel metal2 25480 32816 25480 32816 0 _1209_
rlabel metal2 24360 38248 24360 38248 0 _1210_
rlabel metal3 25144 48104 25144 48104 0 _1211_
rlabel metal3 21896 49784 21896 49784 0 _1212_
rlabel metal3 23688 46872 23688 46872 0 _1213_
rlabel metal3 24584 50568 24584 50568 0 _1214_
rlabel metal2 26040 41664 26040 41664 0 _1215_
rlabel metal2 25704 40600 25704 40600 0 _1216_
rlabel metal2 26152 50512 26152 50512 0 _1217_
rlabel metal2 27384 50904 27384 50904 0 _1218_
rlabel metal2 26544 45304 26544 45304 0 _1219_
rlabel metal3 25480 44072 25480 44072 0 _1220_
rlabel metal2 25480 46368 25480 46368 0 _1221_
rlabel metal2 24248 44968 24248 44968 0 _1222_
rlabel metal2 26712 49336 26712 49336 0 _1223_
rlabel metal2 28056 52360 28056 52360 0 _1224_
rlabel metal2 23688 49000 23688 49000 0 _1225_
rlabel metal2 23576 49784 23576 49784 0 _1226_
rlabel metal2 23800 49896 23800 49896 0 _1227_
rlabel metal3 22624 40936 22624 40936 0 _1228_
rlabel metal3 27776 27944 27776 27944 0 _1229_
rlabel metal3 22400 38920 22400 38920 0 _1230_
rlabel metal3 21728 38696 21728 38696 0 _1231_
rlabel metal2 22680 41048 22680 41048 0 _1232_
rlabel metal2 22568 46368 22568 46368 0 _1233_
rlabel metal3 23184 48328 23184 48328 0 _1234_
rlabel metal3 24024 47320 24024 47320 0 _1235_
rlabel metal3 23800 48216 23800 48216 0 _1236_
rlabel metal2 23408 49560 23408 49560 0 _1237_
rlabel metal3 25928 49896 25928 49896 0 _1238_
rlabel metal3 25200 51128 25200 51128 0 _1239_
rlabel metal2 27944 49392 27944 49392 0 _1240_
rlabel metal2 3304 49168 3304 49168 0 _1241_
rlabel metal2 27272 48944 27272 48944 0 _1242_
rlabel metal2 24136 51576 24136 51576 0 _1243_
rlabel metal2 24584 50456 24584 50456 0 _1244_
rlabel metal2 24920 50064 24920 50064 0 _1245_
rlabel metal3 22680 47432 22680 47432 0 _1246_
rlabel metal3 25256 47432 25256 47432 0 _1247_
rlabel metal2 26152 48048 26152 48048 0 _1248_
rlabel metal2 10472 41496 10472 41496 0 _1249_
rlabel metal2 48440 20440 48440 20440 0 _1250_
rlabel metal2 46760 13328 46760 13328 0 _1251_
rlabel metal2 45864 17192 45864 17192 0 _1252_
rlabel metal2 45752 24696 45752 24696 0 _1253_
rlabel metal3 43904 19320 43904 19320 0 _1254_
rlabel metal2 56560 17640 56560 17640 0 _1255_
rlabel metal2 46984 18592 46984 18592 0 _1256_
rlabel metal2 45472 23128 45472 23128 0 _1257_
rlabel metal2 53368 11928 53368 11928 0 _1258_
rlabel metal3 44296 23128 44296 23128 0 _1259_
rlabel metal3 49280 29400 49280 29400 0 _1260_
rlabel metal2 50064 25704 50064 25704 0 _1261_
rlabel metal2 41608 26488 41608 26488 0 _1262_
rlabel metal3 47208 12936 47208 12936 0 _1263_
rlabel metal2 50008 17192 50008 17192 0 _1264_
rlabel metal2 52248 15344 52248 15344 0 _1265_
rlabel metal3 47712 16856 47712 16856 0 _1266_
rlabel metal2 45528 24696 45528 24696 0 _1267_
rlabel metal2 44744 9128 44744 9128 0 _1268_
rlabel metal2 54152 11312 54152 11312 0 _1269_
rlabel metal3 47992 17360 47992 17360 0 _1270_
rlabel metal3 45472 18984 45472 18984 0 _1271_
rlabel metal2 57960 25760 57960 25760 0 _1272_
rlabel metal3 41384 20776 41384 20776 0 _1273_
rlabel metal2 46648 18984 46648 18984 0 _1274_
rlabel metal3 42056 21000 42056 21000 0 _1275_
rlabel metal2 43176 22624 43176 22624 0 _1276_
rlabel metal3 58184 42504 58184 42504 0 _1277_
rlabel metal2 43792 23128 43792 23128 0 _1278_
rlabel metal2 43288 22904 43288 22904 0 _1279_
rlabel metal2 47544 19656 47544 19656 0 _1280_
rlabel metal2 57568 31752 57568 31752 0 _1281_
rlabel metal2 46760 24752 46760 24752 0 _1282_
rlabel metal2 42168 25928 42168 25928 0 _1283_
rlabel metal3 58128 20104 58128 20104 0 _1284_
rlabel metal2 55272 31808 55272 31808 0 _1285_
rlabel metal4 43064 24304 43064 24304 0 _1286_
rlabel metal2 46200 19824 46200 19824 0 _1287_
rlabel metal2 43176 24304 43176 24304 0 _1288_
rlabel metal2 57680 21560 57680 21560 0 _1289_
rlabel metal2 53480 21896 53480 21896 0 _1290_
rlabel metal2 52920 40936 52920 40936 0 _1291_
rlabel metal2 48608 15624 48608 15624 0 _1292_
rlabel metal2 46200 12824 46200 12824 0 _1293_
rlabel metal2 45584 13720 45584 13720 0 _1294_
rlabel metal3 43624 25256 43624 25256 0 _1295_
rlabel metal3 56392 19096 56392 19096 0 _1296_
rlabel metal2 46088 15848 46088 15848 0 _1297_
rlabel metal2 55720 14056 55720 14056 0 _1298_
rlabel metal2 49672 14056 49672 14056 0 _1299_
rlabel metal3 54992 15064 54992 15064 0 _1300_
rlabel metal2 49336 16128 49336 16128 0 _1301_
rlabel metal2 57848 25984 57848 25984 0 _1302_
rlabel metal3 50456 16072 50456 16072 0 _1303_
rlabel metal2 45864 15960 45864 15960 0 _1304_
rlabel metal4 42728 23744 42728 23744 0 _1305_
rlabel metal2 34888 25424 34888 25424 0 _1306_
rlabel metal3 44352 26264 44352 26264 0 _1307_
rlabel metal2 49336 15512 49336 15512 0 _1308_
rlabel metal2 34216 27496 34216 27496 0 _1309_
rlabel metal2 32424 45192 32424 45192 0 _1310_
rlabel metal2 48720 52136 48720 52136 0 _1311_
rlabel metal2 39816 49336 39816 49336 0 _1312_
rlabel metal3 57148 26824 57148 26824 0 _1313_
rlabel metal2 44408 51688 44408 51688 0 _1314_
rlabel metal2 40712 50120 40712 50120 0 _1315_
rlabel metal2 45640 24360 45640 24360 0 _1316_
rlabel metal2 41552 10808 41552 10808 0 _1317_
rlabel metal2 49840 18648 49840 18648 0 _1318_
rlabel metal2 49392 24696 49392 24696 0 _1319_
rlabel metal2 46088 21560 46088 21560 0 _1320_
rlabel metal2 51576 23968 51576 23968 0 _1321_
rlabel metal3 46256 25480 46256 25480 0 _1322_
rlabel metal3 56896 14504 56896 14504 0 _1323_
rlabel metal2 46984 15680 46984 15680 0 _1324_
rlabel metal2 55328 40152 55328 40152 0 _1325_
rlabel metal2 45080 25032 45080 25032 0 _1326_
rlabel metal2 55160 22848 55160 22848 0 _1327_
rlabel metal3 43064 21784 43064 21784 0 _1328_
rlabel metal2 45192 24696 45192 24696 0 _1329_
rlabel metal2 44968 33880 44968 33880 0 _1330_
rlabel metal2 48328 19712 48328 19712 0 _1331_
rlabel metal2 43400 17976 43400 17976 0 _1332_
rlabel metal2 46424 20776 46424 20776 0 _1333_
rlabel metal3 43400 20776 43400 20776 0 _1334_
rlabel metal3 52136 19992 52136 19992 0 _1335_
rlabel metal2 42504 21336 42504 21336 0 _1336_
rlabel metal3 43960 20664 43960 20664 0 _1337_
rlabel metal3 42896 36232 42896 36232 0 _1338_
rlabel metal2 56448 34216 56448 34216 0 _1339_
rlabel metal2 55496 15736 55496 15736 0 _1340_
rlabel metal2 58016 24920 58016 24920 0 _1341_
rlabel metal2 37464 36680 37464 36680 0 _1342_
rlabel metal3 47600 37800 47600 37800 0 _1343_
rlabel metal2 47768 34272 47768 34272 0 _1344_
rlabel metal3 40320 31080 40320 31080 0 _1345_
rlabel metal2 57680 16856 57680 16856 0 _1346_
rlabel metal2 46536 31864 46536 31864 0 _1347_
rlabel metal3 46088 20216 46088 20216 0 _1348_
rlabel metal3 44968 32536 44968 32536 0 _1349_
rlabel metal2 33544 24528 33544 24528 0 _1350_
rlabel metal2 39088 16072 39088 16072 0 _1351_
rlabel metal3 40488 22344 40488 22344 0 _1352_
rlabel metal2 57512 23632 57512 23632 0 _1353_
rlabel metal3 48384 23688 48384 23688 0 _1354_
rlabel metal2 43848 30408 43848 30408 0 _1355_
rlabel metal2 44184 32760 44184 32760 0 _1356_
rlabel metal2 53480 17696 53480 17696 0 _1357_
rlabel metal2 44520 39200 44520 39200 0 _1358_
rlabel metal2 48104 48608 48104 48608 0 _1359_
rlabel metal3 55776 15736 55776 15736 0 _1360_
rlabel metal2 55608 16744 55608 16744 0 _1361_
rlabel metal2 54656 9240 54656 9240 0 _1362_
rlabel metal3 39424 16184 39424 16184 0 _1363_
rlabel metal2 43120 26264 43120 26264 0 _1364_
rlabel metal2 42784 16856 42784 16856 0 _1365_
rlabel metal2 50848 20888 50848 20888 0 _1366_
rlabel metal2 53368 43176 53368 43176 0 _1367_
rlabel metal3 55944 15848 55944 15848 0 _1368_
rlabel metal4 47936 21672 47936 21672 0 _1369_
rlabel metal2 55496 19600 55496 19600 0 _1370_
rlabel metal2 55552 20216 55552 20216 0 _1371_
rlabel metal2 47656 16352 47656 16352 0 _1372_
rlabel metal2 54992 17080 54992 17080 0 _1373_
rlabel metal3 54880 22344 54880 22344 0 _1374_
rlabel metal3 39760 34888 39760 34888 0 _1375_
rlabel metal2 55720 22456 55720 22456 0 _1376_
rlabel metal3 57064 7672 57064 7672 0 _1377_
rlabel metal2 55608 44912 55608 44912 0 _1378_
rlabel metal2 53592 16800 53592 16800 0 _1379_
rlabel metal2 53480 42168 53480 42168 0 _1380_
rlabel metal2 51576 47824 51576 47824 0 _1381_
rlabel metal2 41720 47880 41720 47880 0 _1382_
rlabel metal2 36960 46760 36960 46760 0 _1383_
rlabel metal3 33096 46536 33096 46536 0 _1384_
rlabel metal2 3360 45304 3360 45304 0 _1385_
rlabel metal2 35112 43064 35112 43064 0 _1386_
rlabel metal2 43848 53200 43848 53200 0 _1387_
rlabel metal2 40824 29288 40824 29288 0 _1388_
rlabel metal4 48664 19376 48664 19376 0 _1389_
rlabel metal2 49840 10808 49840 10808 0 _1390_
rlabel metal3 48608 25032 48608 25032 0 _1391_
rlabel metal2 48664 28560 48664 28560 0 _1392_
rlabel metal2 46760 31696 46760 31696 0 _1393_
rlabel metal3 43008 24360 43008 24360 0 _1394_
rlabel metal2 38864 23352 38864 23352 0 _1395_
rlabel metal2 44296 31360 44296 31360 0 _1396_
rlabel metal2 46368 32760 46368 32760 0 _1397_
rlabel metal2 49672 12320 49672 12320 0 _1398_
rlabel metal2 47656 20496 47656 20496 0 _1399_
rlabel metal3 39984 25480 39984 25480 0 _1400_
rlabel metal2 47544 30408 47544 30408 0 _1401_
rlabel metal2 41832 33320 41832 33320 0 _1402_
rlabel metal2 48776 13440 48776 13440 0 _1403_
rlabel metal2 38696 15624 38696 15624 0 _1404_
rlabel metal2 41664 33320 41664 33320 0 _1405_
rlabel metal3 49672 22344 49672 22344 0 _1406_
rlabel metal2 50008 34384 50008 34384 0 _1407_
rlabel metal4 40600 28280 40600 28280 0 _1408_
rlabel metal2 41608 33096 41608 33096 0 _1409_
rlabel metal2 46760 36064 46760 36064 0 _1410_
rlabel metal3 40432 19880 40432 19880 0 _1411_
rlabel metal2 43064 36848 43064 36848 0 _1412_
rlabel metal2 43176 35952 43176 35952 0 _1413_
rlabel metal2 41608 47992 41608 47992 0 _1414_
rlabel metal2 39144 52976 39144 52976 0 _1415_
rlabel metal2 49504 51352 49504 51352 0 _1416_
rlabel metal3 47656 50456 47656 50456 0 _1417_
rlabel metal2 42504 50456 42504 50456 0 _1418_
rlabel metal2 42784 51240 42784 51240 0 _1419_
rlabel metal2 46816 34104 46816 34104 0 _1420_
rlabel metal2 46424 34552 46424 34552 0 _1421_
rlabel metal2 46088 35112 46088 35112 0 _1422_
rlabel metal2 50232 44352 50232 44352 0 _1423_
rlabel metal3 53704 48216 53704 48216 0 _1424_
rlabel metal2 35336 20496 35336 20496 0 _1425_
rlabel metal2 49784 26096 49784 26096 0 _1426_
rlabel metal2 50344 25480 50344 25480 0 _1427_
rlabel metal2 49952 27720 49952 27720 0 _1428_
rlabel metal3 57456 18648 57456 18648 0 _1429_
rlabel metal2 57120 24024 57120 24024 0 _1430_
rlabel metal2 57624 28616 57624 28616 0 _1431_
rlabel metal3 18256 6664 18256 6664 0 _1432_
rlabel metal3 58408 16744 58408 16744 0 _1433_
rlabel metal3 57624 28504 57624 28504 0 _1434_
rlabel metal2 56168 28952 56168 28952 0 _1435_
rlabel metal3 55384 48104 55384 48104 0 _1436_
rlabel metal3 54264 47432 54264 47432 0 _1437_
rlabel metal2 45808 51240 45808 51240 0 _1438_
rlabel metal3 44632 50008 44632 50008 0 _1439_
rlabel metal3 50400 8904 50400 8904 0 _1440_
rlabel metal2 51016 22456 51016 22456 0 _1441_
rlabel metal2 44464 22120 44464 22120 0 _1442_
rlabel metal3 16968 7448 16968 7448 0 _1443_
rlabel metal2 16856 854 16856 854 0 addI[0]
rlabel metal2 22904 2058 22904 2058 0 addI[1]
rlabel metal3 57666 20216 57666 20216 0 addI[2]
rlabel metal3 28840 3416 28840 3416 0 addI[3]
rlabel metal3 57666 54488 57666 54488 0 addI[4]
rlabel metal3 58856 56168 58856 56168 0 addI[5]
rlabel metal2 19544 57722 19544 57722 0 addQ[0]
rlabel metal2 25760 56168 25760 56168 0 addQ[1]
rlabel metal2 40376 2058 40376 2058 0 addQ[2]
rlabel metal3 1358 22904 1358 22904 0 addQ[3]
rlabel metal3 1358 57176 1358 57176 0 addQ[4]
rlabel metal2 56056 25872 56056 25872 0 addQ[5]
rlabel metal3 40880 12712 40880 12712 0 bit2symb.regi
rlabel metal2 42168 5824 42168 5824 0 clknet_0_CLK
rlabel metal2 40824 5208 40824 5208 0 clknet_1_0__leaf_CLK
rlabel metal3 49112 3640 49112 3640 0 clknet_1_1__leaf_CLK
rlabel metal3 2352 17752 2352 17752 0 net1
rlabel metal3 47936 56056 47936 56056 0 net10
rlabel metal2 34216 4200 34216 4200 0 net11
rlabel metal2 56168 43792 56168 43792 0 net12
rlabel metal2 56168 8456 56168 8456 0 net13
rlabel metal2 20216 3808 20216 3808 0 net14
rlabel metal2 2408 39928 2408 39928 0 net15
rlabel metal2 2968 29120 2968 29120 0 net16
rlabel metal2 23688 55496 23688 55496 0 net17
rlabel metal2 29960 55664 29960 55664 0 net18
rlabel metal2 2352 48328 2352 48328 0 net19
rlabel metal2 34888 16520 34888 16520 0 net2
rlabel metal3 42448 50680 42448 50680 0 net20
rlabel metal2 9800 46984 9800 46984 0 net21
rlabel metal2 2408 3976 2408 3976 0 net22
rlabel metal2 2800 12712 2800 12712 0 net23
rlabel metal2 45416 42000 45416 42000 0 net24
rlabel metal2 8904 53200 8904 53200 0 net25
rlabel metal2 2408 6160 2408 6160 0 net26
rlabel metal3 51688 3528 51688 3528 0 net27
rlabel metal2 27160 55216 27160 55216 0 net28
rlabel metal2 58240 41608 58240 41608 0 net29
rlabel metal3 41328 7336 41328 7336 0 net3
rlabel metal2 19320 3752 19320 3752 0 net30
rlabel metal2 25368 3696 25368 3696 0 net31
rlabel metal2 49112 7336 49112 7336 0 net32
rlabel metal2 40264 4872 40264 4872 0 net33
rlabel metal3 54768 55272 54768 55272 0 net34
rlabel metal3 56896 53816 56896 53816 0 net35
rlabel metal2 21056 56056 21056 56056 0 net36
rlabel metal3 27664 55944 27664 55944 0 net37
rlabel metal2 24920 4368 24920 4368 0 net38
rlabel metal2 2632 4928 2632 4928 0 net39
rlabel metal2 2408 45584 2408 45584 0 net4
rlabel metal3 3808 55048 3808 55048 0 net40
rlabel metal3 54880 26264 54880 26264 0 net41
rlabel metal3 41440 15176 41440 15176 0 net42
rlabel metal2 49560 45248 49560 45248 0 net43
rlabel metal3 29344 23800 29344 23800 0 net44
rlabel metal2 4200 30800 4200 30800 0 net45
rlabel metal2 21784 6272 21784 6272 0 net46
rlabel metal3 56896 35448 56896 35448 0 net47
rlabel metal2 5768 44072 5768 44072 0 net48
rlabel metal2 25144 34104 25144 34104 0 net49
rlabel metal2 55944 4200 55944 4200 0 net5
rlabel metal3 12376 45080 12376 45080 0 net50
rlabel metal2 44800 6104 44800 6104 0 net51
rlabel metal2 41048 10360 41048 10360 0 net52
rlabel metal2 46200 3752 46200 3752 0 net53
rlabel metal2 48328 7280 48328 7280 0 net54
rlabel metal2 48328 9800 48328 9800 0 net55
rlabel metal2 45640 5600 45640 5600 0 net56
rlabel metal2 38752 43736 38752 43736 0 net57
rlabel metal2 50008 49616 50008 49616 0 net58
rlabel metal2 41944 4872 41944 4872 0 net59
rlabel metal2 56168 4368 56168 4368 0 net6
rlabel metal3 57008 39368 57008 39368 0 net7
rlabel metal2 4200 56168 4200 56168 0 net8
rlabel metal2 2408 52808 2408 52808 0 net9
rlabel metal2 49672 39928 49672 39928 0 p_shaping_I.bit_in
rlabel metal2 49896 40712 49896 40712 0 p_shaping_I.bit_in_1
rlabel metal3 53032 45752 53032 45752 0 p_shaping_I.bit_in_2
rlabel metal3 39088 51240 39088 51240 0 p_shaping_I.counter\[0\]
rlabel metal2 39424 46648 39424 46648 0 p_shaping_I.counter\[1\]
rlabel metal3 32144 34664 32144 34664 0 p_shaping_I.ctl_1
rlabel metal2 24920 35056 24920 35056 0 p_shaping_Q.bit_in_1
rlabel metal2 24136 35336 24136 35336 0 p_shaping_Q.bit_in_2
rlabel metal2 6384 44184 6384 44184 0 p_shaping_Q.counter\[0\]
rlabel metal2 8568 44576 8568 44576 0 p_shaping_Q.counter\[1\]
rlabel metal2 27720 31304 27720 31304 0 p_shaping_Q.ctl_1
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
