VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OQPSK_PS_RCOSINE2
  CLASS BLOCK ;
  FOREIGN OQPSK_PS_RCOSINE2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 300.000 BY 300.000 ;
  PIN BitIn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 84.000 4.000 84.560 ;
    END
  END BitIn
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1.000 229.040 4.000 ;
    END
  END CLK
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 296.000 158.480 299.000 ;
    END
  END EN
  PIN I[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.480 4.000 229.040 ;
    END
  END I[0]
  PIN I[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 285.600 1.000 286.160 4.000 ;
    END
  END I[10]
  PIN I[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 13.440 299.000 14.000 ;
    END
  END I[11]
  PIN I[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 184.800 299.000 185.360 ;
    END
  END I[12]
  PIN I[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 13.440 296.000 14.000 299.000 ;
    END
  END I[1]
  PIN I[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.720 4.000 259.280 ;
    END
  END I[2]
  PIN I[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 296.000 242.480 299.000 ;
    END
  END I[3]
  PIN I[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1.000 171.920 4.000 ;
    END
  END I[4]
  PIN I[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 215.040 299.000 215.600 ;
    END
  END I[5]
  PIN I[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 40.320 299.000 40.880 ;
    END
  END I[6]
  PIN I[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 1.000 57.680 4.000 ;
    END
  END I[7]
  PIN I[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 198.240 4.000 198.800 ;
    END
  END I[8]
  PIN I[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 141.120 4.000 141.680 ;
    END
  END I[9]
  PIN Q[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 296.000 185.360 299.000 ;
    END
  END Q[0]
  PIN Q[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 296.000 272.720 299.000 ;
    END
  END Q[10]
  PIN Q[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 171.360 4.000 171.920 ;
    END
  END Q[11]
  PIN Q[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 241.920 299.000 242.480 ;
    END
  END Q[12]
  PIN Q[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 70.560 296.000 71.120 299.000 ;
    END
  END Q[1]
  PIN Q[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END Q[2]
  PIN Q[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 57.120 4.000 57.680 ;
    END
  END Q[3]
  PIN Q[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 157.920 299.000 158.480 ;
    END
  END Q[4]
  PIN Q[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 296.000 40.880 299.000 ;
    END
  END Q[5]
  PIN Q[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.880 4.000 27.440 ;
    END
  END Q[6]
  PIN Q[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1.000 259.280 4.000 ;
    END
  END Q[7]
  PIN Q[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 215.040 296.000 215.600 299.000 ;
    END
  END Q[8]
  PIN Q[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 70.560 299.000 71.120 ;
    END
  END Q[9]
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1.000 27.440 4.000 ;
    END
  END RST
  PIN addI[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1.000 84.560 4.000 ;
    END
  END addI[0]
  PIN addI[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1.000 114.800 4.000 ;
    END
  END addI[1]
  PIN addI[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 100.800 299.000 101.360 ;
    END
  END addI[2]
  PIN addI[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 1.000 141.680 4.000 ;
    END
  END addI[3]
  PIN addI[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 272.160 299.000 272.720 ;
    END
  END addI[4]
  PIN addI[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 296.000 299.600 299.000 ;
    END
  END addI[5]
  PIN addQ[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 296.000 98.000 299.000 ;
    END
  END addQ[0]
  PIN addQ[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 296.000 128.240 299.000 ;
    END
  END addQ[1]
  PIN addQ[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 1.000 202.160 4.000 ;
    END
  END addQ[2]
  PIN addQ[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 114.240 4.000 114.800 ;
    END
  END addQ[3]
  PIN addQ[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 285.600 4.000 286.160 ;
    END
  END addQ[4]
  PIN addQ[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 296.000 127.680 299.000 128.240 ;
    END
  END addQ[5]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 282.540 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 282.540 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 282.540 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 298.390 283.210 ;
      LAYER Metal2 ;
        RECT 0.140 295.700 13.140 296.000 ;
        RECT 14.300 295.700 40.020 296.000 ;
        RECT 41.180 295.700 70.260 296.000 ;
        RECT 71.420 295.700 97.140 296.000 ;
        RECT 98.300 295.700 127.380 296.000 ;
        RECT 128.540 295.700 157.620 296.000 ;
        RECT 158.780 295.700 184.500 296.000 ;
        RECT 185.660 295.700 214.740 296.000 ;
        RECT 215.900 295.700 241.620 296.000 ;
        RECT 242.780 295.700 271.860 296.000 ;
        RECT 273.020 295.700 298.740 296.000 ;
        RECT 0.140 4.300 299.460 295.700 ;
        RECT 0.860 3.500 26.580 4.300 ;
        RECT 27.740 3.500 56.820 4.300 ;
        RECT 57.980 3.500 83.700 4.300 ;
        RECT 84.860 3.500 113.940 4.300 ;
        RECT 115.100 3.500 140.820 4.300 ;
        RECT 141.980 3.500 171.060 4.300 ;
        RECT 172.220 3.500 201.300 4.300 ;
        RECT 202.460 3.500 228.180 4.300 ;
        RECT 229.340 3.500 258.420 4.300 ;
        RECT 259.580 3.500 285.300 4.300 ;
        RECT 286.460 3.500 299.460 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 285.300 0.700 286.020 ;
        RECT 4.300 285.300 299.510 286.020 ;
        RECT 0.090 273.020 299.510 285.300 ;
        RECT 0.090 271.860 295.700 273.020 ;
        RECT 299.300 271.860 299.510 273.020 ;
        RECT 0.090 259.580 299.510 271.860 ;
        RECT 0.090 258.420 0.700 259.580 ;
        RECT 4.300 258.420 299.510 259.580 ;
        RECT 0.090 242.780 299.510 258.420 ;
        RECT 0.090 241.620 295.700 242.780 ;
        RECT 299.300 241.620 299.510 242.780 ;
        RECT 0.090 229.340 299.510 241.620 ;
        RECT 0.090 228.180 0.700 229.340 ;
        RECT 4.300 228.180 299.510 229.340 ;
        RECT 0.090 215.900 299.510 228.180 ;
        RECT 0.090 214.740 295.700 215.900 ;
        RECT 299.300 214.740 299.510 215.900 ;
        RECT 0.090 199.100 299.510 214.740 ;
        RECT 0.090 197.940 0.700 199.100 ;
        RECT 4.300 197.940 299.510 199.100 ;
        RECT 0.090 185.660 299.510 197.940 ;
        RECT 0.090 184.500 295.700 185.660 ;
        RECT 299.300 184.500 299.510 185.660 ;
        RECT 0.090 172.220 299.510 184.500 ;
        RECT 0.090 171.060 0.700 172.220 ;
        RECT 4.300 171.060 299.510 172.220 ;
        RECT 0.090 158.780 299.510 171.060 ;
        RECT 0.090 157.620 295.700 158.780 ;
        RECT 299.300 157.620 299.510 158.780 ;
        RECT 0.090 141.980 299.510 157.620 ;
        RECT 0.090 140.820 0.700 141.980 ;
        RECT 4.300 140.820 299.510 141.980 ;
        RECT 0.090 128.540 299.510 140.820 ;
        RECT 0.090 127.380 295.700 128.540 ;
        RECT 299.300 127.380 299.510 128.540 ;
        RECT 0.090 115.100 299.510 127.380 ;
        RECT 0.090 113.940 0.700 115.100 ;
        RECT 4.300 113.940 299.510 115.100 ;
        RECT 0.090 101.660 299.510 113.940 ;
        RECT 0.090 100.500 295.700 101.660 ;
        RECT 299.300 100.500 299.510 101.660 ;
        RECT 0.090 84.860 299.510 100.500 ;
        RECT 0.090 83.700 0.700 84.860 ;
        RECT 4.300 83.700 299.510 84.860 ;
        RECT 0.090 71.420 299.510 83.700 ;
        RECT 0.090 70.260 295.700 71.420 ;
        RECT 299.300 70.260 299.510 71.420 ;
        RECT 0.090 57.980 299.510 70.260 ;
        RECT 0.090 56.820 0.700 57.980 ;
        RECT 4.300 56.820 299.510 57.980 ;
        RECT 0.090 41.180 299.510 56.820 ;
        RECT 0.090 40.020 295.700 41.180 ;
        RECT 299.300 40.020 299.510 41.180 ;
        RECT 0.090 27.740 299.510 40.020 ;
        RECT 0.090 26.580 0.700 27.740 ;
        RECT 4.300 26.580 299.510 27.740 ;
        RECT 0.090 14.300 299.510 26.580 ;
        RECT 0.090 13.140 295.700 14.300 ;
        RECT 299.300 13.140 299.510 14.300 ;
        RECT 0.090 6.300 299.510 13.140 ;
      LAYER Metal4 ;
        RECT 10.220 15.080 21.940 279.910 ;
        RECT 24.140 15.080 98.740 279.910 ;
        RECT 100.940 15.080 175.540 279.910 ;
        RECT 177.740 15.080 252.340 279.910 ;
        RECT 254.540 15.080 288.820 279.910 ;
        RECT 10.220 7.370 288.820 15.080 ;
  END
END OQPSK_PS_RCOSINE2
END LIBRARY

